module real_aes_6421_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_0), .A2(n_76), .B1(n_391), .B2(n_393), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_1), .A2(n_175), .B1(n_311), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_2), .A2(n_41), .B1(n_481), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_3), .A2(n_258), .B1(n_572), .B2(n_662), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_4), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_5), .A2(n_266), .B1(n_355), .B2(n_358), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_6), .A2(n_99), .B1(n_388), .B2(n_389), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_7), .A2(n_125), .B1(n_522), .B2(n_526), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_8), .A2(n_130), .B1(n_492), .B2(n_599), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_9), .A2(n_101), .B1(n_381), .B2(n_744), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_10), .A2(n_230), .B1(n_479), .B2(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_11), .Y(n_873) );
INVx1_ASAP7_75t_L g753 ( .A(n_12), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_13), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_14), .A2(n_32), .B1(n_441), .B2(n_481), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g849 ( .A1(n_15), .A2(n_127), .B1(n_850), .B2(n_851), .C(n_852), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_16), .A2(n_145), .B1(n_741), .B2(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_17), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_18), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_19), .A2(n_132), .B1(n_375), .B2(n_376), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_20), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_21), .A2(n_153), .B1(n_680), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_22), .A2(n_28), .B1(n_481), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_23), .A2(n_131), .B1(n_342), .B2(n_572), .Y(n_794) );
AO22x2_ASAP7_75t_L g294 ( .A1(n_24), .A2(n_93), .B1(n_295), .B2(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g819 ( .A(n_24), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_25), .A2(n_83), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_26), .A2(n_44), .B1(n_355), .B2(n_672), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_27), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_29), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_30), .A2(n_216), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_31), .A2(n_259), .B1(n_389), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_33), .A2(n_192), .B1(n_393), .B2(n_440), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_34), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_35), .A2(n_136), .B1(n_362), .B2(n_365), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_36), .A2(n_43), .B1(n_357), .B2(n_396), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_37), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_38), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_39), .A2(n_166), .B1(n_364), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_40), .A2(n_241), .B1(n_391), .B2(n_445), .Y(n_882) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_42), .A2(n_95), .B1(n_295), .B2(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g820 ( .A(n_42), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_45), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_46), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_47), .A2(n_222), .B1(n_473), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_48), .A2(n_212), .B1(n_357), .B2(n_448), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_49), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_50), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_51), .A2(n_195), .B1(n_391), .B2(n_520), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_52), .A2(n_213), .B1(n_365), .B2(n_451), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_53), .A2(n_244), .B1(n_439), .B2(n_443), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_54), .A2(n_91), .B1(n_341), .B2(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_55), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_56), .A2(n_158), .B1(n_164), .B2(n_292), .C1(n_329), .C2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_57), .A2(n_105), .B1(n_347), .B2(n_349), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_58), .A2(n_80), .B1(n_398), .B2(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_59), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_60), .A2(n_229), .B1(n_306), .B2(n_311), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_61), .A2(n_235), .B1(n_355), .B2(n_358), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_62), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_63), .A2(n_178), .B1(n_383), .B2(n_384), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_64), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_65), .Y(n_509) );
INVxp67_ASAP7_75t_L g864 ( .A(n_66), .Y(n_864) );
XNOR2x1_ASAP7_75t_L g866 ( .A(n_66), .B(n_867), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_67), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_68), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_69), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_70), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_71), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_72), .A2(n_119), .B1(n_515), .B2(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_73), .A2(n_137), .B1(n_375), .B2(n_515), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_74), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_75), .A2(n_134), .B1(n_341), .B2(n_767), .Y(n_803) );
XNOR2x2_ASAP7_75t_L g658 ( .A(n_77), .B(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_78), .A2(n_202), .B1(n_796), .B2(n_798), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_79), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_81), .B(n_425), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_82), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_84), .A2(n_96), .B1(n_355), .B2(n_693), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_85), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_86), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_87), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_88), .A2(n_116), .B1(n_443), .B2(n_445), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_89), .A2(n_189), .B1(n_391), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_90), .A2(n_156), .B1(n_333), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_92), .A2(n_159), .B1(n_364), .B2(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_94), .Y(n_791) );
AND2x2_ASAP7_75t_L g277 ( .A(n_97), .B(n_278), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_98), .A2(n_193), .B1(n_622), .B2(n_696), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_100), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_102), .A2(n_616), .B1(n_652), .B2(n_653), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_102), .Y(n_652) );
INVx1_ASAP7_75t_L g274 ( .A(n_103), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_104), .A2(n_243), .B1(n_669), .B2(n_670), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_106), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_107), .A2(n_115), .B1(n_481), .B2(n_526), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_108), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_109), .A2(n_263), .B1(n_307), .B2(n_376), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_110), .A2(n_238), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_111), .A2(n_190), .B1(n_669), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_112), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_113), .A2(n_245), .B1(n_381), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_114), .A2(n_228), .B1(n_339), .B2(n_389), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_117), .A2(n_121), .B1(n_376), .B2(n_384), .Y(n_565) );
OA22x2_ASAP7_75t_L g552 ( .A1(n_118), .A2(n_553), .B1(n_554), .B2(n_574), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_118), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_120), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_122), .B(n_592), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_123), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_124), .B(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_126), .Y(n_708) );
AOI22xp5_ASAP7_75t_SL g748 ( .A1(n_128), .A2(n_749), .B1(n_750), .B2(n_772), .Y(n_748) );
INVx1_ASAP7_75t_L g772 ( .A(n_128), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_129), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_133), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_135), .A2(n_260), .B1(n_307), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_138), .A2(n_252), .B1(n_622), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_139), .A2(n_174), .B1(n_723), .B2(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_140), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_141), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_142), .B(n_379), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_143), .Y(n_713) );
XNOR2x2_ASAP7_75t_L g718 ( .A(n_144), .B(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_146), .A2(n_167), .B1(n_439), .B2(n_440), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_147), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_148), .Y(n_836) );
INVx2_ASAP7_75t_L g278 ( .A(n_149), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_150), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_151), .A2(n_176), .B1(n_607), .B2(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_152), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_154), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_155), .B(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_157), .A2(n_160), .B1(n_349), .B2(n_664), .Y(n_663) );
AOI222xp33_ASAP7_75t_L g855 ( .A1(n_161), .A2(n_221), .B1(n_250), .B2(n_419), .C1(n_425), .C2(n_736), .Y(n_855) );
AND2x6_ASAP7_75t_L g273 ( .A(n_162), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_162), .Y(n_813) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_163), .A2(n_225), .B1(n_295), .B2(n_299), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_165), .A2(n_199), .B1(n_448), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_168), .A2(n_240), .B1(n_740), .B2(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_169), .B(n_381), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_170), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_171), .Y(n_423) );
INVx1_ASAP7_75t_L g431 ( .A(n_172), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_173), .A2(n_823), .B1(n_824), .B2(n_856), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_173), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_177), .A2(n_242), .B1(n_450), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_179), .A2(n_255), .B1(n_364), .B2(n_522), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_180), .A2(n_187), .B1(n_329), .B2(n_333), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_181), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_182), .A2(n_206), .B1(n_357), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_183), .A2(n_248), .B1(n_538), .B2(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_184), .A2(n_269), .B1(n_339), .B2(n_342), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_185), .A2(n_219), .B1(n_621), .B2(n_622), .Y(n_620) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_186), .A2(n_246), .B1(n_295), .B2(n_296), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_188), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_191), .B(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_194), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_196), .A2(n_226), .B1(n_396), .B2(n_398), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_197), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_198), .A2(n_247), .B1(n_329), .B2(n_375), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_200), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_201), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_203), .A2(n_251), .B1(n_800), .B2(n_801), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_204), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_205), .A2(n_223), .B1(n_375), .B2(n_376), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_207), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_208), .A2(n_686), .B1(n_715), .B2(n_716), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_208), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_209), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_210), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_211), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_214), .Y(n_464) );
INVx1_ASAP7_75t_L g674 ( .A(n_215), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_217), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_218), .B(n_317), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_220), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_224), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_225), .B(n_818), .Y(n_817) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_227), .A2(n_271), .B(n_279), .C(n_821), .Y(n_270) );
INVx1_ASAP7_75t_L g533 ( .A(n_231), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_232), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_233), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_234), .B(n_564), .Y(n_675) );
INVx1_ASAP7_75t_L g527 ( .A(n_236), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_237), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_239), .Y(n_367) );
INVx1_ASAP7_75t_L g816 ( .A(n_246), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_249), .Y(n_841) );
OA22x2_ASAP7_75t_SL g402 ( .A1(n_253), .A2(n_403), .B1(n_404), .B2(n_452), .Y(n_402) );
INVx1_ASAP7_75t_L g452 ( .A(n_253), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_254), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_256), .Y(n_588) );
INVx1_ASAP7_75t_L g295 ( .A(n_257), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_261), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_262), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_264), .Y(n_877) );
OA22x2_ASAP7_75t_L g456 ( .A1(n_265), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_265), .Y(n_457) );
AOI22x1_ASAP7_75t_L g580 ( .A1(n_267), .A2(n_581), .B1(n_608), .B2(n_609), .Y(n_580) );
INVx1_ASAP7_75t_L g608 ( .A(n_267), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_268), .Y(n_512) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_274), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_275), .A2(n_811), .B(n_863), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_656), .B1(n_806), .B2(n_807), .C(n_808), .Y(n_279) );
INVx1_ASAP7_75t_L g806 ( .A(n_280), .Y(n_806) );
AOI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_613), .B1(n_654), .B2(n_655), .Y(n_280) );
INVx1_ASAP7_75t_L g654 ( .A(n_281), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_453), .B1(n_611), .B2(n_612), .Y(n_281) );
INVx2_ASAP7_75t_SL g611 ( .A(n_282), .Y(n_611) );
XNOR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_402), .Y(n_282) );
OAI22x1_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_368), .B2(n_401), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
XOR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_367), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_336), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_315), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_305), .Y(n_288) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g587 ( .A(n_291), .Y(n_587) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g372 ( .A(n_292), .Y(n_372) );
INVx4_ASAP7_75t_L g420 ( .A(n_292), .Y(n_420) );
BUFx3_ASAP7_75t_L g468 ( .A(n_292), .Y(n_468) );
INVx2_ASAP7_75t_L g704 ( .A(n_292), .Y(n_704) );
AND2x6_ASAP7_75t_L g292 ( .A(n_293), .B(n_300), .Y(n_292) );
AND2x4_ASAP7_75t_L g312 ( .A(n_293), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g434 ( .A(n_293), .Y(n_434) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
AND2x2_ASAP7_75t_L g310 ( .A(n_294), .B(n_302), .Y(n_310) );
INVx2_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_297), .Y(n_299) );
OR2x2_ASAP7_75t_L g322 ( .A(n_298), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_298), .B(n_323), .Y(n_327) );
INVx2_ASAP7_75t_L g332 ( .A(n_298), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
AND2x6_ASAP7_75t_L g341 ( .A(n_300), .B(n_321), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_300), .B(n_345), .Y(n_348) );
AND2x4_ASAP7_75t_L g357 ( .A(n_300), .B(n_327), .Y(n_357) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_L g320 ( .A(n_301), .B(n_304), .Y(n_320) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_314), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_302), .B(n_304), .Y(n_352) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g309 ( .A(n_304), .Y(n_309) );
INVx1_ASAP7_75t_L g314 ( .A(n_304), .Y(n_314) );
BUFx3_ASAP7_75t_L g425 ( .A(n_306), .Y(n_425) );
BUFx2_ASAP7_75t_L g646 ( .A(n_306), .Y(n_646) );
INVx2_ASAP7_75t_L g790 ( .A(n_306), .Y(n_790) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_307), .Y(n_375) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_307), .Y(n_592) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g331 ( .A(n_309), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g330 ( .A(n_310), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g333 ( .A(n_310), .B(n_334), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_310), .B(n_366), .Y(n_430) );
BUFx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_SL g376 ( .A(n_312), .Y(n_376) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_312), .Y(n_548) );
BUFx3_ASAP7_75t_L g875 ( .A(n_312), .Y(n_875) );
INVx1_ASAP7_75t_L g435 ( .A(n_313), .Y(n_435) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_324), .C(n_328), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
INVx5_ASAP7_75t_L g564 ( .A(n_318), .Y(n_564) );
INVx2_ASAP7_75t_L g744 ( .A(n_318), .Y(n_744) );
INVx4_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x6_ASAP7_75t_L g326 ( .A(n_320), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g364 ( .A(n_320), .B(n_345), .Y(n_364) );
INVx1_ASAP7_75t_L g411 ( .A(n_320), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_320), .B(n_327), .Y(n_416) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g410 ( .A(n_322), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g345 ( .A(n_323), .B(n_332), .Y(n_345) );
BUFx4f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g381 ( .A(n_326), .Y(n_381) );
INVx1_ASAP7_75t_SL g562 ( .A(n_326), .Y(n_562) );
BUFx2_ASAP7_75t_L g851 ( .A(n_326), .Y(n_851) );
AND2x2_ASAP7_75t_L g360 ( .A(n_327), .B(n_344), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g835 ( .A(n_327), .B(n_344), .Y(n_835) );
INVx1_ASAP7_75t_L g589 ( .A(n_329), .Y(n_589) );
BUFx4f_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_330), .Y(n_383) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_330), .Y(n_473) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_330), .Y(n_515) );
BUFx2_ASAP7_75t_L g707 ( .A(n_330), .Y(n_707) );
INVx1_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
BUFx3_ASAP7_75t_L g384 ( .A(n_333), .Y(n_384) );
INVx1_ASAP7_75t_L g678 ( .A(n_333), .Y(n_678) );
BUFx2_ASAP7_75t_L g759 ( .A(n_333), .Y(n_759) );
BUFx2_ASAP7_75t_L g788 ( .A(n_333), .Y(n_788) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x6_ASAP7_75t_L g399 ( .A(n_335), .B(n_352), .Y(n_399) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_353), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_346), .Y(n_337) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx5_ASAP7_75t_SL g388 ( .A(n_340), .Y(n_388) );
INVx1_ASAP7_75t_L g492 ( .A(n_340), .Y(n_492) );
INVx2_ASAP7_75t_L g662 ( .A(n_340), .Y(n_662) );
INVx11_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx11_ASAP7_75t_L g444 ( .A(n_341), .Y(n_444) );
BUFx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
BUFx3_ASAP7_75t_L g520 ( .A(n_343), .Y(n_520) );
BUFx3_ASAP7_75t_L g670 ( .A(n_343), .Y(n_670) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_344), .B(n_345), .Y(n_497) );
AND2x4_ASAP7_75t_L g350 ( .A(n_345), .B(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g439 ( .A(n_347), .Y(n_439) );
BUFx3_ASAP7_75t_L g599 ( .A(n_347), .Y(n_599) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_347), .Y(n_669) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_348), .Y(n_486) );
BUFx2_ASAP7_75t_SL g767 ( .A(n_348), .Y(n_767) );
INVx2_ASAP7_75t_L g802 ( .A(n_349), .Y(n_802) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g393 ( .A(n_350), .Y(n_393) );
BUFx3_ASAP7_75t_L g445 ( .A(n_350), .Y(n_445) );
BUFx2_ASAP7_75t_SL g489 ( .A(n_350), .Y(n_489) );
BUFx2_ASAP7_75t_L g522 ( .A(n_350), .Y(n_522) );
BUFx3_ASAP7_75t_L g634 ( .A(n_350), .Y(n_634) );
BUFx2_ASAP7_75t_SL g723 ( .A(n_350), .Y(n_723) );
AND2x2_ASAP7_75t_L g365 ( .A(n_351), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_361), .Y(n_353) );
INVxp67_ASAP7_75t_L g842 ( .A(n_355), .Y(n_842) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g572 ( .A(n_356), .Y(n_572) );
INVx2_ASAP7_75t_L g626 ( .A(n_356), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_356), .A2(n_495), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g770 ( .A(n_356), .Y(n_770) );
INVx6_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g542 ( .A(n_357), .Y(n_542) );
BUFx3_ASAP7_75t_L g605 ( .A(n_357), .Y(n_605) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx4_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
INVx5_ASAP7_75t_L g451 ( .A(n_359), .Y(n_451) );
INVx1_ASAP7_75t_L g479 ( .A(n_359), .Y(n_479) );
INVx2_ASAP7_75t_L g672 ( .A(n_359), .Y(n_672) );
INVx8_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g441 ( .A(n_364), .Y(n_441) );
BUFx3_ASAP7_75t_L g526 ( .A(n_364), .Y(n_526) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_364), .Y(n_666) );
BUFx3_ASAP7_75t_L g886 ( .A(n_364), .Y(n_886) );
INVx3_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
XOR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_400), .Y(n_368) );
NAND2x1_ASAP7_75t_SL g369 ( .A(n_370), .B(n_385), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_377), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B(n_374), .Y(n_371) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_372), .A2(n_734), .B(n_735), .Y(n_733) );
INVx2_ASAP7_75t_L g756 ( .A(n_375), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .C(n_382), .Y(n_377) );
INVx2_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
INVx4_ASAP7_75t_L g737 ( .A(n_383), .Y(n_737) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_394), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g727 ( .A(n_388), .Y(n_727) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_388), .Y(n_847) );
BUFx3_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g537 ( .A(n_392), .Y(n_537) );
BUFx2_ASAP7_75t_L g602 ( .A(n_393), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_396), .Y(n_696) );
INVx2_ASAP7_75t_L g797 ( .A(n_396), .Y(n_797) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx6_ASAP7_75t_SL g482 ( .A(n_399), .Y(n_482) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_SL g404 ( .A(n_405), .B(n_436), .Y(n_404) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_417), .C(n_426), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_412), .B2(n_413), .Y(n_406) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g462 ( .A(n_409), .Y(n_462) );
INVx1_ASAP7_75t_SL g712 ( .A(n_409), .Y(n_712) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g504 ( .A(n_410), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_410), .A2(n_415), .B1(n_545), .B2(n_546), .C(n_547), .Y(n_544) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_410), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_410), .A2(n_506), .B1(n_870), .B2(n_871), .Y(n_869) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_413), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g714 ( .A(n_415), .Y(n_714) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g507 ( .A(n_416), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B1(n_422), .B2(n_423), .C(n_424), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_418), .A2(n_642), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g752 ( .A1(n_418), .A2(n_753), .B(n_754), .Y(n_752) );
OAI21xp33_ASAP7_75t_SL g785 ( .A1(n_418), .A2(n_786), .B(n_787), .Y(n_785) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g508 ( .A1(n_420), .A2(n_509), .B(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_431), .B2(n_432), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_428), .A2(n_706), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_SL g700 ( .A(n_429), .Y(n_700) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_430), .A2(n_512), .B1(n_513), .B2(n_516), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_430), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_430), .A2(n_433), .B1(n_853), .B2(n_854), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_432), .A2(n_475), .B1(n_594), .B2(n_595), .Y(n_593) );
OAI22xp5_ASAP7_75t_SL g789 ( .A1(n_432), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_789) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g640 ( .A(n_433), .Y(n_640) );
OR2x6_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_446), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_442), .Y(n_437) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g631 ( .A(n_441), .Y(n_631) );
INVx4_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx4_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
INVx2_ASAP7_75t_SL g600 ( .A(n_444), .Y(n_600) );
INVx3_ASAP7_75t_L g764 ( .A(n_444), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g612 ( .A(n_453), .Y(n_612) );
XOR2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_529), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_498), .B1(n_499), .B2(n_528), .Y(n_455) );
INVx2_ASAP7_75t_L g528 ( .A(n_456), .Y(n_528) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_476), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .C(n_470), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_462), .A2(n_506), .B1(n_584), .B2(n_585), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_469), .Y(n_465) );
OAI21xp5_ASAP7_75t_SL g549 ( .A1(n_467), .A2(n_550), .B(n_551), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g556 ( .A1(n_467), .A2(n_557), .B(n_558), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_467), .A2(n_873), .B(n_874), .Y(n_872) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_474), .B2(n_475), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_483), .C(n_490), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_479), .Y(n_621) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx4f_ASAP7_75t_SL g607 ( .A(n_482), .Y(n_607) );
BUFx2_ASAP7_75t_L g622 ( .A(n_482), .Y(n_622) );
BUFx2_ASAP7_75t_L g798 ( .A(n_482), .Y(n_798) );
BUFx2_ASAP7_75t_L g838 ( .A(n_482), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_487), .B2(n_488), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g628 ( .A(n_496), .Y(n_628) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
XOR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_527), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_517), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .C(n_511), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_502) );
OA211x2_ASAP7_75t_L g673 ( .A1(n_506), .A2(n_674), .B(n_675), .C(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g651 ( .A(n_507), .Y(n_651) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g643 ( .A(n_514), .Y(n_643) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
INVx1_ASAP7_75t_L g694 ( .A(n_520), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_577), .B1(n_578), .B2(n_610), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g610 ( .A(n_531), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_552), .B1(n_575), .B2(n_576), .Y(n_531) );
INVx2_ASAP7_75t_SL g575 ( .A(n_532), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_532), .A2(n_575), .B1(n_579), .B2(n_580), .Y(n_578) );
XNOR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NOR4xp75_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .C(n_544), .D(n_549), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_539), .Y(n_535) );
INVxp67_ASAP7_75t_L g830 ( .A(n_537), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_SL g742 ( .A(n_548), .Y(n_742) );
INVx1_ASAP7_75t_L g576 ( .A(n_552), .Y(n_576) );
INVx1_ASAP7_75t_L g574 ( .A(n_554), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_566), .Y(n_554) );
NOR2xp67_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .C(n_565), .Y(n_559) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_564), .Y(n_850) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g609 ( .A(n_581), .Y(n_609) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_596), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .C(n_593), .Y(n_582) );
OAI221xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_590), .C(n_591), .Y(n_586) );
BUFx4f_ASAP7_75t_L g680 ( .A(n_592), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g655 ( .A(n_613), .Y(n_655) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g653 ( .A(n_616), .Y(n_653) );
AND2x2_ASAP7_75t_SL g616 ( .A(n_617), .B(n_635), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_623), .C(n_629), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_623) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_628), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_631), .A2(n_845), .B1(n_846), .B2(n_848), .Y(n_844) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_641), .C(n_647), .Y(n_635) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g702 ( .A(n_640), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_647) );
INVx1_ASAP7_75t_L g783 ( .A(n_649), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_651), .A2(n_781), .B1(n_782), .B2(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g807 ( .A(n_656), .Y(n_807) );
AOI22xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_775), .B1(n_804), .B2(n_805), .Y(n_656) );
INVx1_ASAP7_75t_L g804 ( .A(n_657), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_681), .B1(n_773), .B2(n_774), .Y(n_657) );
INVx1_ASAP7_75t_L g773 ( .A(n_658), .Y(n_773) );
NAND4xp75_ASAP7_75t_L g659 ( .A(n_660), .B(n_667), .C(n_673), .D(n_679), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_665), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
INVx4_ASAP7_75t_L g800 ( .A(n_665), .Y(n_800) );
INVx4_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
BUFx4f_ASAP7_75t_SL g765 ( .A(n_670), .Y(n_765) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g740 ( .A(n_678), .Y(n_740) );
INVx1_ASAP7_75t_L g774 ( .A(n_681), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_745), .B2(n_746), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_717), .B2(n_718), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g716 ( .A(n_686), .Y(n_716) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_687), .B(n_697), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR3xp33_ASAP7_75t_SL g697 ( .A(n_698), .B(n_703), .C(n_710), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_708), .C(n_709), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_720), .B(n_732), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_725), .C(n_729), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_738), .Y(n_732) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_761), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_757), .Y(n_751) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_768), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g805 ( .A(n_775), .Y(n_805) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
XNOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_793), .Y(n_778) );
NOR3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_785), .C(n_789), .Y(n_779) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND4x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .C(n_799), .D(n_803), .Y(n_793) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_802), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_828) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
NOR2x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
OR2x2_ASAP7_75t_SL g889 ( .A(n_810), .B(n_815), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_812), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_812), .B(n_860), .Y(n_863) );
CKINVDCx16_ASAP7_75t_R g860 ( .A(n_813), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
OAI322xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_857), .A3(n_858), .B1(n_861), .B2(n_864), .C1(n_865), .C2(n_887), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND4x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_839), .C(n_849), .D(n_855), .Y(n_826) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_828), .B(n_832), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_836), .B2(n_837), .Y(n_832) );
BUFx2_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
INVxp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_879), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .C(n_876), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
endmodule