module real_aes_16875_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1121 ( .A1(n_0), .A2(n_3), .B1(n_864), .B2(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1158 ( .A1(n_0), .A2(n_240), .B1(n_1159), .B2(n_1160), .Y(n_1158) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1), .Y(n_1039) );
INVx1_ASAP7_75t_L g439 ( .A(n_2), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_3), .A2(n_241), .B1(n_830), .B2(n_1159), .Y(n_1163) );
XNOR2xp5_ASAP7_75t_L g758 ( .A(n_4), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g949 ( .A(n_5), .Y(n_949) );
OAI211xp5_ASAP7_75t_L g881 ( .A1(n_6), .A2(n_569), .B(n_624), .C(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g893 ( .A(n_6), .Y(n_893) );
INVx1_ASAP7_75t_L g295 ( .A(n_7), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_7), .B(n_305), .Y(n_459) );
INVx1_ASAP7_75t_L g1137 ( .A(n_8), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_8), .A2(n_28), .B1(n_1149), .B2(n_1150), .Y(n_1148) );
INVx1_ASAP7_75t_L g898 ( .A(n_9), .Y(n_898) );
INVx1_ASAP7_75t_L g841 ( .A(n_10), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_11), .A2(n_181), .B1(n_297), .B2(n_407), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1062 ( .A1(n_11), .A2(n_181), .B1(n_315), .B2(n_324), .Y(n_1062) );
OAI211xp5_ASAP7_75t_L g1074 ( .A1(n_12), .A2(n_643), .B(n_1075), .C(n_1077), .Y(n_1074) );
INVx1_ASAP7_75t_L g1085 ( .A(n_12), .Y(n_1085) );
INVx1_ASAP7_75t_L g1143 ( .A(n_13), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_14), .B(n_1176), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_14), .B(n_102), .Y(n_1178) );
INVx2_ASAP7_75t_L g1182 ( .A(n_14), .Y(n_1182) );
OAI22xp33_ASAP7_75t_SL g1032 ( .A1(n_15), .A2(n_17), .B1(n_563), .B2(n_935), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_15), .A2(n_17), .B1(n_357), .B2(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1396 ( .A(n_16), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g1461 ( .A1(n_18), .A2(n_127), .B1(n_1418), .B2(n_1462), .Y(n_1461) );
OAI22xp33_ASAP7_75t_L g1470 ( .A1(n_18), .A2(n_127), .B1(n_297), .B2(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1093 ( .A(n_19), .Y(n_1093) );
INVx1_ASAP7_75t_L g1050 ( .A(n_20), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_21), .A2(n_214), .B1(n_551), .B2(n_1005), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_21), .A2(n_233), .B1(n_517), .B2(n_1018), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_22), .A2(n_156), .B1(n_407), .B2(n_684), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_22), .A2(n_269), .B1(n_317), .B2(n_640), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g1186 ( .A1(n_23), .A2(n_185), .B1(n_1183), .B2(n_1187), .Y(n_1186) );
XNOR2xp5_ASAP7_75t_L g1384 ( .A(n_23), .B(n_1385), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_23), .A2(n_1431), .B1(n_1433), .B2(n_1477), .Y(n_1430) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_24), .A2(n_172), .B1(n_1177), .B2(n_1183), .Y(n_1193) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_25), .Y(n_660) );
XNOR2x2_ASAP7_75t_SL g1070 ( .A(n_26), .B(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_26), .A2(n_205), .B1(n_1173), .B2(n_1180), .Y(n_1227) );
INVx1_ASAP7_75t_L g958 ( .A(n_27), .Y(n_958) );
INVx1_ASAP7_75t_L g1140 ( .A(n_28), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_29), .A2(n_207), .B1(n_401), .B2(n_634), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_29), .A2(n_96), .B1(n_317), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g1079 ( .A(n_30), .Y(n_1079) );
OAI211xp5_ASAP7_75t_L g1083 ( .A1(n_30), .A2(n_751), .B(n_905), .C(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g957 ( .A(n_31), .Y(n_957) );
INVx1_ASAP7_75t_L g423 ( .A(n_32), .Y(n_423) );
INVx1_ASAP7_75t_L g710 ( .A(n_33), .Y(n_710) );
INVx1_ASAP7_75t_L g778 ( .A(n_34), .Y(n_778) );
INVx1_ASAP7_75t_L g1144 ( .A(n_35), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_36), .Y(n_666) );
INVx1_ASAP7_75t_L g1443 ( .A(n_37), .Y(n_1443) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_38), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g880 ( .A1(n_39), .A2(n_120), .B1(n_684), .B2(n_851), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_39), .A2(n_52), .B1(n_359), .B2(n_640), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_40), .A2(n_213), .B1(n_1173), .B2(n_1183), .Y(n_1200) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_41), .A2(n_97), .B1(n_1173), .B2(n_1180), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_42), .A2(n_159), .B1(n_407), .B2(n_634), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_42), .A2(n_115), .B1(n_317), .B2(n_355), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_43), .A2(n_277), .B1(n_317), .B2(n_356), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_43), .A2(n_45), .B1(n_684), .B2(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g766 ( .A(n_44), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_45), .A2(n_175), .B1(n_359), .B2(n_640), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_46), .A2(n_106), .B1(n_1173), .B2(n_1180), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_47), .A2(n_80), .B1(n_1005), .B2(n_1007), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_47), .A2(n_88), .B1(n_595), .B2(n_1016), .Y(n_1019) );
INVx1_ASAP7_75t_L g803 ( .A(n_48), .Y(n_803) );
OAI211xp5_ASAP7_75t_L g809 ( .A1(n_48), .A2(n_643), .B(n_810), .C(n_811), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_49), .A2(n_133), .B1(n_315), .B2(n_324), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_49), .A2(n_133), .B1(n_297), .B2(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g321 ( .A(n_50), .Y(n_321) );
INVx1_ASAP7_75t_L g337 ( .A(n_50), .Y(n_337) );
INVx1_ASAP7_75t_L g988 ( .A(n_51), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_51), .A2(n_100), .B1(n_603), .B2(n_997), .C(n_998), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_52), .A2(n_211), .B1(n_634), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_53), .A2(n_73), .B1(n_864), .B2(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1157 ( .A(n_53), .Y(n_1157) );
INVx1_ASAP7_75t_L g1398 ( .A(n_54), .Y(n_1398) );
INVx1_ASAP7_75t_L g783 ( .A(n_55), .Y(n_783) );
INVx1_ASAP7_75t_L g741 ( .A(n_56), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g754 ( .A1(n_56), .A2(n_158), .B1(n_407), .B2(n_634), .Y(n_754) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_57), .A2(n_478), .B(n_624), .C(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g647 ( .A(n_57), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_58), .A2(n_204), .B1(n_511), .B2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_58), .A2(n_212), .B1(n_547), .B2(n_551), .Y(n_554) );
INVx1_ASAP7_75t_L g288 ( .A(n_59), .Y(n_288) );
INVx2_ASAP7_75t_L g323 ( .A(n_60), .Y(n_323) );
INVx1_ASAP7_75t_L g1052 ( .A(n_61), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_62), .A2(n_244), .B1(n_736), .B2(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_62), .A2(n_177), .B1(n_866), .B2(n_868), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_63), .A2(n_85), .B1(n_1180), .B2(n_1187), .Y(n_1201) );
INVx1_ASAP7_75t_L g840 ( .A(n_64), .Y(n_840) );
INVx1_ASAP7_75t_L g884 ( .A(n_65), .Y(n_884) );
INVx1_ASAP7_75t_L g706 ( .A(n_66), .Y(n_706) );
INVx1_ASAP7_75t_L g838 ( .A(n_67), .Y(n_838) );
INVx1_ASAP7_75t_L g1100 ( .A(n_68), .Y(n_1100) );
OAI222xp33_ASAP7_75t_L g499 ( .A1(n_69), .A2(n_105), .B1(n_238), .B2(n_500), .C1(n_502), .C2(n_503), .Y(n_499) );
OAI222xp33_ASAP7_75t_L g566 ( .A1(n_69), .A2(n_105), .B1(n_238), .B2(n_389), .C1(n_567), .C2(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g901 ( .A(n_70), .Y(n_901) );
INVx1_ASAP7_75t_L g1133 ( .A(n_71), .Y(n_1133) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_72), .A2(n_96), .B1(n_396), .B2(n_407), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_72), .A2(n_207), .B1(n_356), .B2(n_359), .Y(n_648) );
INVxp67_ASAP7_75t_SL g1162 ( .A(n_73), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g1463 ( .A1(n_74), .A2(n_339), .B(n_1464), .C(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1474 ( .A(n_74), .Y(n_1474) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_75), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_76), .A2(n_278), .B1(n_520), .B2(n_523), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_76), .A2(n_132), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_77), .A2(n_132), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_77), .A2(n_278), .B1(n_547), .B2(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g952 ( .A(n_78), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_79), .A2(n_276), .B1(n_532), .B2(n_825), .C(n_826), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_79), .A2(n_130), .B1(n_557), .B2(n_871), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_80), .A2(n_191), .B1(n_1014), .B2(n_1016), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1197 ( .A1(n_81), .A2(n_123), .B1(n_1173), .B2(n_1180), .Y(n_1197) );
INVx1_ASAP7_75t_L g1453 ( .A(n_82), .Y(n_1453) );
OAI211xp5_ASAP7_75t_L g1411 ( .A1(n_83), .A2(n_1027), .B(n_1028), .C(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1422 ( .A(n_83), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_84), .A2(n_174), .B1(n_563), .B2(n_748), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_84), .A2(n_174), .B1(n_939), .B2(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1138 ( .A(n_86), .Y(n_1138) );
INVx1_ASAP7_75t_L g711 ( .A(n_87), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_88), .A2(n_191), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_89), .Y(n_802) );
INVx1_ASAP7_75t_L g577 ( .A(n_90), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g1205 ( .A1(n_90), .A2(n_121), .B1(n_1173), .B2(n_1180), .Y(n_1205) );
INVx1_ASAP7_75t_L g1441 ( .A(n_91), .Y(n_1441) );
INVx1_ASAP7_75t_L g431 ( .A(n_92), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_93), .A2(n_216), .B1(n_684), .B2(n_851), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_93), .A2(n_216), .B1(n_356), .B2(n_359), .Y(n_999) );
AOI22xp5_ASAP7_75t_SL g1204 ( .A1(n_94), .A2(n_260), .B1(n_1183), .B2(n_1187), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_95), .Y(n_290) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_95), .B(n_288), .Y(n_1174) );
INVx1_ASAP7_75t_L g1099 ( .A(n_98), .Y(n_1099) );
INVx1_ASAP7_75t_L g1030 ( .A(n_99), .Y(n_1030) );
INVx1_ASAP7_75t_L g991 ( .A(n_100), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g1215 ( .A1(n_101), .A2(n_108), .B1(n_1177), .B2(n_1183), .Y(n_1215) );
INVx1_ASAP7_75t_L g1176 ( .A(n_102), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_102), .B(n_1182), .Y(n_1184) );
INVx1_ASAP7_75t_L g777 ( .A(n_103), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_104), .A2(n_273), .B1(n_1173), .B2(n_1177), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_107), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_109), .A2(n_228), .B1(n_496), .B2(n_497), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_109), .A2(n_228), .B1(n_563), .B2(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g366 ( .A(n_110), .Y(n_366) );
INVx1_ASAP7_75t_L g447 ( .A(n_110), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_111), .Y(n_585) );
INVx1_ASAP7_75t_L g904 ( .A(n_112), .Y(n_904) );
INVx1_ASAP7_75t_L g1095 ( .A(n_113), .Y(n_1095) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_114), .A2(n_236), .B1(n_1173), .B2(n_1180), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_115), .A2(n_122), .B1(n_563), .B2(n_805), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_116), .Y(n_590) );
XNOR2xp5_ASAP7_75t_L g1022 ( .A(n_117), .B(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1413 ( .A(n_118), .Y(n_1413) );
INVx1_ASAP7_75t_L g491 ( .A(n_119), .Y(n_491) );
OAI22xp5_ASAP7_75t_SL g888 ( .A1(n_120), .A2(n_211), .B1(n_317), .B2(n_356), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_122), .A2(n_159), .B1(n_324), .B2(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g453 ( .A(n_124), .Y(n_453) );
INVx1_ASAP7_75t_L g908 ( .A(n_125), .Y(n_908) );
INVx1_ASAP7_75t_L g1389 ( .A(n_126), .Y(n_1389) );
INVx1_ASAP7_75t_L g714 ( .A(n_128), .Y(n_714) );
INVx1_ASAP7_75t_L g1450 ( .A(n_129), .Y(n_1450) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_130), .A2(n_219), .B1(n_532), .B2(n_825), .C(n_828), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_131), .A2(n_235), .B1(n_317), .B2(n_1081), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_131), .A2(n_235), .B1(n_407), .B2(n_634), .Y(n_1088) );
XOR2xp5_ASAP7_75t_L g487 ( .A(n_134), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g1390 ( .A(n_135), .Y(n_1390) );
INVx1_ASAP7_75t_L g1394 ( .A(n_136), .Y(n_1394) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_137), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_138), .A2(n_250), .B1(n_1183), .B2(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1106 ( .A(n_139), .Y(n_1106) );
INVx1_ASAP7_75t_L g906 ( .A(n_140), .Y(n_906) );
AOI31xp33_ASAP7_75t_L g819 ( .A1(n_141), .A2(n_820), .A3(n_834), .B(n_844), .Y(n_819) );
NAND2xp33_ASAP7_75t_SL g861 ( .A(n_141), .B(n_862), .Y(n_861) );
INVxp67_ASAP7_75t_SL g875 ( .A(n_141), .Y(n_875) );
INVx1_ASAP7_75t_L g982 ( .A(n_142), .Y(n_982) );
INVx1_ASAP7_75t_L g1044 ( .A(n_143), .Y(n_1044) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_144), .A2(n_247), .B1(n_297), .B2(n_886), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_144), .A2(n_247), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
INVx1_ASAP7_75t_L g739 ( .A(n_145), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_145), .A2(n_257), .B1(n_563), .B2(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g734 ( .A(n_146), .Y(n_734) );
OA211x2_ASAP7_75t_L g750 ( .A1(n_146), .A2(n_569), .B(n_751), .C(n_752), .Y(n_750) );
BUFx3_ASAP7_75t_L g319 ( .A(n_147), .Y(n_319) );
INVx1_ASAP7_75t_L g1120 ( .A(n_148), .Y(n_1120) );
INVx1_ASAP7_75t_L g899 ( .A(n_149), .Y(n_899) );
INVx1_ASAP7_75t_L g421 ( .A(n_150), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_151), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_152), .Y(n_667) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_153), .A2(n_695), .B1(n_745), .B2(n_756), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_153), .B(n_696), .C(n_716), .D(n_728), .Y(n_695) );
INVx1_ASAP7_75t_L g1467 ( .A(n_154), .Y(n_1467) );
OAI211xp5_ASAP7_75t_L g1472 ( .A1(n_154), .A2(n_379), .B(n_928), .C(n_1473), .Y(n_1472) );
XOR2xp5_ASAP7_75t_L g1434 ( .A(n_155), .B(n_1435), .Y(n_1434) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_156), .A2(n_274), .B1(n_356), .B2(n_359), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_157), .Y(n_664) );
INVx1_ASAP7_75t_L g738 ( .A(n_158), .Y(n_738) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_160), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_161), .A2(n_212), .B1(n_511), .B2(n_517), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_204), .B1(n_539), .B2(n_543), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_162), .Y(n_655) );
INVx1_ASAP7_75t_L g781 ( .A(n_163), .Y(n_781) );
INVx1_ASAP7_75t_L g1047 ( .A(n_164), .Y(n_1047) );
XOR2x2_ASAP7_75t_L g877 ( .A(n_165), .B(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g427 ( .A(n_166), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g799 ( .A1(n_167), .A2(n_751), .B(n_800), .C(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g812 ( .A(n_167), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_168), .A2(n_199), .B1(n_297), .B2(n_407), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g945 ( .A1(n_168), .A2(n_199), .B1(n_315), .B2(n_324), .Y(n_945) );
INVx1_ASAP7_75t_L g349 ( .A(n_169), .Y(n_349) );
INVx1_ASAP7_75t_L g832 ( .A(n_170), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_170), .A2(n_244), .B1(n_544), .B2(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g1103 ( .A(n_171), .Y(n_1103) );
INVx1_ASAP7_75t_L g1107 ( .A(n_173), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_175), .Y(n_848) );
INVx1_ASAP7_75t_L g1134 ( .A(n_176), .Y(n_1134) );
INVx1_ASAP7_75t_L g831 ( .A(n_177), .Y(n_831) );
INVx1_ASAP7_75t_L g768 ( .A(n_178), .Y(n_768) );
INVx1_ASAP7_75t_L g701 ( .A(n_179), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g924 ( .A(n_180), .B(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g1036 ( .A(n_182), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_183), .A2(n_201), .B1(n_356), .B2(n_357), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_183), .A2(n_201), .B1(n_396), .B2(n_805), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_184), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_186), .A2(n_192), .B1(n_1177), .B2(n_1183), .Y(n_1226) );
INVx1_ASAP7_75t_L g909 ( .A(n_187), .Y(n_909) );
OAI211xp5_ASAP7_75t_SL g927 ( .A1(n_188), .A2(n_751), .B(n_928), .C(n_930), .Y(n_927) );
INVx1_ASAP7_75t_L g944 ( .A(n_188), .Y(n_944) );
INVx1_ASAP7_75t_L g950 ( .A(n_189), .Y(n_950) );
OAI211xp5_ASAP7_75t_SL g331 ( .A1(n_190), .A2(n_332), .B(n_339), .C(n_343), .Y(n_331) );
INVx1_ASAP7_75t_L g393 ( .A(n_190), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_193), .Y(n_659) );
INVx1_ASAP7_75t_L g703 ( .A(n_194), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_195), .Y(n_588) );
INVx1_ASAP7_75t_L g1414 ( .A(n_196), .Y(n_1414) );
OAI211xp5_ASAP7_75t_L g1420 ( .A1(n_196), .A2(n_332), .B(n_339), .C(n_1421), .Y(n_1420) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_197), .A2(n_263), .B1(n_355), .B2(n_357), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_197), .A2(n_263), .B1(n_395), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_L g700 ( .A(n_198), .Y(n_700) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
INVx1_ASAP7_75t_L g1448 ( .A(n_202), .Y(n_1448) );
INVx1_ASAP7_75t_L g1452 ( .A(n_203), .Y(n_1452) );
INVx1_ASAP7_75t_L g1401 ( .A(n_206), .Y(n_1401) );
INVx1_ASAP7_75t_L g681 ( .A(n_208), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_208), .A2(n_450), .B(n_643), .C(n_688), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_209), .Y(n_583) );
INVx1_ASAP7_75t_L g883 ( .A(n_210), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1020 ( .A1(n_214), .A2(n_261), .B1(n_826), .B2(n_830), .C(n_1018), .Y(n_1020) );
INVx1_ASAP7_75t_L g1104 ( .A(n_215), .Y(n_1104) );
INVx1_ASAP7_75t_L g902 ( .A(n_217), .Y(n_902) );
INVx1_ASAP7_75t_L g932 ( .A(n_218), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_219), .A2(n_276), .B1(n_866), .B2(n_868), .Y(n_865) );
INVx1_ASAP7_75t_L g1031 ( .A(n_220), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1063 ( .A1(n_220), .A2(n_332), .B(n_339), .C(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1444 ( .A(n_221), .Y(n_1444) );
INVx1_ASAP7_75t_L g983 ( .A(n_222), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_223), .Y(n_629) );
INVx1_ASAP7_75t_L g954 ( .A(n_224), .Y(n_954) );
INVx1_ASAP7_75t_L g1393 ( .A(n_225), .Y(n_1393) );
BUFx3_ASAP7_75t_L g305 ( .A(n_226), .Y(n_305) );
INVx1_ASAP7_75t_L g398 ( .A(n_226), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_227), .A2(n_265), .B1(n_563), .B2(n_935), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_227), .A2(n_265), .B1(n_939), .B2(n_940), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_229), .A2(n_259), .B1(n_355), .B2(n_1424), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_229), .A2(n_259), .B1(n_563), .B2(n_1476), .Y(n_1475) );
XOR2x2_ASAP7_75t_L g311 ( .A(n_230), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g733 ( .A(n_231), .Y(n_733) );
INVx1_ASAP7_75t_L g715 ( .A(n_232), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_233), .A2(n_261), .B1(n_556), .B2(n_557), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_234), .A2(n_478), .B(n_624), .C(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g689 ( .A(n_234), .Y(n_689) );
INVx1_ASAP7_75t_L g441 ( .A(n_237), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_239), .Y(n_596) );
INVxp67_ASAP7_75t_SL g1124 ( .A(n_240), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_241), .Y(n_1125) );
INVx1_ASAP7_75t_L g371 ( .A(n_242), .Y(n_371) );
INVx1_ASAP7_75t_L g446 ( .A(n_242), .Y(n_446) );
INVx2_ASAP7_75t_L g458 ( .A(n_242), .Y(n_458) );
INVx1_ASAP7_75t_L g763 ( .A(n_243), .Y(n_763) );
INVx1_ASAP7_75t_L g1078 ( .A(n_245), .Y(n_1078) );
INVx1_ASAP7_75t_L g1119 ( .A(n_246), .Y(n_1119) );
INVx1_ASAP7_75t_L g1466 ( .A(n_248), .Y(n_1466) );
XNOR2xp5_ASAP7_75t_L g978 ( .A(n_249), .B(n_979), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_249), .A2(n_251), .B1(n_1180), .B2(n_1183), .Y(n_1179) );
XNOR2xp5_ASAP7_75t_L g1115 ( .A(n_252), .B(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g933 ( .A(n_253), .Y(n_933) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_253), .A2(n_332), .B(n_339), .C(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g1041 ( .A(n_254), .Y(n_1041) );
INVx1_ASAP7_75t_L g772 ( .A(n_255), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_256), .Y(n_987) );
INVx1_ASAP7_75t_L g743 ( .A(n_257), .Y(n_743) );
INVx1_ASAP7_75t_L g1400 ( .A(n_258), .Y(n_1400) );
INVx1_ASAP7_75t_L g1440 ( .A(n_262), .Y(n_1440) );
INVx1_ASAP7_75t_L g449 ( .A(n_264), .Y(n_449) );
INVx1_ASAP7_75t_L g735 ( .A(n_266), .Y(n_735) );
XNOR2xp5_ASAP7_75t_L g650 ( .A(n_267), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_268), .A2(n_374), .B(n_379), .C(n_384), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_269), .A2(n_274), .B1(n_401), .B2(n_634), .Y(n_682) );
INVx1_ASAP7_75t_L g493 ( .A(n_270), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_271), .Y(n_604) );
INVx1_ASAP7_75t_L g962 ( .A(n_272), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g1026 ( .A1(n_275), .A2(n_1027), .B(n_1028), .C(n_1029), .Y(n_1026) );
INVx1_ASAP7_75t_L g1065 ( .A(n_275), .Y(n_1065) );
INVx1_ASAP7_75t_L g846 ( .A(n_277), .Y(n_846) );
INVx1_ASAP7_75t_L g632 ( .A(n_279), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_279), .A2(n_450), .B(n_643), .C(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g1042 ( .A(n_280), .Y(n_1042) );
AOI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_306), .B(n_1167), .Y(n_281) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_285), .B(n_294), .Y(n_1429) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1432 ( .A(n_287), .B(n_290), .Y(n_1432) );
INVx1_ASAP7_75t_L g1478 ( .A(n_287), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_290), .B(n_1478), .Y(n_1480) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g412 ( .A(n_294), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g481 ( .A(n_295), .B(n_305), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_296), .A2(n_408), .B1(n_491), .B2(n_493), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_296), .A2(n_408), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
AND2x4_ASAP7_75t_SL g1428 ( .A(n_296), .B(n_1429), .Y(n_1428) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
OR2x6_ASAP7_75t_L g396 ( .A(n_298), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g684 ( .A(n_298), .B(n_397), .Y(n_684) );
BUFx4f_ASAP7_75t_L g722 ( .A(n_298), .Y(n_722) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_299), .Y(n_464) );
INVx3_ASAP7_75t_L g635 ( .A(n_299), .Y(n_635) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_301), .B(n_302), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_301), .B(n_302), .Y(n_383) );
INVx1_ASAP7_75t_L g392 ( .A(n_301), .Y(n_392) );
INVx2_ASAP7_75t_L g405 ( .A(n_301), .Y(n_405) );
AND2x2_ASAP7_75t_L g409 ( .A(n_301), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g473 ( .A(n_301), .Y(n_473) );
BUFx2_ASAP7_75t_L g387 ( .A(n_302), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_302), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g410 ( .A(n_302), .Y(n_410) );
OR2x2_ASAP7_75t_L g472 ( .A(n_302), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g542 ( .A(n_302), .Y(n_542) );
AND2x2_ASAP7_75t_L g545 ( .A(n_302), .B(n_405), .Y(n_545) );
OR2x6_ASAP7_75t_L g634 ( .A(n_303), .B(n_635), .Y(n_634) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g381 ( .A(n_304), .Y(n_381) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g386 ( .A(n_305), .Y(n_386) );
AND2x4_ASAP7_75t_L g390 ( .A(n_305), .B(n_391), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_918), .B2(n_919), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
XNOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_572), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_485), .B2(n_486), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_372), .C(n_415), .Y(n_312) );
OAI31xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_331), .A3(n_354), .B(n_362), .Y(n_313) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_316), .A2(n_325), .B1(n_1143), .B2(n_1144), .Y(n_1151) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g492 ( .A(n_317), .Y(n_492) );
INVx1_ASAP7_75t_L g742 ( .A(n_317), .Y(n_742) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_317), .Y(n_1418) );
OR2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
OR2x4_ASAP7_75t_L g356 ( .A(n_318), .B(n_326), .Y(n_356) );
BUFx3_ASAP7_75t_L g422 ( .A(n_318), .Y(n_422) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_318), .Y(n_584) );
INVx2_ASAP7_75t_L g601 ( .A(n_318), .Y(n_601) );
BUFx3_ASAP7_75t_L g789 ( .A(n_318), .Y(n_789) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g330 ( .A(n_319), .Y(n_330) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_319), .Y(n_338) );
AND2x4_ASAP7_75t_L g341 ( .A(n_319), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_319), .B(n_337), .Y(n_361) );
INVx1_ASAP7_75t_L g516 ( .A(n_320), .Y(n_516) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g329 ( .A(n_321), .Y(n_329) );
INVx1_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
AND2x4_ASAP7_75t_L g340 ( .A(n_322), .B(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g359 ( .A(n_322), .B(n_360), .Y(n_359) );
NAND3x1_ASAP7_75t_L g444 ( .A(n_322), .B(n_445), .C(n_447), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_322), .B(n_447), .Y(n_606) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
NAND2xp33_ASAP7_75t_SL g419 ( .A(n_323), .B(n_366), .Y(n_419) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_325), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_490) );
INVx2_ASAP7_75t_L g1081 ( .A(n_325), .Y(n_1081) );
INVx1_ASAP7_75t_L g1419 ( .A(n_325), .Y(n_1419) );
INVx1_ASAP7_75t_L g1462 ( .A(n_325), .Y(n_1462) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g641 ( .A(n_326), .B(n_327), .Y(n_641) );
INVx2_ASAP7_75t_L g589 ( .A(n_327), .Y(n_589) );
INVx2_ASAP7_75t_L g794 ( .A(n_327), .Y(n_794) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_327), .Y(n_825) );
INVx2_ASAP7_75t_L g1156 ( .A(n_327), .Y(n_1156) );
INVx1_ASAP7_75t_L g1449 ( .A(n_327), .Y(n_1449) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_328), .Y(n_430) );
INVx2_ASAP7_75t_L g522 ( .A(n_328), .Y(n_522) );
BUFx8_ASAP7_75t_L g709 ( .A(n_328), .Y(n_709) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g515 ( .A(n_330), .B(n_516), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_332), .A2(n_950), .B1(n_958), .B2(n_973), .Y(n_972) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g502 ( .A(n_333), .Y(n_502) );
INVx1_ASAP7_75t_L g790 ( .A(n_333), .Y(n_790) );
INVx1_ASAP7_75t_L g810 ( .A(n_333), .Y(n_810) );
INVx1_ASAP7_75t_L g916 ( .A(n_333), .Y(n_916) );
INVx4_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_334), .Y(n_670) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g452 ( .A(n_335), .Y(n_452) );
BUFx3_ASAP7_75t_L g603 ( .A(n_335), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
BUFx2_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g342 ( .A(n_337), .Y(n_342) );
BUFx2_ASAP7_75t_L g348 ( .A(n_338), .Y(n_348) );
AND2x4_ASAP7_75t_L g525 ( .A(n_338), .B(n_526), .Y(n_525) );
CKINVDCx8_ASAP7_75t_R g339 ( .A(n_340), .Y(n_339) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_340), .B(n_495), .C(n_499), .Y(n_494) );
CKINVDCx8_ASAP7_75t_R g643 ( .A(n_340), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_340), .B(n_731), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g995 ( .A(n_340), .B(n_996), .C(n_999), .Y(n_995) );
AOI211xp5_ASAP7_75t_L g1146 ( .A1(n_340), .A2(n_1138), .B(n_1147), .C(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g518 ( .A(n_341), .Y(n_518) );
BUFx2_ASAP7_75t_L g529 ( .A(n_341), .Y(n_529) );
BUFx2_ASAP7_75t_L g736 ( .A(n_341), .Y(n_736) );
BUFx3_ASAP7_75t_L g830 ( .A(n_341), .Y(n_830) );
BUFx2_ASAP7_75t_L g891 ( .A(n_341), .Y(n_891) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_341), .Y(n_1160) );
INVx1_ASAP7_75t_L g526 ( .A(n_342), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_349), .B1(n_350), .B2(n_353), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_344), .A2(n_350), .B1(n_1413), .B2(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1465 ( .A1(n_344), .A2(n_350), .B1(n_1466), .B2(n_1467), .Y(n_1465) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g943 ( .A(n_345), .Y(n_943) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AND2x4_ASAP7_75t_L g351 ( .A(n_346), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g501 ( .A(n_346), .B(n_348), .Y(n_501) );
AND2x4_ASAP7_75t_L g645 ( .A(n_346), .B(n_348), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_346), .B(n_352), .Y(n_646) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND3x4_ASAP7_75t_L g508 ( .A(n_347), .B(n_366), .C(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_349), .A2(n_385), .B1(n_388), .B2(n_393), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_350), .A2(n_932), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_350), .A2(n_943), .B1(n_1030), .B2(n_1065), .Y(n_1064) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g503 ( .A(n_351), .Y(n_503) );
AOI222xp33_ASAP7_75t_L g732 ( .A1(n_351), .A2(n_645), .B1(n_733), .B2(n_734), .C1(n_735), .C2(n_736), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_351), .A2(n_501), .B1(n_802), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_351), .A2(n_501), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g496 ( .A(n_356), .Y(n_496) );
INVx2_ASAP7_75t_SL g744 ( .A(n_356), .Y(n_744) );
BUFx2_ASAP7_75t_L g939 ( .A(n_356), .Y(n_939) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_358), .A2(n_641), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g498 ( .A(n_359), .Y(n_498) );
BUFx3_ASAP7_75t_L g814 ( .A(n_359), .Y(n_814) );
INVx1_ASAP7_75t_L g1425 ( .A(n_359), .Y(n_1425) );
BUFx3_ASAP7_75t_L g440 ( .A(n_360), .Y(n_440) );
INVx1_ASAP7_75t_L g598 ( .A(n_360), .Y(n_598) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g434 ( .A(n_361), .Y(n_434) );
BUFx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI31xp33_ASAP7_75t_L g937 ( .A1(n_363), .A2(n_938), .A3(n_941), .B(n_945), .Y(n_937) );
OAI31xp33_ASAP7_75t_L g1061 ( .A1(n_363), .A2(n_1062), .A3(n_1063), .B(n_1066), .Y(n_1061) );
OAI31xp33_ASAP7_75t_L g1416 ( .A1(n_363), .A2(n_1417), .A3(n_1420), .B(n_1423), .Y(n_1416) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_364), .B(n_367), .Y(n_363) );
AND2x4_ASAP7_75t_L g505 ( .A(n_364), .B(n_367), .Y(n_505) );
AND2x2_ASAP7_75t_L g649 ( .A(n_364), .B(n_367), .Y(n_649) );
AND2x2_ASAP7_75t_L g815 ( .A(n_364), .B(n_367), .Y(n_815) );
AND2x2_ASAP7_75t_L g843 ( .A(n_364), .B(n_367), .Y(n_843) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g418 ( .A(n_369), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g483 ( .A(n_369), .Y(n_483) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_369), .B(n_481), .Y(n_621) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_394), .A3(n_406), .B(n_411), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_376), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_376), .A2(n_617), .B1(n_1099), .B2(n_1103), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_376), .A2(n_617), .B1(n_1095), .B2(n_1107), .Y(n_1113) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g570 ( .A(n_377), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_377), .A2(n_585), .B1(n_604), .B2(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_377), .A2(n_614), .B1(n_659), .B2(n_660), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_377), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
BUFx2_ASAP7_75t_SL g1407 ( .A(n_377), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_377), .A2(n_956), .B1(n_1441), .B2(n_1453), .Y(n_1458) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_378), .Y(n_476) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR3xp33_ASAP7_75t_L g561 ( .A(n_380), .B(n_562), .C(n_566), .Y(n_561) );
INVx3_ASAP7_75t_L g751 ( .A(n_380), .Y(n_751) );
INVx1_ASAP7_75t_L g1028 ( .A(n_380), .Y(n_1028) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g625 ( .A(n_381), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g628 ( .A(n_381), .B(n_387), .Y(n_628) );
OR2x2_ASAP7_75t_L g851 ( .A(n_381), .B(n_403), .Y(n_851) );
BUFx3_ASAP7_75t_L g868 ( .A(n_382), .Y(n_868) );
BUFx6f_ASAP7_75t_L g1141 ( .A(n_382), .Y(n_1141) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g553 ( .A(n_383), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g1084 ( .A1(n_385), .A2(n_1078), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g402 ( .A(n_386), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g568 ( .A(n_386), .B(n_387), .Y(n_568) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_386), .B(n_873), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_388), .A2(n_568), .B1(n_733), .B2(n_735), .Y(n_752) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g1086 ( .A(n_389), .Y(n_1086) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g631 ( .A(n_390), .Y(n_631) );
BUFx3_ASAP7_75t_L g680 ( .A(n_390), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_390), .A2(n_628), .B1(n_838), .B2(n_840), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_390), .A2(n_628), .B1(n_987), .B2(n_988), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_390), .A2(n_568), .B1(n_1413), .B2(n_1414), .Y(n_1412) );
AOI22xp33_ASAP7_75t_SL g1473 ( .A1(n_390), .A2(n_568), .B1(n_1466), .B2(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_396), .Y(n_563) );
AND2x4_ASAP7_75t_L g408 ( .A(n_397), .B(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_400), .A2(n_1132), .B1(n_1133), .B2(n_1134), .C(n_1135), .Y(n_1131) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_401), .Y(n_935) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g565 ( .A(n_402), .Y(n_565) );
INVx2_ASAP7_75t_L g749 ( .A(n_402), .Y(n_749) );
INVx8_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
BUFx2_ASAP7_75t_L g723 ( .A(n_403), .Y(n_723) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_408), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_408), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
INVx4_ASAP7_75t_L g886 ( .A(n_408), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_408), .A2(n_847), .B1(n_982), .B2(n_983), .Y(n_981) );
INVx3_ASAP7_75t_SL g1471 ( .A(n_408), .Y(n_1471) );
INVx2_ASAP7_75t_L g550 ( .A(n_409), .Y(n_550) );
BUFx6f_ASAP7_75t_L g867 ( .A(n_409), .Y(n_867) );
OAI31xp33_ASAP7_75t_L g1024 ( .A1(n_411), .A2(n_1025), .A3(n_1026), .B(n_1032), .Y(n_1024) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g571 ( .A(n_412), .Y(n_571) );
BUFx2_ASAP7_75t_L g637 ( .A(n_412), .Y(n_637) );
OAI31xp33_ASAP7_75t_L g879 ( .A1(n_412), .A2(n_880), .A3(n_881), .B(n_885), .Y(n_879) );
BUFx2_ASAP7_75t_SL g1089 ( .A(n_412), .Y(n_1089) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_454), .Y(n_415) );
OAI33xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .A3(n_426), .B1(n_435), .B2(n_442), .B3(n_448), .Y(n_416) );
OAI33xp33_ASAP7_75t_L g697 ( .A1(n_417), .A2(n_698), .A3(n_702), .B1(n_707), .B2(n_712), .B3(n_713), .Y(n_697) );
OAI33xp33_ASAP7_75t_L g1091 ( .A1(n_417), .A2(n_712), .A3(n_1092), .B1(n_1098), .B2(n_1101), .B3(n_1105), .Y(n_1091) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_417), .A2(n_1155), .B1(n_1161), .B2(n_1164), .Y(n_1154) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx4f_ASAP7_75t_L g581 ( .A(n_418), .Y(n_581) );
BUFx8_ASAP7_75t_L g785 ( .A(n_418), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_449), .B1(n_461), .B2(n_465), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_422), .A2(n_449), .B1(n_450), .B2(n_453), .Y(n_448) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_422), .A2(n_670), .B1(n_714), .B2(n_715), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_422), .A2(n_949), .B1(n_957), .B2(n_968), .Y(n_967) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_422), .A2(n_1050), .B1(n_1051), .B2(n_1052), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_422), .A2(n_1389), .B1(n_1390), .B2(n_1391), .Y(n_1388) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_422), .A2(n_968), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
OAI22xp33_ASAP7_75t_L g1439 ( .A1(n_422), .A2(n_1391), .B1(n_1440), .B2(n_1441), .Y(n_1439) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_422), .A2(n_916), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_423), .A2(n_453), .B1(n_469), .B2(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g586 ( .A(n_425), .Y(n_586) );
INVx2_ASAP7_75t_L g797 ( .A(n_425), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_431), .B2(n_432), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_427), .A2(n_439), .B1(n_469), .B2(n_474), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_428), .A2(n_432), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1442 ( .A1(n_428), .A2(n_1443), .B1(n_1444), .B2(n_1445), .Y(n_1442) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx8_ASAP7_75t_L g1046 ( .A(n_429), .Y(n_1046) );
INVx5_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
INVx2_ASAP7_75t_SL g673 ( .A(n_430), .Y(n_673) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_430), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_431), .A2(n_441), .B1(n_461), .B2(n_465), .Y(n_484) );
OAI22xp33_ASAP7_75t_SL g793 ( .A1(n_432), .A2(n_772), .B1(n_783), .B2(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_432), .A2(n_1448), .B1(n_1449), .B2(n_1450), .Y(n_1447) );
CKINVDCx8_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g591 ( .A(n_433), .Y(n_591) );
INVx3_ASAP7_75t_L g674 ( .A(n_433), .Y(n_674) );
INVx3_ASAP7_75t_L g914 ( .A(n_433), .Y(n_914) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g705 ( .A(n_434), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_438), .A2(n_591), .B1(n_901), .B2(n_908), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_440), .A2(n_768), .B1(n_781), .B2(n_792), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_440), .A2(n_952), .B1(n_962), .B2(n_970), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_440), .A2(n_589), .B1(n_954), .B2(n_965), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_440), .A2(n_589), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_440), .A2(n_1044), .B1(n_1045), .B2(n_1047), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1155 ( .A1(n_440), .A2(n_1119), .B1(n_1156), .B2(n_1157), .C(n_1158), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_440), .A2(n_1396), .B1(n_1397), .B2(n_1398), .Y(n_1395) );
INVx1_ASAP7_75t_L g533 ( .A(n_442), .Y(n_533) );
OAI33xp33_ASAP7_75t_L g966 ( .A1(n_442), .A2(n_785), .A3(n_967), .B1(n_969), .B2(n_971), .B3(n_972), .Y(n_966) );
OAI33xp33_ASAP7_75t_L g1387 ( .A1(n_442), .A2(n_785), .A3(n_1388), .B1(n_1392), .B2(n_1395), .B3(n_1399), .Y(n_1387) );
OAI33xp33_ASAP7_75t_L g1438 ( .A1(n_442), .A2(n_785), .A3(n_1439), .B1(n_1442), .B2(n_1447), .B3(n_1451), .Y(n_1438) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g795 ( .A(n_443), .Y(n_795) );
INVx2_ASAP7_75t_L g1048 ( .A(n_443), .Y(n_1048) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g1166 ( .A(n_444), .Y(n_1166) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g1097 ( .A(n_452), .Y(n_1097) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_460), .A3(n_468), .B1(n_477), .B2(n_479), .B3(n_484), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
INVx2_ASAP7_75t_L g608 ( .A(n_456), .Y(n_608) );
INVx4_ASAP7_75t_L g720 ( .A(n_456), .Y(n_720) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
OR2x2_ASAP7_75t_L g605 ( .A(n_457), .B(n_606), .Y(n_605) );
OR2x6_ASAP7_75t_L g712 ( .A(n_457), .B(n_606), .Y(n_712) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_461), .A2(n_1036), .B1(n_1050), .B2(n_1055), .Y(n_1054) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g610 ( .A(n_464), .Y(n_610) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_464), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_465), .A2(n_780), .B1(n_949), .B2(n_950), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_465), .A2(n_961), .B1(n_1394), .B2(n_1398), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1459 ( .A1(n_465), .A2(n_780), .B1(n_1444), .B2(n_1450), .Y(n_1459) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g612 ( .A(n_467), .Y(n_612) );
INVx4_ASAP7_75t_L g619 ( .A(n_467), .Y(n_619) );
INVx2_ASAP7_75t_SL g656 ( .A(n_467), .Y(n_656) );
INVx2_ASAP7_75t_L g782 ( .A(n_467), .Y(n_782) );
INVx1_ASAP7_75t_L g964 ( .A(n_467), .Y(n_964) );
INVx1_ASAP7_75t_L g1055 ( .A(n_467), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_469), .A2(n_701), .B1(n_715), .B2(n_725), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_469), .A2(n_569), .B1(n_1393), .B2(n_1396), .Y(n_1405) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g614 ( .A(n_471), .Y(n_614) );
INVx2_ASAP7_75t_L g953 ( .A(n_471), .Y(n_953) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g617 ( .A(n_472), .Y(n_617) );
BUFx2_ASAP7_75t_L g771 ( .A(n_472), .Y(n_771) );
INVx1_ASAP7_75t_L g776 ( .A(n_472), .Y(n_776) );
AND2x2_ASAP7_75t_L g541 ( .A(n_473), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_475), .Y(n_478) );
INVx2_ASAP7_75t_L g615 ( .A(n_475), .Y(n_615) );
INVx1_ASAP7_75t_L g725 ( .A(n_475), .Y(n_725) );
INVx2_ASAP7_75t_L g800 ( .A(n_475), .Y(n_800) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_476), .Y(n_663) );
BUFx4f_ASAP7_75t_L g773 ( .A(n_476), .Y(n_773) );
BUFx4f_ASAP7_75t_L g905 ( .A(n_476), .Y(n_905) );
OAI33xp33_ASAP7_75t_L g761 ( .A1(n_479), .A2(n_720), .A3(n_762), .B1(n_767), .B2(n_774), .B3(n_779), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
AOI33xp33_ASAP7_75t_L g534 ( .A1(n_480), .A2(n_535), .A3(n_538), .B1(n_546), .B2(n_554), .B3(n_555), .Y(n_534) );
INVx2_ASAP7_75t_L g959 ( .A(n_480), .Y(n_959) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_481), .B(n_482), .Y(n_1129) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND4xp25_ASAP7_75t_SL g488 ( .A(n_489), .B(n_506), .C(n_534), .D(n_559), .Y(n_488) );
AO21x1_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_494), .B(n_504), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_492), .A2(n_641), .B1(n_982), .B2(n_983), .Y(n_994) );
INVx1_ASAP7_75t_L g1153 ( .A(n_496), .Y(n_1153) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g940 ( .A(n_498), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g1152 ( .A1(n_498), .A2(n_1133), .B1(n_1134), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_502), .A2(n_1036), .B1(n_1037), .B2(n_1039), .Y(n_1035) );
AOI31xp33_ASAP7_75t_L g729 ( .A1(n_504), .A2(n_730), .A3(n_737), .B(n_740), .Y(n_729) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AOI33xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .A3(n_519), .B1(n_527), .B2(n_530), .B3(n_533), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g826 ( .A(n_508), .Y(n_826) );
BUFx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_513), .A2(n_829), .B1(n_831), .B2(n_832), .C(n_833), .Y(n_828) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx8_ASAP7_75t_L g823 ( .A(n_515), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_517), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g1147 ( .A(n_518), .Y(n_1147) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_521), .A2(n_703), .B1(n_704), .B2(n_706), .Y(n_702) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g531 ( .A(n_522), .Y(n_531) );
INVx3_ASAP7_75t_L g595 ( .A(n_522), .Y(n_595) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g532 ( .A(n_524), .Y(n_532) );
INVx5_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx12f_ASAP7_75t_L g1016 ( .A(n_525), .Y(n_1016) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g1397 ( .A(n_531), .Y(n_1397) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_536), .A2(n_1118), .B1(n_1123), .B2(n_1129), .Y(n_1117) );
OAI33xp33_ASAP7_75t_L g1402 ( .A1(n_536), .A2(n_959), .A3(n_1403), .B1(n_1405), .B2(n_1406), .B3(n_1408), .Y(n_1402) );
OAI33xp33_ASAP7_75t_L g1454 ( .A1(n_536), .A2(n_959), .A3(n_1455), .B1(n_1456), .B2(n_1458), .B3(n_1459), .Y(n_1454) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI33xp33_ASAP7_75t_L g653 ( .A1(n_537), .A2(n_620), .A3(n_654), .B1(n_658), .B2(n_661), .B3(n_665), .Y(n_653) );
OAI33xp33_ASAP7_75t_L g896 ( .A1(n_537), .A2(n_620), .A3(n_897), .B1(n_900), .B2(n_903), .B3(n_907), .Y(n_896) );
OAI33xp33_ASAP7_75t_L g1053 ( .A1(n_537), .A2(n_959), .A3(n_1054), .B1(n_1056), .B2(n_1057), .B3(n_1060), .Y(n_1053) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_SL g556 ( .A(n_540), .Y(n_556) );
INVx2_ASAP7_75t_L g864 ( .A(n_540), .Y(n_864) );
INVx1_ASAP7_75t_L g1010 ( .A(n_540), .Y(n_1010) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_541), .Y(n_873) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g558 ( .A(n_545), .Y(n_558) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_545), .Y(n_1011) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g990 ( .A(n_552), .Y(n_990) );
INVx2_ASAP7_75t_L g1007 ( .A(n_552), .Y(n_1007) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g626 ( .A(n_553), .Y(n_626) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g1122 ( .A(n_558), .Y(n_1122) );
AO21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_571), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_568), .A2(n_630), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_568), .A2(n_680), .B1(n_883), .B2(n_884), .Y(n_882) );
BUFx3_ASAP7_75t_L g931 ( .A(n_568), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_569), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_569), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_569), .A2(n_956), .B1(n_1041), .B2(n_1044), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_569), .A2(n_1039), .B1(n_1052), .B2(n_1058), .Y(n_1057) );
INVx5_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AO21x1_ASAP7_75t_L g844 ( .A1(n_571), .A2(n_845), .B(n_849), .Y(n_844) );
AO21x1_ASAP7_75t_L g980 ( .A1(n_571), .A2(n_981), .B(n_984), .Y(n_980) );
AOI21xp33_ASAP7_75t_L g1130 ( .A1(n_571), .A2(n_1131), .B(n_1142), .Y(n_1130) );
XOR2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_691), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
XNOR2x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_650), .Y(n_575) );
XNOR2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND3x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_622), .C(n_638), .Y(n_578) );
NOR2xp33_ASAP7_75t_SL g579 ( .A(n_580), .B(n_607), .Y(n_579) );
OAI33xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .A3(n_587), .B1(n_592), .B2(n_599), .B3(n_605), .Y(n_580) );
OAI33xp33_ASAP7_75t_L g668 ( .A1(n_581), .A2(n_605), .A3(n_669), .B1(n_671), .B2(n_672), .B3(n_675), .Y(n_668) );
OAI33xp33_ASAP7_75t_L g910 ( .A1(n_581), .A2(n_605), .A3(n_911), .B1(n_912), .B2(n_913), .B3(n_915), .Y(n_910) );
OAI33xp33_ASAP7_75t_L g1034 ( .A1(n_581), .A2(n_1035), .A3(n_1040), .B1(n_1043), .B2(n_1048), .B3(n_1049), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_583), .A2(n_602), .B1(n_610), .B2(n_611), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g915 ( .A1(n_584), .A2(n_899), .B1(n_906), .B2(n_916), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_586), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_588), .A2(n_593), .B1(n_614), .B2(n_615), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_589), .A2(n_591), .B1(n_659), .B2(n_666), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_589), .A2(n_902), .B1(n_909), .B2(n_914), .Y(n_913) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_589), .A2(n_914), .B1(n_1120), .B2(n_1162), .C(n_1163), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_590), .A2(n_596), .B1(n_610), .B2(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_596), .B2(n_597), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g792 ( .A(n_595), .Y(n_792) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g1446 ( .A(n_598), .Y(n_1446) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_600), .A2(n_655), .B1(n_662), .B2(n_670), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_600), .A2(n_603), .B1(n_657), .B2(n_664), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_600), .A2(n_603), .B1(n_898), .B2(n_904), .Y(n_911) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx3_ASAP7_75t_L g699 ( .A(n_601), .Y(n_699) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_603), .Y(n_968) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_603), .Y(n_1051) );
INVx2_ASAP7_75t_L g1076 ( .A(n_603), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_603), .A2(n_699), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_603), .Y(n_1391) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .A3(n_613), .B1(n_616), .B2(n_618), .B3(n_620), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_610), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_610), .A2(n_611), .B1(n_666), .B2(n_667), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_610), .A2(n_611), .B1(n_898), .B2(n_899), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_610), .A2(n_656), .B1(n_908), .B2(n_909), .Y(n_907) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_614), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_614), .A2(n_663), .B1(n_901), .B2(n_902), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_614), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_617), .A2(n_703), .B1(n_710), .B2(n_725), .Y(n_724) );
OAI33xp33_ASAP7_75t_L g717 ( .A1(n_620), .A2(n_718), .A3(n_721), .B1(n_724), .B2(n_726), .B3(n_727), .Y(n_717) );
OAI33xp33_ASAP7_75t_L g1108 ( .A1(n_620), .A2(n_720), .A3(n_1109), .B1(n_1112), .B2(n_1113), .B3(n_1114), .Y(n_1108) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI33xp33_ASAP7_75t_L g862 ( .A1(n_621), .A2(n_719), .A3(n_863), .B1(n_865), .B2(n_869), .B3(n_870), .Y(n_862) );
AOI33xp33_ASAP7_75t_L g1001 ( .A1(n_621), .A2(n_1002), .A3(n_1003), .B1(n_1004), .B2(n_1008), .B3(n_1009), .Y(n_1001) );
OAI31xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_633), .A3(n_636), .B(n_637), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g857 ( .A(n_625), .Y(n_857) );
INVx1_ASAP7_75t_L g856 ( .A(n_626), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_630), .B2(n_632), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_628), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_628), .A2(n_630), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_629), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_630), .A2(n_931), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g847 ( .A(n_634), .Y(n_847) );
BUFx3_ASAP7_75t_L g780 ( .A(n_635), .Y(n_780) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_635), .Y(n_1111) );
OAI31xp33_ASAP7_75t_L g676 ( .A1(n_637), .A2(n_677), .A3(n_682), .B(n_683), .Y(n_676) );
INVx1_ASAP7_75t_L g755 ( .A(n_637), .Y(n_755) );
OAI31xp33_ASAP7_75t_L g798 ( .A1(n_637), .A2(n_799), .A3(n_804), .B(n_806), .Y(n_798) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_637), .A2(n_927), .A3(n_934), .B(n_936), .Y(n_926) );
OAI31xp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_642), .A3(n_648), .B(n_649), .Y(n_638) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g836 ( .A(n_643), .B(n_837), .C(n_839), .Y(n_836) );
NAND3xp33_ASAP7_75t_SL g889 ( .A(n_643), .B(n_890), .C(n_892), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_645), .A2(n_646), .B1(n_679), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_645), .A2(n_646), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_645), .A2(n_646), .B1(n_883), .B2(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_645), .B(n_987), .Y(n_998) );
INVx1_ASAP7_75t_L g1149 ( .A(n_645), .Y(n_1149) );
INVx1_ASAP7_75t_L g997 ( .A(n_646), .Y(n_997) );
INVxp67_ASAP7_75t_L g1150 ( .A(n_646), .Y(n_1150) );
OAI31xp33_ASAP7_75t_SL g685 ( .A1(n_649), .A2(n_686), .A3(n_687), .B(n_690), .Y(n_685) );
AND3x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_676), .C(n_685), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_668), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_656), .A2(n_706), .B1(n_711), .B2(n_722), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_656), .A2(n_763), .B1(n_764), .B2(n_766), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_656), .A2(n_1100), .B1(n_1104), .B2(n_1110), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_660), .A2(n_667), .B1(n_673), .B2(n_674), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_663), .A2(n_956), .B1(n_1124), .B2(n_1125), .C(n_1126), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_674), .A2(n_792), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_680), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_817), .B2(n_917), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_757), .B1(n_758), .B2(n_816), .Y(n_693) );
INVx1_ASAP7_75t_L g816 ( .A(n_694), .Y(n_816) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR4xp25_ASAP7_75t_L g756 ( .A(n_697), .B(n_717), .C(n_729), .D(n_745), .Y(n_756) );
BUFx4f_ASAP7_75t_SL g1094 ( .A(n_699), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_700), .A2(n_714), .B1(n_722), .B2(n_723), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_704), .A2(n_708), .B1(n_710), .B2(n_711), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_704), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1101) );
BUFx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_709), .Y(n_1102) );
INVx1_ASAP7_75t_L g833 ( .A(n_712), .Y(n_833) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OAI33xp33_ASAP7_75t_L g947 ( .A1(n_720), .A2(n_948), .A3(n_951), .B1(n_955), .B2(n_959), .B3(n_960), .Y(n_947) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_720), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_723), .A2(n_1093), .B1(n_1106), .B2(n_1110), .Y(n_1109) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx2_ASAP7_75t_L g1067 ( .A(n_744), .Y(n_1067) );
AOI31xp67_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_750), .A3(n_753), .B(n_755), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_SL g805 ( .A(n_749), .Y(n_805) );
INVx1_ASAP7_75t_L g1476 ( .A(n_749), .Y(n_1476) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_798), .C(n_807), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_784), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_763), .A2(n_777), .B1(n_787), .B2(n_790), .Y(n_786) );
INVx3_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g961 ( .A(n_765), .Y(n_961) );
INVx2_ASAP7_75t_L g1404 ( .A(n_765), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_766), .A2(n_778), .B1(n_787), .B2(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_769), .B1(n_772), .B2(n_773), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g956 ( .A(n_770), .Y(n_956) );
INVx4_ASAP7_75t_L g1457 ( .A(n_770), .Y(n_1457) );
INVx4_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g929 ( .A(n_773), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_775), .A2(n_905), .B1(n_1119), .B2(n_1120), .C(n_1121), .Y(n_1118) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_779) );
OAI33xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .A3(n_791), .B1(n_793), .B2(n_795), .B3(n_796), .Y(n_784) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g974 ( .A(n_789), .Y(n_974) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_789), .Y(n_1038) );
OAI31xp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .A3(n_813), .B(n_815), .Y(n_807) );
OAI31xp33_ASAP7_75t_L g1460 ( .A1(n_815), .A2(n_1461), .A3(n_1463), .B(n_1468), .Y(n_1460) );
INVx2_ASAP7_75t_L g917 ( .A(n_817), .Y(n_917) );
XNOR2x1_ASAP7_75t_L g817 ( .A(n_818), .B(n_877), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_858), .Y(n_818) );
INVx1_ASAP7_75t_L g860 ( .A(n_820), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_824), .B(n_827), .Y(n_820) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx8_ASAP7_75t_L g1018 ( .A(n_823), .Y(n_1018) );
INVx3_ASAP7_75t_L g1159 ( .A(n_823), .Y(n_1159) );
INVx1_ASAP7_75t_L g970 ( .A(n_825), .Y(n_970) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI32xp33_ASAP7_75t_L g1012 ( .A1(n_833), .A2(n_1013), .A3(n_1017), .B1(n_1019), .B2(n_1020), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_834), .B(n_844), .Y(n_859) );
OAI31xp33_ASAP7_75t_SL g834 ( .A1(n_835), .A2(n_836), .A3(n_842), .B(n_843), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_841), .B(n_855), .Y(n_854) );
OAI31xp33_ASAP7_75t_SL g887 ( .A1(n_843), .A2(n_888), .A3(n_889), .B(n_894), .Y(n_887) );
INVx1_ASAP7_75t_L g1000 ( .A(n_843), .Y(n_1000) );
OAI31xp33_ASAP7_75t_L g1072 ( .A1(n_843), .A2(n_1073), .A3(n_1074), .B(n_1080), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_852), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .C(n_857), .Y(n_852) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_857), .B(n_986), .C(n_989), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g1135 ( .A(n_857), .B(n_1136), .C(n_1139), .Y(n_1135) );
OAI31xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .A3(n_861), .B(n_874), .Y(n_858) );
INVx1_ASAP7_75t_L g876 ( .A(n_862), .Y(n_876) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g1006 ( .A(n_867), .Y(n_1006) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
NAND3xp33_ASAP7_75t_SL g878 ( .A(n_879), .B(n_887), .C(n_895), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_884), .B(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_910), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_905), .A2(n_1443), .B1(n_1448), .B2(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_921), .B1(n_1068), .B2(n_1069), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
XNOR2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_975), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_937), .C(n_946), .Y(n_925) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NOR2xp33_ASAP7_75t_SL g946 ( .A(n_947), .B(n_966), .Y(n_946) );
INVx1_ASAP7_75t_L g1059 ( .A(n_953), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_956), .A2(n_1390), .B1(n_1401), .B2(n_1407), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_962), .B1(n_963), .B2(n_965), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_961), .A2(n_963), .B1(n_1042), .B2(n_1047), .Y(n_1060) );
BUFx3_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_1021), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
NAND4xp75_ASAP7_75t_L g979 ( .A(n_980), .B(n_993), .C(n_1001), .D(n_1012), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_992), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
AO21x1_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .B(n_1000), .Y(n_993) );
AOI31xp33_ASAP7_75t_L g1145 ( .A1(n_1000), .A2(n_1146), .A3(n_1151), .B(n_1152), .Y(n_1145) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1011), .Y(n_1128) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
AND3x1_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1033), .C(n_1061), .Y(n_1023) );
NOR2xp33_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1053), .Y(n_1033) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1403 ( .A1(n_1055), .A2(n_1389), .B1(n_1400), .B2(n_1404), .Y(n_1403) );
OAI22xp33_ASAP7_75t_L g1455 ( .A1(n_1055), .A2(n_1404), .B1(n_1440), .B2(n_1452), .Y(n_1455) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
XNOR2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1115), .Y(n_1069) );
NAND3xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1082), .C(n_1090), .Y(n_1071) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
OAI31xp33_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1087), .A3(n_1088), .B(n_1089), .Y(n_1082) );
OAI31xp33_ASAP7_75t_L g1409 ( .A1(n_1089), .A2(n_1410), .A3(n_1411), .B(n_1415), .Y(n_1409) );
OAI31xp33_ASAP7_75t_L g1469 ( .A1(n_1089), .A2(n_1470), .A3(n_1472), .B(n_1475), .Y(n_1469) );
NOR2xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1108), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1092) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1097), .Y(n_1464) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NOR4xp25_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1130), .C(n_1145), .D(n_1154), .Y(n_1116) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OAI221xp5_ASAP7_75t_SL g1167 ( .A1(n_1168), .A2(n_1381), .B1(n_1383), .B2(n_1426), .C(n_1430), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1272), .B(n_1293), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1189), .B(n_1220), .C(n_1258), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1185), .Y(n_1170) );
INVx3_ASAP7_75t_L g1229 ( .A(n_1171), .Y(n_1229) );
INVx3_ASAP7_75t_L g1269 ( .A(n_1171), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1271 ( .A(n_1171), .B(n_1246), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1171), .B(n_1292), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1171), .B(n_1314), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1171), .B(n_1185), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1171), .B(n_1238), .Y(n_1338) );
AND2x4_ASAP7_75t_SL g1171 ( .A(n_1172), .B(n_1179), .Y(n_1171) );
AND2x6_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1174), .B(n_1178), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1174), .B(n_1181), .Y(n_1180) );
AND2x6_ASAP7_75t_L g1183 ( .A(n_1174), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1174), .B(n_1178), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1174), .B(n_1178), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1176), .B(n_1182), .Y(n_1181) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1177), .Y(n_1382) );
OAI21xp5_ASAP7_75t_L g1477 ( .A1(n_1178), .A2(n_1478), .B(n_1479), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1185), .B(n_1214), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1185), .B(n_1269), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1185), .B(n_1213), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1185), .B(n_1214), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1185), .B(n_1300), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1188), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1233 ( .A(n_1186), .B(n_1188), .Y(n_1233) );
AOI211xp5_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1198), .B(n_1206), .C(n_1211), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1190), .B(n_1250), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1190), .B(n_1245), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1190), .B(n_1210), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1194), .Y(n_1190) );
INVx3_ASAP7_75t_L g1209 ( .A(n_1191), .Y(n_1209) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1191), .Y(n_1242) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1191), .B(n_1194), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1191), .B(n_1326), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1191), .B(n_1213), .Y(n_1341) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1191), .B(n_1362), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1194), .B(n_1237), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1194), .B(n_1219), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g1254 ( .A(n_1194), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1194), .B(n_1253), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1194), .B(n_1260), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1194), .B(n_1250), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1197), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1195), .B(n_1197), .Y(n_1222) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1198), .Y(n_1245) );
NOR2xp33_ASAP7_75t_L g1345 ( .A(n_1198), .B(n_1209), .Y(n_1345) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1202), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1199), .B(n_1202), .Y(n_1210) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1199), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1199), .B(n_1203), .Y(n_1250) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1199), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1201), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1202), .B(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1202), .Y(n_1237) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1203), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1205), .Y(n_1203) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1210), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1208), .B(n_1236), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1208), .B(n_1238), .Y(n_1255) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1209), .B(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1209), .B(n_1210), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1209), .B(n_1265), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1209), .B(n_1305), .Y(n_1327) );
OAI21xp33_ASAP7_75t_L g1330 ( .A1(n_1209), .A2(n_1321), .B(n_1331), .Y(n_1330) );
NOR2xp33_ASAP7_75t_L g1349 ( .A(n_1209), .B(n_1350), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1209), .B(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1210), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1210), .B(n_1276), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1217), .Y(n_1211) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1212), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1213), .B(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1214), .Y(n_1247) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1214), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
NOR3xp33_ASAP7_75t_L g1340 ( .A(n_1217), .B(n_1269), .C(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1218), .B(n_1254), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1218), .B(n_1338), .Y(n_1337) );
OAI32xp33_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1224), .A3(n_1228), .B1(n_1230), .B2(n_1256), .Y(n_1220) );
AOI332xp33_ASAP7_75t_L g1346 ( .A1(n_1221), .A2(n_1229), .A3(n_1286), .B1(n_1292), .B2(n_1314), .B3(n_1347), .C1(n_1349), .C2(n_1351), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1222), .B(n_1245), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1222), .B(n_1290), .Y(n_1321) );
AOI22xp5_ASAP7_75t_SL g1231 ( .A1(n_1223), .A2(n_1232), .B1(n_1234), .B2(n_1238), .Y(n_1231) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1224), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1224), .B(n_1229), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_1224), .A2(n_1225), .B1(n_1360), .B2(n_1368), .Y(n_1359) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AOI211xp5_ASAP7_75t_L g1274 ( .A1(n_1225), .A2(n_1275), .B(n_1277), .C(n_1278), .Y(n_1274) );
O2A1O1Ixp33_ASAP7_75t_SL g1316 ( .A1(n_1225), .A2(n_1317), .B(n_1318), .C(n_1319), .Y(n_1316) );
O2A1O1Ixp33_ASAP7_75t_L g1323 ( .A1(n_1225), .A2(n_1324), .B(n_1334), .C(n_1342), .Y(n_1323) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1225), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1228), .B(n_1257), .Y(n_1256) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1272 ( .A1(n_1229), .A2(n_1273), .B1(n_1274), .B2(n_1281), .C(n_1282), .Y(n_1272) );
AOI22xp5_ASAP7_75t_L g1357 ( .A1(n_1229), .A2(n_1358), .B1(n_1359), .B2(n_1372), .Y(n_1357) );
INVxp67_ASAP7_75t_SL g1273 ( .A(n_1230), .Y(n_1273) );
NAND4xp25_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1239), .C(n_1248), .D(n_1251), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1232), .B(n_1249), .Y(n_1248) );
NAND2xp5_ASAP7_75t_SL g1262 ( .A(n_1232), .B(n_1242), .Y(n_1262) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1232), .Y(n_1317) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1233), .Y(n_1292) );
CKINVDCx6p67_ASAP7_75t_R g1297 ( .A(n_1233), .Y(n_1297) );
NOR2xp33_ASAP7_75t_L g1351 ( .A(n_1233), .B(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
AOI21xp33_ASAP7_75t_L g1366 ( .A1(n_1235), .A2(n_1241), .B(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1236), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1237), .B(n_1254), .Y(n_1265) );
CKINVDCx14_ASAP7_75t_R g1367 ( .A(n_1238), .Y(n_1367) );
OAI21xp5_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1244), .B(n_1246), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_1240), .A2(n_1329), .B1(n_1330), .B2(n_1332), .Y(n_1328) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1243), .Y(n_1241) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1242), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1242), .B(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_SL g1356 ( .A(n_1242), .B(n_1245), .Y(n_1356) );
CKINVDCx14_ASAP7_75t_R g1306 ( .A(n_1243), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1336 ( .A(n_1244), .Y(n_1336) );
OAI21xp5_ASAP7_75t_L g1251 ( .A1(n_1245), .A2(n_1252), .B(n_1255), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1245), .B(n_1276), .Y(n_1275) );
OAI21xp5_ASAP7_75t_L g1319 ( .A1(n_1245), .A2(n_1255), .B(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1246), .Y(n_1280) );
OAI21xp33_ASAP7_75t_L g1353 ( .A1(n_1246), .A2(n_1291), .B(n_1354), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1246), .B(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
OAI21xp5_ASAP7_75t_SL g1311 ( .A1(n_1247), .A2(n_1312), .B(n_1313), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1249), .B(n_1280), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1250), .B(n_1254), .Y(n_1305) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1250), .Y(n_1362) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1252), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1254), .B(n_1290), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1254), .B(n_1345), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1254), .B(n_1356), .Y(n_1355) );
A2O1A1Ixp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1261), .B(n_1263), .C(n_1266), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1260), .B(n_1276), .Y(n_1318) );
INVxp67_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1270), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1269), .B(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1277), .B(n_1310), .Y(n_1309) );
A2O1A1Ixp33_ASAP7_75t_L g1324 ( .A1(n_1277), .A2(n_1325), .B(n_1327), .C(n_1328), .Y(n_1324) );
INVx2_ASAP7_75t_SL g1365 ( .A(n_1277), .Y(n_1365) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AOI211xp5_ASAP7_75t_L g1294 ( .A1(n_1281), .A2(n_1295), .B(n_1316), .C(n_1322), .Y(n_1294) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1286), .B1(n_1288), .B2(n_1291), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1284), .B(n_1289), .Y(n_1322) );
OAI211xp5_ASAP7_75t_SL g1342 ( .A1(n_1284), .A2(n_1343), .B(n_1346), .C(n_1353), .Y(n_1342) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1285), .Y(n_1348) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1363 ( .A(n_1290), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1291), .Y(n_1335) );
A2O1A1Ixp33_ASAP7_75t_L g1372 ( .A1(n_1292), .A2(n_1315), .B(n_1373), .C(n_1374), .Y(n_1372) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_1292), .A2(n_1365), .B1(n_1375), .B2(n_1376), .C(n_1379), .Y(n_1374) );
NAND3xp33_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1323), .C(n_1357), .Y(n_1293) );
OAI211xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1298), .B(n_1302), .C(n_1311), .Y(n_1295) );
CKINVDCx6p67_ASAP7_75t_R g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
AOI211xp5_ASAP7_75t_L g1368 ( .A1(n_1299), .A2(n_1314), .B(n_1369), .C(n_1370), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1301), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1300), .B(n_1350), .Y(n_1369) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1301), .Y(n_1310) );
AOI21xp5_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1307), .B(n_1309), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1306), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1305), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1327), .Y(n_1375) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
OAI211xp5_ASAP7_75t_L g1334 ( .A1(n_1335), .A2(n_1336), .B(n_1337), .C(n_1339), .Y(n_1334) );
INVxp67_ASAP7_75t_SL g1339 ( .A(n_1340), .Y(n_1339) );
NAND2xp5_ASAP7_75t_SL g1376 ( .A(n_1343), .B(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AOI211xp5_ASAP7_75t_L g1360 ( .A1(n_1348), .A2(n_1361), .B(n_1363), .C(n_1366), .Y(n_1360) );
INVxp67_ASAP7_75t_L g1358 ( .A(n_1351), .Y(n_1358) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1370), .Y(n_1373) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx4_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
BUFx2_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
AND3x1_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1409), .C(n_1416), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1402), .Y(n_1386) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
BUFx3_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
BUFx3_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVxp33_ASAP7_75t_SL g1433 ( .A(n_1434), .Y(n_1433) );
HB1xp67_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
NAND3xp33_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1460), .C(n_1469), .Y(n_1436) );
NOR2xp33_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1454), .Y(n_1437) );
INVx3_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
endmodule