module fake_netlist_1_4235_n_523 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_523);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_523;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g74 ( .A(n_36), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_33), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_55), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_16), .Y(n_77) );
CKINVDCx14_ASAP7_75t_R g78 ( .A(n_14), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_61), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_64), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_53), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_7), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_57), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_47), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_2), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_39), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_37), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_27), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_5), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_17), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_65), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_45), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_13), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_6), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_51), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_22), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_31), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_78), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_89), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_79), .B(n_0), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_84), .B(n_0), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_75), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_97), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_97), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_97), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_82), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_82), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_115), .B(n_76), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_123), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_119), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_111), .B(n_76), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_123), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_132), .A2(n_105), .B1(n_106), .B2(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
INVxp67_ASAP7_75t_SL g142 ( .A(n_115), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_116), .A2(n_110), .B(n_83), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_112), .B(n_88), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_119), .B(n_84), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_126), .A2(n_110), .B(n_83), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_119), .B(n_85), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_111), .B(n_85), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
OAI22xp33_ASAP7_75t_L g156 ( .A1(n_132), .A2(n_98), .B1(n_77), .B2(n_100), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_121), .B(n_101), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_142), .B(n_74), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_139), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_142), .B(n_74), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_155), .B(n_113), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_145), .Y(n_165) );
BUFx8_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_155), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_134), .A2(n_122), .B1(n_113), .B2(n_114), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_134), .Y(n_170) );
AO22x1_ASAP7_75t_L g171 ( .A1(n_134), .A2(n_90), .B1(n_87), .B2(n_103), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_134), .B(n_144), .Y(n_172) );
OAI21xp33_ASAP7_75t_L g173 ( .A1(n_152), .A2(n_114), .B(n_131), .Y(n_173) );
OR2x6_ASAP7_75t_L g174 ( .A(n_145), .B(n_77), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_139), .B(n_98), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_146), .B(n_108), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
NOR2x1p5_ASAP7_75t_L g185 ( .A(n_156), .B(n_102), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_144), .B(n_125), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_144), .B(n_125), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_146), .B(n_124), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_134), .Y(n_189) );
BUFx10_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_166), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_185), .A2(n_134), .B1(n_148), .B2(n_144), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_170), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_170), .B(n_158), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_185), .A2(n_148), .B1(n_144), .B2(n_156), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_190), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_167), .B(n_148), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_190), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_189), .B(n_148), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_177), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
NOR2xp33_ASAP7_75t_SL g205 ( .A(n_166), .B(n_136), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
CKINVDCx11_ASAP7_75t_R g207 ( .A(n_177), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g208 ( .A(n_178), .B(n_136), .Y(n_208) );
AOI221xp5_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_148), .B1(n_100), .B2(n_158), .C(n_128), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_190), .Y(n_210) );
NOR2x1_ASAP7_75t_L g211 ( .A(n_172), .B(n_137), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_180), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_186), .A2(n_151), .B(n_152), .C(n_154), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_177), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_172), .A2(n_177), .B1(n_167), .B2(n_178), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_189), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_177), .B(n_158), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_172), .A2(n_158), .B1(n_137), .B2(n_136), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_160), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_204), .Y(n_223) );
BUFx12f_ASAP7_75t_L g224 ( .A(n_207), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_195), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_219), .B(n_159), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_196), .B(n_163), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_204), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_216), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_214), .A2(n_187), .B(n_186), .Y(n_230) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_191), .B(n_172), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_219), .A2(n_161), .B1(n_165), .B2(n_174), .Y(n_232) );
CKINVDCx6p67_ASAP7_75t_R g233 ( .A(n_219), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_191), .Y(n_235) );
INVx4_ASAP7_75t_SL g236 ( .A(n_191), .Y(n_236) );
OAI221xp5_ASAP7_75t_L g237 ( .A1(n_193), .A2(n_165), .B1(n_174), .B2(n_163), .C(n_168), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_219), .A2(n_174), .B1(n_183), .B2(n_188), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_195), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_213), .Y(n_240) );
OAI221xp5_ASAP7_75t_L g241 ( .A1(n_209), .A2(n_174), .B1(n_181), .B2(n_164), .C(n_188), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_219), .B(n_176), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
AO221x2_ASAP7_75t_L g245 ( .A1(n_199), .A2(n_171), .B1(n_101), .B2(n_91), .C(n_93), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_217), .A2(n_164), .B1(n_184), .B2(n_174), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_209), .B(n_171), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_202), .A2(n_184), .B1(n_180), .B2(n_187), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_245), .A2(n_203), .B1(n_222), .B2(n_202), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_230), .A2(n_199), .B(n_202), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_223), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_242), .B(n_202), .Y(n_252) );
BUFx5_ASAP7_75t_L g253 ( .A(n_242), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_228), .B(n_211), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_227), .A2(n_131), .A3(n_127), .B(n_129), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_235), .Y(n_256) );
AOI221xp5_ASAP7_75t_SL g257 ( .A1(n_241), .A2(n_173), .B1(n_221), .B2(n_151), .C(n_128), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_245), .A2(n_198), .B1(n_192), .B2(n_205), .Y(n_259) );
AOI31xp33_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_192), .A3(n_211), .B(n_208), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g261 ( .A1(n_232), .A2(n_198), .B1(n_205), .B2(n_173), .C(n_133), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_240), .B(n_220), .Y(n_262) );
OAI211xp5_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_101), .B(n_133), .C(n_93), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_235), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_236), .B(n_201), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_245), .A2(n_195), .B1(n_201), .B2(n_158), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_246), .A2(n_195), .B1(n_194), .B2(n_201), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_265), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_261), .A2(n_233), .B1(n_226), .B2(n_229), .Y(n_272) );
OAI21xp5_ASAP7_75t_SL g273 ( .A1(n_259), .A2(n_225), .B(n_239), .Y(n_273) );
AOI22xp33_ASAP7_75t_SL g274 ( .A1(n_268), .A2(n_224), .B1(n_229), .B2(n_225), .Y(n_274) );
INVxp67_ASAP7_75t_SL g275 ( .A(n_264), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_268), .B(n_224), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_261), .A2(n_239), .B1(n_237), .B2(n_226), .Y(n_277) );
OAI31xp33_ASAP7_75t_L g278 ( .A1(n_269), .A2(n_247), .A3(n_244), .B(n_243), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_265), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_251), .B(n_248), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_260), .A2(n_195), .B1(n_201), .B2(n_194), .Y(n_281) );
AOI31xp33_ASAP7_75t_L g282 ( .A1(n_259), .A2(n_107), .A3(n_87), .B(n_104), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_251), .B(n_149), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g284 ( .A1(n_260), .A2(n_208), .B1(n_212), .B2(n_220), .Y(n_284) );
OAI321xp33_ASAP7_75t_L g285 ( .A1(n_269), .A2(n_91), .A3(n_94), .B1(n_95), .B2(n_96), .C(n_99), .Y(n_285) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_263), .A2(n_107), .B(n_95), .C(n_96), .Y(n_286) );
NAND4xp25_ASAP7_75t_L g287 ( .A(n_249), .B(n_94), .C(n_99), .D(n_103), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_253), .B(n_109), .Y(n_288) );
INVx5_ASAP7_75t_L g289 ( .A(n_256), .Y(n_289) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_257), .A2(n_127), .B1(n_129), .B2(n_130), .C(n_104), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_267), .A2(n_208), .B1(n_212), .B2(n_220), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_292), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_253), .B1(n_252), .B2(n_264), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_292), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_280), .B(n_252), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_280), .B(n_255), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_255), .Y(n_299) );
AOI21xp5_ASAP7_75t_SL g300 ( .A1(n_281), .A2(n_266), .B(n_265), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g303 ( .A1(n_287), .A2(n_257), .B1(n_263), .B2(n_254), .C(n_264), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_282), .B(n_256), .Y(n_304) );
OR2x2_ASAP7_75t_SL g305 ( .A(n_278), .B(n_258), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_255), .Y(n_306) );
OAI221xp5_ASAP7_75t_SL g307 ( .A1(n_286), .A2(n_254), .B1(n_258), .B2(n_250), .C(n_270), .Y(n_307) );
AOI211x1_ASAP7_75t_SL g308 ( .A1(n_291), .A2(n_258), .B(n_250), .C(n_262), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_289), .B(n_255), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_289), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_289), .Y(n_311) );
NOR3xp33_ASAP7_75t_L g312 ( .A(n_274), .B(n_270), .C(n_256), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_277), .B(n_255), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_286), .A2(n_253), .B1(n_256), .B2(n_270), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_273), .A2(n_270), .B1(n_262), .B2(n_266), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AOI33xp33_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_130), .A3(n_153), .B1(n_154), .B2(n_140), .B3(n_141), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_276), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_296), .B(n_255), .Y(n_322) );
INVx3_ASAP7_75t_SL g323 ( .A(n_302), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_296), .B(n_255), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_295), .Y(n_326) );
NOR2x1_ASAP7_75t_L g327 ( .A(n_302), .B(n_266), .Y(n_327) );
NOR3xp33_ASAP7_75t_L g328 ( .A(n_304), .B(n_288), .C(n_157), .Y(n_328) );
NAND3xp33_ASAP7_75t_SL g329 ( .A(n_321), .B(n_153), .C(n_4), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_297), .B(n_253), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_297), .B(n_309), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_315), .B(n_253), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_321), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_316), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_300), .A2(n_266), .B(n_157), .C(n_5), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_314), .A2(n_253), .B1(n_236), .B2(n_212), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_253), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_306), .B(n_253), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_315), .B(n_253), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_299), .B(n_253), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_299), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_298), .B(n_236), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_315), .B(n_253), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_301), .B(n_1), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_306), .B(n_4), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_300), .A2(n_200), .B(n_206), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_301), .B(n_6), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_298), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_314), .B(n_7), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_8), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_302), .B(n_236), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_318), .A2(n_220), .B1(n_157), .B2(n_218), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_318), .A2(n_307), .B1(n_313), .B2(n_303), .C(n_317), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_305), .Y(n_361) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_319), .B(n_8), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_9), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_310), .B(n_9), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_334), .B(n_310), .Y(n_366) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_329), .B(n_317), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_333), .B(n_10), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_365), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_345), .B(n_308), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_294), .B1(n_312), .B2(n_308), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_352), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_354), .B(n_320), .C(n_157), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_331), .B(n_11), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_362), .A2(n_157), .B1(n_150), .B2(n_140), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_364), .B(n_11), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_364), .B(n_12), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_365), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_352), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_335), .A2(n_200), .B(n_206), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_345), .B(n_12), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_331), .B(n_13), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_341), .B(n_14), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_15), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_339), .A2(n_210), .B1(n_197), .B2(n_200), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_344), .B(n_16), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_325), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_360), .B(n_18), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_330), .B(n_19), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_349), .B(n_19), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_326), .B(n_150), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_330), .B(n_20), .Y(n_394) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_327), .B(n_150), .Y(n_395) );
AO22x2_ASAP7_75t_L g396 ( .A1(n_361), .A2(n_135), .B1(n_141), .B2(n_138), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_349), .B(n_135), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_323), .B(n_206), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_342), .B(n_21), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g401 ( .A(n_323), .B(n_357), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_361), .B(n_135), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_342), .B(n_23), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_361), .B(n_138), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g405 ( .A(n_360), .Y(n_405) );
OR2x6_ASAP7_75t_L g406 ( .A(n_327), .B(n_210), .Y(n_406) );
NAND2xp33_ASAP7_75t_SL g407 ( .A(n_357), .B(n_206), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_338), .Y(n_408) );
NAND2x1_ASAP7_75t_SL g409 ( .A(n_357), .B(n_143), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_322), .B(n_143), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_353), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_351), .B(n_24), .Y(n_412) );
NOR2x1p5_ASAP7_75t_L g413 ( .A(n_360), .B(n_143), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_407), .A2(n_358), .B(n_357), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_413), .B(n_346), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_408), .B(n_348), .Y(n_418) );
NOR4xp25_ASAP7_75t_L g419 ( .A(n_371), .B(n_359), .C(n_351), .D(n_356), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_379), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_411), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_389), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
XNOR2x1_ASAP7_75t_SL g424 ( .A(n_374), .B(n_363), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
NOR2xp33_ASAP7_75t_SL g426 ( .A(n_401), .B(n_346), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_405), .B(n_353), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_369), .B(n_355), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_378), .B(n_363), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_390), .B(n_346), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_381), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_370), .A2(n_356), .B(n_324), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_384), .B(n_332), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_385), .B(n_336), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
XOR2x2_ASAP7_75t_L g438 ( .A(n_368), .B(n_328), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_391), .B(n_337), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_390), .B(n_346), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_410), .B(n_347), .Y(n_441) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_371), .A2(n_339), .B(n_350), .C(n_343), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_383), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_386), .B(n_337), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_402), .Y(n_445) );
AOI211x1_ASAP7_75t_L g446 ( .A1(n_392), .A2(n_25), .B(n_28), .C(n_29), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_367), .A2(n_412), .B(n_375), .Y(n_447) );
OAI211xp5_ASAP7_75t_SL g448 ( .A1(n_376), .A2(n_340), .B(n_143), .C(n_182), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_388), .B(n_340), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g450 ( .A(n_377), .B(n_30), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_373), .A2(n_143), .B1(n_136), .B2(n_182), .C(n_179), .Y(n_452) );
XOR2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_394), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_401), .A2(n_182), .B1(n_179), .B2(n_175), .C1(n_162), .C2(n_218), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_400), .B(n_32), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_393), .Y(n_458) );
NOR4xp25_ASAP7_75t_L g459 ( .A(n_404), .B(n_179), .C(n_175), .D(n_162), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_396), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_398), .B(n_34), .Y(n_462) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_403), .B(n_35), .Y(n_463) );
NAND4xp75_ASAP7_75t_L g464 ( .A(n_382), .B(n_38), .C(n_40), .D(n_42), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_396), .B(n_46), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_387), .B(n_206), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_406), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_406), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_406), .B(n_50), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_371), .A2(n_197), .B1(n_210), .B2(n_180), .Y(n_471) );
XNOR2xp5_ASAP7_75t_L g472 ( .A(n_374), .B(n_52), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_372), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_372), .Y(n_474) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_413), .A2(n_197), .B(n_56), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_381), .Y(n_476) );
AO22x2_ASAP7_75t_L g477 ( .A1(n_408), .A2(n_54), .B1(n_58), .B2(n_60), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_370), .B(n_62), .Y(n_478) );
NAND2xp33_ASAP7_75t_R g479 ( .A(n_381), .B(n_63), .Y(n_479) );
AOI31xp33_ASAP7_75t_L g480 ( .A1(n_374), .A2(n_66), .A3(n_67), .B(n_69), .Y(n_480) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_374), .B(n_70), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_374), .Y(n_482) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_367), .A2(n_71), .B(n_72), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_453), .A2(n_475), .B(n_483), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_432), .A2(n_440), .B1(n_476), .B2(n_433), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_432), .A2(n_482), .B1(n_468), .B2(n_417), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_438), .A2(n_425), .B1(n_453), .B2(n_434), .Y(n_487) );
OAI211xp5_ASAP7_75t_SL g488 ( .A1(n_447), .A2(n_425), .B(n_471), .C(n_442), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_419), .A2(n_418), .B(n_428), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_479), .A2(n_431), .B1(n_426), .B2(n_438), .C(n_443), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_465), .B(n_461), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_480), .B(n_478), .C(n_448), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_478), .B(n_452), .C(n_466), .Y(n_493) );
AOI31xp33_ASAP7_75t_L g494 ( .A1(n_481), .A2(n_472), .A3(n_463), .B(n_470), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_469), .A2(n_415), .B1(n_424), .B2(n_431), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_450), .B(n_424), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_467), .A2(n_418), .B(n_437), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_427), .B(n_429), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_439), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_420), .Y(n_500) );
OAI211xp5_ASAP7_75t_SL g501 ( .A1(n_489), .A2(n_430), .B(n_455), .C(n_466), .Y(n_501) );
AOI221x1_ASAP7_75t_L g502 ( .A1(n_495), .A2(n_477), .B1(n_474), .B2(n_473), .C(n_414), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_484), .B(n_446), .C(n_451), .D(n_457), .Y(n_503) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_487), .B(n_437), .Y(n_504) );
AOI22x1_ASAP7_75t_L g505 ( .A1(n_497), .A2(n_477), .B1(n_455), .B2(n_436), .Y(n_505) );
AOI211xp5_ASAP7_75t_L g506 ( .A1(n_490), .A2(n_459), .B(n_460), .C(n_444), .Y(n_506) );
XNOR2x1_ASAP7_75t_L g507 ( .A(n_496), .B(n_477), .Y(n_507) );
OAI211xp5_ASAP7_75t_L g508 ( .A1(n_488), .A2(n_435), .B(n_449), .C(n_441), .Y(n_508) );
AOI211xp5_ASAP7_75t_L g509 ( .A1(n_486), .A2(n_454), .B(n_445), .C(n_458), .Y(n_509) );
AO22x2_ASAP7_75t_L g510 ( .A1(n_507), .A2(n_485), .B1(n_491), .B2(n_492), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_508), .Y(n_511) );
NOR2xp67_ASAP7_75t_L g512 ( .A(n_503), .B(n_499), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_506), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_502), .B(n_493), .C(n_494), .D(n_462), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_512), .A2(n_504), .B1(n_505), .B2(n_509), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_514), .B(n_501), .C(n_494), .Y(n_516) );
OAI222xp33_ASAP7_75t_L g517 ( .A1(n_511), .A2(n_498), .B1(n_500), .B2(n_456), .C1(n_423), .C2(n_416), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_516), .A2(n_510), .B1(n_513), .B2(n_464), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_515), .Y(n_519) );
AND3x4_ASAP7_75t_L g520 ( .A(n_518), .B(n_517), .C(n_421), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_520), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_521), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_522), .A2(n_519), .B(n_422), .Y(n_523) );
endmodule