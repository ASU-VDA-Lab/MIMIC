module fake_jpeg_15035_n_363 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_363);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_76),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_25),
.B(n_37),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_79),
.B1(n_27),
.B2(n_35),
.Y(n_109)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_35),
.B1(n_31),
.B2(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_29),
.Y(n_86)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_93),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_49),
.C(n_22),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_22),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_49),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_100),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_38),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_55),
.B1(n_47),
.B2(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_81),
.B1(n_74),
.B2(n_57),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_33),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_23),
.Y(n_141)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_24),
.B1(n_29),
.B2(n_32),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_110),
.B1(n_104),
.B2(n_93),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_18),
.B(n_13),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_70),
.B1(n_68),
.B2(n_62),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_116),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_120),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_87),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_123),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_135),
.C(n_19),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_31),
.B(n_21),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_128),
.B1(n_101),
.B2(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_68),
.B1(n_81),
.B2(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_129),
.B1(n_143),
.B2(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_24),
.B1(n_32),
.B2(n_36),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_37),
.B(n_1),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_106),
.B(n_102),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_39),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_54),
.B1(n_37),
.B2(n_36),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_88),
.B(n_92),
.C(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_36),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_150),
.B1(n_158),
.B2(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_99),
.B1(n_111),
.B2(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_111),
.B1(n_99),
.B2(n_89),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_164),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_90),
.B(n_37),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_174),
.B1(n_127),
.B2(n_137),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_163),
.B(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_116),
.B1(n_115),
.B2(n_105),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_126),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_122),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_182),
.C(n_190),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_122),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_192),
.Y(n_205)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_124),
.B1(n_135),
.B2(n_129),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_200),
.B1(n_146),
.B2(n_160),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_138),
.C(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_123),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_131),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_199),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_125),
.B1(n_118),
.B2(n_142),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_198),
.B1(n_202),
.B2(n_164),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_128),
.B1(n_144),
.B2(n_125),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_133),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_125),
.B1(n_118),
.B2(n_142),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_158),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_221),
.B1(n_186),
.B2(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_150),
.C(n_165),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_209),
.B(n_229),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_161),
.C(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_162),
.B1(n_159),
.B2(n_155),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_162),
.B1(n_161),
.B2(n_166),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_162),
.B(n_154),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_231),
.B(n_214),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_169),
.B1(n_167),
.B2(n_154),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_170),
.B1(n_157),
.B2(n_171),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_148),
.B1(n_134),
.B2(n_145),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_153),
.B(n_2),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_226),
.B(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_39),
.B(n_19),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_19),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_34),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_78),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_0),
.Y(n_256)
);

NAND2x1p5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_78),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_186),
.B(n_183),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_233),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_236),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_244),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_224),
.B(n_226),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_222),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_197),
.B1(n_187),
.B2(n_196),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_197),
.B(n_187),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_245),
.C(n_34),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_196),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_134),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_252),
.B1(n_2),
.B2(n_4),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_252)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_20),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_234),
.B(n_5),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_6),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_6),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_257),
.B(n_249),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_235),
.B1(n_257),
.B2(n_253),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_233),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_276),
.Y(n_292)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_246),
.C(n_243),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_20),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_238),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_280),
.C(n_281),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_253),
.B1(n_245),
.B2(n_250),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_259),
.B1(n_258),
.B2(n_266),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_277),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_296),
.B(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_250),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_260),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_310),
.C(n_313),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_312),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_297),
.B1(n_286),
.B2(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_274),
.B1(n_268),
.B2(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_299),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_292),
.A2(n_283),
.B1(n_284),
.B2(n_274),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_287),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_299),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_285),
.B(n_289),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_317),
.A2(n_304),
.B(n_310),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_325),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_311),
.A2(n_298),
.B1(n_262),
.B2(n_275),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_9),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_291),
.B(n_294),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_9),
.B(n_10),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_328),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_302),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_11),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_34),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_321),
.A2(n_313),
.B(n_10),
.Y(n_332)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_34),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_327),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_325),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_336),
.B(n_340),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_339),
.B(n_11),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_10),
.C(n_11),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_341),
.B(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_348),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_347),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_324),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_337),
.B(n_339),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_354),
.C(n_355),
.Y(n_356)
);

O2A1O1Ixp33_ASAP7_75t_SL g353 ( 
.A1(n_346),
.A2(n_334),
.B(n_319),
.C(n_330),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_12),
.B(n_16),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_322),
.Y(n_355)
);

NAND4xp25_ASAP7_75t_SL g357 ( 
.A(n_350),
.B(n_349),
.C(n_16),
.D(n_17),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_358),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_351),
.B(n_356),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_360),
.A2(n_351),
.B(n_20),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_20),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_20),
.B(n_34),
.Y(n_363)
);


endmodule