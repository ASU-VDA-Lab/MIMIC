module fake_jpeg_29265_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_7),
.B(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_50),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_27),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_51),
.B(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_65),
.Y(n_115)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_82),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_13),
.B1(n_11),
.B2(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_38),
.B1(n_20),
.B2(n_28),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_46),
.B1(n_37),
.B2(n_33),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_99),
.B(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_120),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_25),
.B(n_26),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_114),
.B(n_137),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_22),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_38),
.B1(n_20),
.B2(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_34),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_44),
.B(n_39),
.C(n_22),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_25),
.B1(n_41),
.B2(n_45),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_124),
.A2(n_127),
.B1(n_132),
.B2(n_29),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_34),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_79),
.A2(n_25),
.B1(n_41),
.B2(n_45),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_32),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_120),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_41),
.B1(n_45),
.B2(n_24),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_18),
.B(n_26),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_84),
.Y(n_169)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_146),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_163),
.Y(n_204)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_88),
.B1(n_78),
.B2(n_72),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_67),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_39),
.B1(n_44),
.B2(n_57),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_160),
.A2(n_164),
.B1(n_172),
.B2(n_177),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_26),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_162),
.B(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_123),
.A2(n_45),
.B1(n_18),
.B2(n_28),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_137),
.B1(n_102),
.B2(n_114),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_180),
.B(n_183),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_99),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_181),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_116),
.A2(n_18),
.B1(n_37),
.B2(n_49),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_100),
.B(n_75),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_188),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_77),
.B1(n_89),
.B2(n_82),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_136),
.A2(n_91),
.B1(n_74),
.B2(n_40),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_101),
.B(n_11),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_185),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_106),
.B(n_29),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_190),
.B1(n_151),
.B2(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_130),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_95),
.A2(n_29),
.B1(n_11),
.B2(n_2),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_140),
.B1(n_136),
.B2(n_94),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_195),
.A2(n_197),
.B1(n_207),
.B2(n_212),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_119),
.B1(n_94),
.B2(n_140),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_198),
.A2(n_183),
.B1(n_147),
.B2(n_182),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_110),
.C(n_105),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_190),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_205),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_144),
.A2(n_109),
.B1(n_95),
.B2(n_117),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_104),
.B(n_97),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_176),
.B(n_158),
.C(n_183),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_109),
.B1(n_93),
.B2(n_118),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_149),
.A2(n_118),
.B1(n_93),
.B2(n_133),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_178),
.B1(n_143),
.B2(n_184),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_104),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_131),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_151),
.A2(n_131),
.B1(n_133),
.B2(n_126),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_170),
.B1(n_154),
.B2(n_156),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_170),
.A2(n_97),
.B(n_126),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_174),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_233),
.A2(n_254),
.B1(n_260),
.B2(n_267),
.Y(n_277)
);

OR2x2_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_176),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_234),
.Y(n_281)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_236),
.A2(n_266),
.B(n_209),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_162),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_188),
.C(n_161),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_255),
.C(n_209),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_205),
.B(n_210),
.C(n_223),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_261),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_97),
.B1(n_113),
.B2(n_142),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_259),
.B1(n_265),
.B2(n_142),
.Y(n_271)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_249),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_246),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_176),
.B(n_179),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_251),
.Y(n_284)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_193),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_158),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_192),
.B(n_145),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_257),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_173),
.B1(n_166),
.B2(n_152),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_153),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx2_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_175),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_204),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_213),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_150),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_192),
.B(n_113),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_261),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_272),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_278),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_208),
.C(n_197),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_293),
.C(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_207),
.B(n_201),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_283),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_240),
.A2(n_198),
.B(n_220),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_246),
.A2(n_220),
.B1(n_219),
.B2(n_227),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_290),
.B1(n_292),
.B2(n_302),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_233),
.A2(n_195),
.B1(n_221),
.B2(n_212),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_230),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_267),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_228),
.B1(n_196),
.B2(n_206),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_219),
.C(n_227),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_191),
.C(n_206),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_191),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_262),
.A2(n_196),
.B1(n_232),
.B2(n_216),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_194),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_250),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_306),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_254),
.B1(n_247),
.B2(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_314),
.A2(n_326),
.B(n_289),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_244),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_328),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_251),
.B1(n_242),
.B2(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_323),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_284),
.B(n_279),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_321),
.B(n_322),
.Y(n_338)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_194),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_324),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_202),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_330),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_283),
.A2(n_236),
.B(n_234),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g328 ( 
.A(n_287),
.B(n_236),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_298),
.A2(n_236),
.B(n_216),
.C(n_249),
.D(n_199),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_331),
.A2(n_286),
.B1(n_241),
.B2(n_299),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_259),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_294),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_309),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_335),
.B(n_343),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_337),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_278),
.C(n_295),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_349),
.C(n_352),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_341),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_274),
.C(n_281),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_315),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_280),
.C(n_293),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_292),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_355),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_302),
.C(n_291),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_277),
.C(n_276),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_306),
.C(n_317),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_304),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_316),
.A2(n_286),
.B1(n_299),
.B2(n_199),
.Y(n_357)
);

AOI21xp33_ASAP7_75t_L g364 ( 
.A1(n_357),
.A2(n_305),
.B(n_332),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_308),
.B1(n_309),
.B2(n_307),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_359),
.A2(n_290),
.B1(n_347),
.B2(n_356),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_362),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_285),
.C(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_366),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_364),
.A2(n_350),
.B1(n_330),
.B2(n_324),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_334),
.B(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_370),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_326),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_378),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_323),
.C(n_329),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_377),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_320),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_277),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_353),
.C(n_352),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_382),
.C(n_383),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_358),
.B(n_336),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_385),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_348),
.C(n_355),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_348),
.C(n_343),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_370),
.B1(n_369),
.B2(n_372),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_335),
.B1(n_344),
.B2(n_347),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_359),
.A2(n_356),
.B(n_346),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_394),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_371),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_396),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_397),
.Y(n_408)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_391),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_404),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_402),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_373),
.C(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_379),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_394),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_376),
.C(n_375),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_407),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_341),
.C(n_313),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_393),
.Y(n_410)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_398),
.A2(n_311),
.B1(n_386),
.B2(n_388),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_385),
.B1(n_398),
.B2(n_403),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_399),
.B(n_383),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_417),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_406),
.A2(n_387),
.B(n_382),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_270),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_416),
.A2(n_403),
.B(n_404),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_419),
.A2(n_0),
.B(n_6),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_420),
.B1(n_424),
.B2(n_427),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_425),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_248),
.C(n_270),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_426),
.C(n_415),
.Y(n_429)
);

AO21x1_ASAP7_75t_L g424 ( 
.A1(n_410),
.A2(n_417),
.B(n_408),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_0),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_412),
.B(n_215),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_121),
.C(n_1),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_430),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_423),
.A2(n_426),
.B1(n_1),
.B2(n_4),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);

NOR3xp33_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_6),
.C(n_8),
.Y(n_435)
);

OAI321xp33_ASAP7_75t_L g438 ( 
.A1(n_435),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_428),
.C(n_436),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_429),
.C(n_433),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_438),
.C(n_8),
.Y(n_440)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_440),
.Y(n_441)
);


endmodule