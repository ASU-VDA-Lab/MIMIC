module fake_jpeg_26496_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_48),
.B1(n_19),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_33),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_26),
.B1(n_16),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_30),
.B1(n_27),
.B2(n_17),
.Y(n_64)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_60),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_67),
.Y(n_98)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_70),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_19),
.B1(n_18),
.B2(n_28),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_27),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_75),
.B(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_74),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_76),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_22),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_33),
.A3(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_101),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_57),
.C(n_36),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_100),
.C(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_44),
.B1(n_41),
.B2(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_117),
.B1(n_82),
.B2(n_88),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_42),
.C(n_39),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_39),
.Y(n_101)
);

OAI22x1_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_29),
.B1(n_22),
.B2(n_33),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_103),
.B1(n_110),
.B2(n_102),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_33),
.B(n_80),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_24),
.B1(n_98),
.B2(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_86),
.B1(n_89),
.B2(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_138),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_68),
.C(n_72),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_143),
.B1(n_139),
.B2(n_107),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_127),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_33),
.B(n_84),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_137),
.B(n_99),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_86),
.A3(n_73),
.B1(n_28),
.B2(n_24),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_117),
.A3(n_109),
.B1(n_114),
.B2(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_101),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_129),
.B1(n_14),
.B2(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_140),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_111),
.C(n_113),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_79),
.Y(n_138)
);

AOI21x1_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_79),
.B(n_58),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_109),
.B(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_0),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_0),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_2),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_94),
.B(n_118),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_147),
.B(n_151),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_153),
.B1(n_164),
.B2(n_2),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_167),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_2),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_110),
.B1(n_92),
.B2(n_102),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_100),
.B(n_93),
.C(n_103),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_159),
.B(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_124),
.B1(n_120),
.B2(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_173),
.B1(n_145),
.B2(n_141),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_114),
.B1(n_92),
.B2(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_134),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_170),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_125),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_168),
.C(n_159),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_157),
.Y(n_219)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_123),
.B(n_121),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_147),
.B(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_127),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_126),
.B1(n_123),
.B2(n_4),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_191),
.A2(n_182),
.B1(n_148),
.B2(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_14),
.C(n_12),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_162),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_146),
.C(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_8),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_14),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_214),
.B1(n_207),
.B2(n_211),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_218),
.C(n_202),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_158),
.B(n_172),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_160),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_160),
.C(n_157),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_232),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_179),
.C(n_189),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.C(n_231),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_177),
.C(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_184),
.B1(n_185),
.B2(n_199),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_188),
.C(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_187),
.C(n_178),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_191),
.C(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_195),
.C(n_191),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_211),
.B1(n_207),
.B2(n_206),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_152),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_152),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_175),
.C(n_167),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_204),
.CI(n_210),
.CON(n_245),
.SN(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_216),
.B(n_210),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_249),
.B(n_250),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_217),
.B(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

XOR2x1_ASAP7_75t_SL g253 ( 
.A(n_223),
.B(n_212),
.Y(n_253)
);

XOR2x1_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_233),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_225),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_257),
.B1(n_263),
.B2(n_245),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_217),
.B1(n_221),
.B2(n_208),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_242),
.B1(n_241),
.B2(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_224),
.C(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_262),
.C(n_251),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_212),
.C(n_10),
.Y(n_262)
);

FAx1_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_154),
.CI(n_5),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_154),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_251),
.C(n_244),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_255),
.B(n_241),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_248),
.B(n_263),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_260),
.C(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.C(n_11),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_270),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_268),
.B(n_11),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_276),
.B(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_287),
.B(n_11),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.C(n_283),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_292),
.B(n_3),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_284),
.B(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_3),
.C(n_5),
.Y(n_295)
);

OAI321xp33_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_293),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_6),
.Y(n_297)
);


endmodule