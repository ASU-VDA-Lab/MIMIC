module fake_netlist_1_1158_n_614 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_614);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_614;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_49), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_71), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_70), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_18), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_28), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_25), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_20), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_54), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_51), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_31), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_23), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_58), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_50), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_26), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_72), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_59), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_19), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_42), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_35), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_27), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_39), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_53), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_30), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_55), .Y(n_122) );
OR2x2_ASAP7_75t_L g123 ( .A(n_83), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
AND3x2_ASAP7_75t_L g126 ( .A(n_101), .B(n_0), .C(n_1), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_106), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
INVx6_ASAP7_75t_L g130 ( .A(n_113), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_89), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_115), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
NAND2xp33_ASAP7_75t_SL g139 ( .A(n_78), .B(n_2), .Y(n_139) );
INVx5_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
INVx2_ASAP7_75t_SL g149 ( .A(n_118), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_78), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_122), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_93), .B(n_2), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_121), .B(n_3), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_76), .B(n_3), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_77), .B(n_4), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_121), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_93), .B(n_5), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_79), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_82), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_92), .B(n_7), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_99), .B(n_7), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_128), .B(n_120), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
AND3x4_ASAP7_75t_L g167 ( .A(n_156), .B(n_102), .C(n_88), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_156), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_163), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_128), .A2(n_102), .B1(n_88), .B2(n_81), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_130), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_130), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_150), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_163), .B(n_117), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_124), .B(n_99), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_91), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_130), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_137), .A2(n_103), .B1(n_91), .B2(n_109), .Y(n_193) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_103), .B1(n_81), .B2(n_100), .Y(n_195) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_155), .B(n_98), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_129), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_159), .B(n_137), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_164), .A2(n_104), .B1(n_112), .B2(n_108), .Y(n_201) );
BUFx8_ASAP7_75t_SL g202 ( .A(n_164), .Y(n_202) );
BUFx10_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_125), .Y(n_204) );
INVx4_ASAP7_75t_SL g205 ( .A(n_154), .Y(n_205) );
INVxp67_ASAP7_75t_L g206 ( .A(n_127), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_133), .B(n_149), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_132), .B(n_114), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g210 ( .A(n_159), .B(n_105), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_140), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_145), .B(n_80), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_129), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_131), .B(n_96), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_134), .A2(n_97), .B1(n_94), .B2(n_11), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_131), .B(n_8), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_135), .B(n_8), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_189), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_192), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_186), .B(n_123), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_200), .A2(n_143), .B1(n_135), .B2(n_138), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_208), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_204), .B(n_123), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_169), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_186), .B(n_146), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_185), .B(n_144), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_220), .B(n_144), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_200), .Y(n_240) );
INVxp67_ASAP7_75t_SL g241 ( .A(n_206), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_172), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_165), .B(n_146), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_194), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_166), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_190), .B(n_138), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_165), .A2(n_139), .B1(n_158), .B2(n_157), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_174), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_190), .B(n_126), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_200), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_184), .B(n_143), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_165), .B(n_148), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_200), .Y(n_258) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_183), .B(n_133), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_202), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_207), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_209), .B(n_213), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_193), .A2(n_148), .B1(n_157), .B2(n_161), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_183), .B(n_162), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_197), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_202), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_197), .Y(n_268) );
INVx5_ASAP7_75t_L g269 ( .A(n_212), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_182), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_220), .A2(n_162), .B1(n_161), .B2(n_149), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_183), .B(n_162), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_195), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_196), .B(n_161), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_198), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_196), .B(n_140), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_221), .A2(n_152), .B1(n_147), .B2(n_141), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_198), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_270), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_242), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_242), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_270), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_242), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_270), .B(n_181), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_238), .Y(n_289) );
HAxp5_ASAP7_75t_L g290 ( .A(n_275), .B(n_167), .CON(n_290), .SN(n_290) );
BUFx4f_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_259), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g293 ( .A1(n_235), .A2(n_201), .B(n_173), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_223), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_238), .B(n_179), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_223), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_238), .Y(n_298) );
O2A1O1Ixp5_ASAP7_75t_L g299 ( .A1(n_264), .A2(n_168), .B(n_215), .C(n_217), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_230), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g302 ( .A1(n_275), .A2(n_167), .B1(n_216), .B2(n_210), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_236), .A2(n_210), .B1(n_180), .B2(n_187), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
AND2x6_ASAP7_75t_L g307 ( .A(n_237), .B(n_177), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_222), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_258), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_269), .Y(n_310) );
NAND2x1_ASAP7_75t_L g311 ( .A(n_279), .B(n_258), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_222), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_224), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_258), .B(n_203), .Y(n_315) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_229), .A2(n_187), .B1(n_180), .B2(n_178), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_233), .B(n_178), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_254), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_224), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_256), .A2(n_234), .B(n_248), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_236), .B(n_212), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_228), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_240), .B(n_177), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_245), .A2(n_136), .B1(n_147), .B2(n_152), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_228), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_278), .A2(n_171), .B(n_175), .C(n_170), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_248), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_269), .Y(n_331) );
OR2x2_ASAP7_75t_SL g332 ( .A(n_290), .B(n_261), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_302), .A2(n_225), .B1(n_252), .B2(n_241), .Y(n_333) );
BUFx2_ASAP7_75t_R g334 ( .A(n_292), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_321), .A2(n_236), .B1(n_282), .B2(n_229), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_330), .Y(n_336) );
NOR2xp33_ASAP7_75t_SL g337 ( .A(n_292), .B(n_259), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_293), .B(n_225), .Y(n_339) );
AO31x2_ASAP7_75t_L g340 ( .A1(n_314), .A2(n_147), .A3(n_141), .B(n_136), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_286), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_288), .B(n_225), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g344 ( .A1(n_290), .A2(n_271), .B1(n_267), .B2(n_252), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_286), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_286), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_288), .A2(n_252), .B1(n_247), .B2(n_233), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_288), .B(n_254), .Y(n_350) );
AND2x6_ASAP7_75t_L g351 ( .A(n_283), .B(n_260), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_290), .A2(n_267), .B1(n_249), .B2(n_257), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_291), .A2(n_250), .B1(n_263), .B2(n_249), .Y(n_353) );
NOR2xp67_ASAP7_75t_L g354 ( .A(n_283), .B(n_240), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_318), .B(n_274), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_308), .B(n_260), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_313), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_283), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_288), .A2(n_260), .B1(n_262), .B2(n_243), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_295), .A2(n_253), .B1(n_226), .B2(n_265), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_325), .A2(n_272), .B1(n_276), .B2(n_280), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_333), .A2(n_295), .B1(n_328), .B2(n_325), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_342), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_352), .A2(n_295), .B1(n_328), .B2(n_316), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_358), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_358), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_348), .A2(n_327), .B1(n_299), .B2(n_323), .C(n_305), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_337), .A2(n_291), .B1(n_313), .B2(n_320), .Y(n_370) );
A2O1A1Ixp33_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_320), .B(n_291), .C(n_295), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_346), .A2(n_319), .B1(n_307), .B2(n_298), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_336), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_351), .A2(n_319), .B1(n_307), .B2(n_298), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_353), .A2(n_304), .B1(n_301), .B2(n_300), .Y(n_376) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_351), .A2(n_307), .B1(n_312), .B2(n_309), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_297), .B1(n_303), .B2(n_294), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g379 ( .A1(n_339), .A2(n_300), .B1(n_304), .B2(n_301), .C1(n_306), .C2(n_297), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g380 ( .A1(n_356), .A2(n_141), .B(n_136), .C(n_152), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_334), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_306), .B1(n_296), .B2(n_303), .C(n_294), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_351), .A2(n_312), .B1(n_284), .B2(n_285), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_357), .B(n_296), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_336), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_350), .A2(n_317), .B1(n_312), .B2(n_289), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_338), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_351), .A2(n_307), .B1(n_312), .B2(n_309), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_329), .B1(n_287), .B2(n_284), .C(n_285), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_379), .A2(n_338), .B(n_355), .Y(n_390) );
AOI211xp5_ASAP7_75t_SL g391 ( .A1(n_370), .A2(n_341), .B(n_331), .C(n_354), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_381), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_366), .A2(n_361), .B(n_356), .C(n_355), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_371), .A2(n_341), .B(n_349), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_372), .A2(n_350), .B1(n_332), .B2(n_362), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_350), .B1(n_332), .B2(n_362), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_382), .A2(n_351), .B1(n_357), .B2(n_350), .Y(n_397) );
OAI222xp33_ASAP7_75t_L g398 ( .A1(n_373), .A2(n_341), .B1(n_359), .B2(n_349), .C1(n_347), .C2(n_345), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_374), .A2(n_351), .B1(n_359), .B2(n_354), .C1(n_287), .C2(n_345), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_376), .A2(n_347), .B1(n_317), .B2(n_312), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_378), .A2(n_311), .B(n_331), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
OAI31xp33_ASAP7_75t_L g403 ( .A1(n_369), .A2(n_324), .A3(n_322), .B(n_310), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_380), .A2(n_311), .B1(n_324), .B2(n_322), .C(n_310), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_387), .A2(n_351), .B1(n_326), .B2(n_307), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_387), .A2(n_142), .B1(n_151), .B2(n_140), .C(n_170), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_384), .Y(n_407) );
OAI321xp33_ASAP7_75t_L g408 ( .A1(n_386), .A2(n_142), .A3(n_151), .B1(n_219), .B2(n_171), .C(n_175), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_375), .A2(n_151), .B1(n_142), .B2(n_331), .C(n_289), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_307), .B1(n_326), .B2(n_142), .C1(n_151), .C2(n_140), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_199), .B(n_214), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_365), .A2(n_315), .B(n_309), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_385), .B(n_340), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_384), .A2(n_326), .B1(n_307), .B2(n_289), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_367), .B(n_340), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_367), .B(n_340), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_368), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_368), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_377), .A2(n_309), .B1(n_326), .B2(n_140), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_388), .A2(n_151), .B(n_140), .C(n_199), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_397), .A2(n_383), .B1(n_309), .B2(n_140), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_407), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_409), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_415), .A2(n_218), .B(n_214), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_419), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_417), .B(n_340), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_393), .A2(n_188), .A3(n_217), .B(n_218), .Y(n_429) );
OAI31xp33_ASAP7_75t_L g430 ( .A1(n_395), .A2(n_188), .A3(n_217), .B(n_13), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_390), .A2(n_188), .B(n_12), .C(n_13), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_402), .B(n_151), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_417), .B(n_10), .Y(n_434) );
OAI33xp33_ASAP7_75t_L g435 ( .A1(n_396), .A2(n_10), .A3(n_12), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_420), .B(n_14), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_418), .B(n_15), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
OAI33xp33_ASAP7_75t_L g440 ( .A1(n_400), .A2(n_16), .A3(n_281), .B1(n_277), .B2(n_268), .B3(n_266), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_405), .A2(n_309), .B1(n_269), .B2(n_219), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_398), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_413), .B(n_21), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_399), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_403), .B(n_22), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_403), .A2(n_219), .B1(n_203), .B2(n_273), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_410), .A2(n_219), .B1(n_203), .B2(n_273), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_394), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_401), .B(n_24), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_404), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_29), .Y(n_458) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_408), .B(n_273), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_219), .B1(n_273), .B2(n_231), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_392), .A2(n_273), .B1(n_246), .B2(n_244), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_422), .B(n_33), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_408), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_414), .B(n_37), .Y(n_464) );
INVx4_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_393), .A2(n_281), .A3(n_277), .B(n_268), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_427), .B(n_38), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_456), .A2(n_266), .B(n_255), .C(n_251), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_428), .B(n_40), .Y(n_469) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_465), .B(n_427), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_430), .B(n_255), .C(n_251), .D(n_44), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_465), .B(n_41), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_428), .B(n_43), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_434), .B(n_45), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_60), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_434), .B(n_62), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_453), .A2(n_246), .B1(n_244), .B2(n_239), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_428), .B(n_63), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_437), .B(n_65), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_465), .B(n_66), .Y(n_483) );
NAND3xp33_ASAP7_75t_SL g484 ( .A(n_429), .B(n_67), .C(n_73), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_438), .B(n_205), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_439), .B(n_205), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_424), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_205), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_435), .A2(n_231), .B1(n_239), .B2(n_244), .C(n_246), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_446), .B(n_205), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_438), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_446), .B(n_231), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_453), .B(n_231), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_447), .B(n_231), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_454), .B(n_239), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_452), .B(n_246), .Y(n_497) );
AND2x4_ASAP7_75t_SL g498 ( .A(n_448), .B(n_244), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_426), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_433), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_436), .B(n_442), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_426), .B(n_451), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_445), .B(n_451), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_455), .B(n_448), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_426), .B(n_445), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_445), .B(n_443), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_432), .B(n_466), .C(n_458), .D(n_449), .Y(n_509) );
OAI31xp67_ASAP7_75t_L g510 ( .A1(n_440), .A2(n_463), .A3(n_458), .B(n_423), .Y(n_510) );
NAND2x1_ASAP7_75t_SL g511 ( .A(n_452), .B(n_463), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_503), .B(n_464), .C(n_463), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g513 ( .A(n_474), .B(n_464), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_476), .B(n_462), .Y(n_515) );
AND4x1_ASAP7_75t_L g516 ( .A(n_470), .B(n_450), .C(n_460), .D(n_457), .Y(n_516) );
AND3x2_ASAP7_75t_L g517 ( .A(n_472), .B(n_452), .C(n_457), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_487), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_492), .A2(n_462), .B(n_441), .C(n_461), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_494), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_506), .B(n_487), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_469), .B(n_452), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_505), .B(n_459), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_496), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_509), .A2(n_459), .B1(n_471), .B2(n_498), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_483), .B(n_475), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_500), .B(n_493), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_479), .B(n_473), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_467), .B(n_497), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_493), .B(n_495), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_467), .Y(n_531) );
XNOR2x1_ASAP7_75t_L g532 ( .A(n_469), .B(n_481), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_507), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_473), .B(n_502), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_501), .B(n_502), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_501), .B(n_505), .Y(n_536) );
OR2x6_ASAP7_75t_L g537 ( .A(n_511), .B(n_497), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_477), .B(n_508), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_508), .B(n_498), .Y(n_539) );
AOI311xp33_ASAP7_75t_L g540 ( .A1(n_510), .A2(n_489), .A3(n_485), .B(n_511), .C(n_491), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_495), .B(n_491), .Y(n_541) );
NOR3xp33_ASAP7_75t_SL g542 ( .A(n_484), .B(n_510), .C(n_468), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_507), .B(n_490), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_490), .B(n_499), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_482), .B(n_499), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_536), .B(n_504), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_518), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_518), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_543), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_512), .A2(n_482), .B1(n_497), .B2(n_486), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_532), .A2(n_480), .B1(n_486), .B2(n_488), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_540), .B(n_488), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_536), .Y(n_554) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_537), .B(n_539), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_533), .B(n_530), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_533), .A2(n_521), .A3(n_515), .B1(n_529), .B2(n_534), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_527), .B(n_541), .Y(n_558) );
OAI211xp5_ASAP7_75t_L g559 ( .A1(n_525), .A2(n_519), .B(n_542), .C(n_531), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_544), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_513), .B(n_535), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_537), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_545), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_537), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_516), .B(n_517), .C(n_526), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_522), .B(n_528), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_520), .B(n_524), .Y(n_567) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_513), .B(n_532), .Y(n_568) );
NOR3x1_ASAP7_75t_L g569 ( .A(n_521), .B(n_503), .C(n_506), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_543), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_523), .B(n_538), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_521), .B(n_465), .Y(n_572) );
XNOR2xp5_ASAP7_75t_L g573 ( .A(n_532), .B(n_392), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_518), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_542), .A2(n_525), .B(n_512), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_512), .A2(n_525), .B(n_511), .C(n_503), .Y(n_578) );
XOR2xp5_ASAP7_75t_L g579 ( .A(n_513), .B(n_392), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g580 ( .A(n_532), .B(n_392), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_570), .Y(n_581) );
XOR2xp5_ASAP7_75t_L g582 ( .A(n_580), .B(n_573), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_554), .Y(n_583) );
AOI22x1_ASAP7_75t_L g584 ( .A1(n_579), .A2(n_580), .B1(n_573), .B2(n_576), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_563), .B(n_569), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_555), .A2(n_568), .B(n_553), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_561), .A2(n_565), .B1(n_548), .B2(n_574), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_559), .B(n_553), .C(n_578), .Y(n_588) );
NOR2xp33_ASAP7_75t_SL g589 ( .A(n_547), .B(n_572), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_550), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_550), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_579), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_546), .B(n_560), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_586), .A2(n_561), .B1(n_551), .B2(n_575), .Y(n_594) );
AOI211x1_ASAP7_75t_SL g595 ( .A1(n_588), .A2(n_584), .B(n_585), .C(n_587), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_582), .A2(n_568), .B1(n_551), .B2(n_564), .C(n_567), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_581), .Y(n_597) );
NOR4xp25_ASAP7_75t_L g598 ( .A(n_587), .B(n_564), .C(n_549), .D(n_577), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_592), .B(n_552), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_593), .A2(n_558), .B1(n_556), .B2(n_566), .Y(n_600) );
AOI22x1_ASAP7_75t_L g601 ( .A1(n_590), .A2(n_562), .B1(n_556), .B2(n_571), .Y(n_601) );
NAND4xp25_ASAP7_75t_L g602 ( .A(n_595), .B(n_589), .C(n_557), .D(n_562), .Y(n_602) );
NAND2x1p5_ASAP7_75t_SL g603 ( .A(n_601), .B(n_591), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_597), .B(n_583), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_599), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_604), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_605), .A2(n_594), .B1(n_596), .B2(n_598), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_603), .B(n_600), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_608), .Y(n_609) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_607), .B(n_602), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_609), .Y(n_611) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_611), .Y(n_612) );
XNOR2xp5_ASAP7_75t_L g613 ( .A(n_612), .B(n_610), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_613), .A2(n_610), .B(n_606), .Y(n_614) );
endmodule