module fake_jpeg_31186_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_11),
.Y(n_67)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_4),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_34),
.C(n_33),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_46),
.C(n_49),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_1),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_58),
.C(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_55),
.C(n_67),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_77),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_68),
.C(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_80),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_12),
.B(n_15),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_20),
.Y(n_88)
);


endmodule