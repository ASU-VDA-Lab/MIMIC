module fake_jpeg_23004_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_72),
.B1(n_82),
.B2(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_33),
.B1(n_25),
.B2(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_25),
.B1(n_34),
.B2(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_31),
.B1(n_24),
.B2(n_37),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_33),
.B1(n_37),
.B2(n_32),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_87),
.Y(n_125)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_50),
.B1(n_23),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_110),
.B1(n_63),
.B2(n_31),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_29),
.B1(n_35),
.B2(n_27),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_101),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_53),
.B(n_59),
.C(n_23),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_19),
.B(n_21),
.C(n_28),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_92),
.B1(n_111),
.B2(n_94),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_59),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_77),
.B1(n_79),
.B2(n_75),
.Y(n_154)
);

CKINVDCx9p33_ASAP7_75t_R g116 ( 
.A(n_54),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_28),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_55),
.B(n_24),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_106),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_67),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_126),
.A2(n_141),
.B(n_130),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_143),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_105),
.B1(n_95),
.B2(n_122),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_19),
.B(n_22),
.Y(n_184)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_39),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_63),
.B1(n_77),
.B2(n_76),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_146),
.B1(n_97),
.B2(n_100),
.Y(n_189)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_17),
.B1(n_27),
.B2(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_39),
.C(n_41),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_150),
.C(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_46),
.B1(n_66),
.B2(n_58),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_151),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_46),
.C(n_44),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_74),
.C(n_35),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_111),
.B1(n_95),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_164),
.B1(n_168),
.B2(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_161),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_174),
.Y(n_195)
);

XOR2x1_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_102),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_184),
.B(n_129),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_101),
.B1(n_120),
.B2(n_122),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_179),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_148),
.C(n_153),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_11),
.C(n_16),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_102),
.B1(n_120),
.B2(n_109),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_173),
.A2(n_186),
.B1(n_155),
.B2(n_139),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_87),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_98),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_181),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_123),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_87),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_113),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_116),
.C(n_28),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_136),
.B1(n_151),
.B2(n_150),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_30),
.B(n_19),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_132),
.A2(n_19),
.B1(n_114),
.B2(n_109),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_192),
.B1(n_129),
.B2(n_123),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_197),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_138),
.B(n_140),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_214),
.B(n_179),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_134),
.B1(n_156),
.B2(n_158),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_215),
.B1(n_214),
.B2(n_210),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_218),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_186),
.B1(n_160),
.B2(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_98),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_217),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_219),
.C(n_2),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_166),
.B1(n_180),
.B2(n_168),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_22),
.B(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_100),
.C(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_162),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_22),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_170),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_0),
.B(n_2),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_218),
.B(n_200),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_230),
.B(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_162),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_189),
.B1(n_191),
.B2(n_169),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_196),
.A2(n_191),
.B1(n_165),
.B2(n_181),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_178),
.B1(n_165),
.B2(n_181),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_221),
.B1(n_202),
.B2(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_161),
.B1(n_171),
.B2(n_183),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_203),
.B1(n_197),
.B2(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_223),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_246),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_13),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_213),
.C(n_219),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_226),
.B(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_229),
.B1(n_248),
.B2(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_265),
.C(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_228),
.B(n_217),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_257),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_200),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_204),
.B1(n_199),
.B2(n_196),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_262),
.B1(n_266),
.B2(n_267),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_199),
.B1(n_201),
.B2(n_194),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_2),
.C(n_3),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_225),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_8),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_250),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_247),
.C(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_283),
.C(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_282),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_225),
.B1(n_233),
.B2(n_224),
.Y(n_278)
);

AOI21x1_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_231),
.B(n_232),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_254),
.B1(n_263),
.B2(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_245),
.C(n_231),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_246),
.C(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_286),
.B1(n_265),
.B2(n_254),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_268),
.C(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_277),
.C(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_284),
.B1(n_10),
.B2(n_12),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_291),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_250),
.C(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_258),
.C(n_5),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_298),
.B(n_286),
.Y(n_303)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_272),
.B1(n_278),
.B2(n_282),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_272),
.B1(n_270),
.B2(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_297),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_274),
.B(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_298),
.C(n_288),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_298),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_309),
.B1(n_289),
.B2(n_287),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_280),
.B1(n_285),
.B2(n_270),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_292),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_287),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_308),
.B(n_301),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_326),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_311),
.B(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_322),
.B1(n_302),
.B2(n_321),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_303),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_327),
.B1(n_328),
.B2(n_10),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_13),
.B(n_6),
.Y(n_331)
);

AOI32xp33_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_5),
.A3(n_7),
.B1(n_13),
.B2(n_298),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_7),
.Y(n_333)
);


endmodule