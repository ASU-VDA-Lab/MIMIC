module fake_jpeg_26276_n_273 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_64),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_21),
.CON(n_52),
.SN(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_17),
.B(n_22),
.C(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_60),
.B1(n_65),
.B2(n_27),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_24),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_24),
.B1(n_19),
.B2(n_31),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_19),
.B1(n_31),
.B2(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_45),
.B1(n_47),
.B2(n_53),
.Y(n_93)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_43),
.B(n_27),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_80),
.B(n_84),
.Y(n_115)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_44),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_90),
.B1(n_63),
.B2(n_45),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_38),
.B(n_44),
.C(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_63),
.B1(n_45),
.B2(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_89),
.Y(n_92)
);

NOR4xp25_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_59),
.C(n_60),
.D(n_56),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_76),
.A3(n_82),
.B1(n_59),
.B2(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_115),
.B(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_114),
.B1(n_92),
.B2(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_102),
.B1(n_51),
.B2(n_70),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_101),
.Y(n_131)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_49),
.C(n_58),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_105),
.C(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_110),
.Y(n_140)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_49),
.C(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_75),
.B1(n_79),
.B2(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_113),
.B1(n_91),
.B2(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_117),
.A2(n_128),
.B1(n_135),
.B2(n_139),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_136),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_28),
.B(n_34),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_95),
.B1(n_102),
.B2(n_99),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_125),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_4),
.B(n_6),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_70),
.B1(n_68),
.B2(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_34),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_44),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_38),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_19),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_44),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_104),
.C(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_69),
.B1(n_74),
.B2(n_73),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_148),
.B(n_158),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_132),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_146),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_38),
.B(n_98),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_28),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_155),
.Y(n_172)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_157),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_1),
.C(n_2),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_121),
.C(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_160),
.B(n_164),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_3),
.B(n_4),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_3),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_7),
.B(n_8),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_117),
.B1(n_135),
.B2(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_182),
.B1(n_151),
.B2(n_166),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_177),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_168),
.C(n_147),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_185),
.C(n_192),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_147),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_181),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

BUFx12f_ASAP7_75t_SL g179 ( 
.A(n_164),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_191),
.B(n_141),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_155),
.B1(n_157),
.B2(n_159),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_132),
.C(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_120),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_151),
.B1(n_158),
.B2(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_156),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_142),
.C(n_138),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_183),
.B(n_187),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_15),
.C(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_181),
.C(n_170),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_7),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_187),
.B1(n_171),
.B2(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_207),
.Y(n_217)
);

BUFx4f_ASAP7_75t_SL g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_203),
.B(n_210),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_222),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_227),
.Y(n_229)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_177),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_9),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_177),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_202),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_235),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_233),
.B(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_194),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_237),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_212),
.B(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_200),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_205),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_232),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_224),
.C(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_248),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_237),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_206),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_247),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_209),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_214),
.C(n_216),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_228),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_214),
.C(n_230),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_197),
.B(n_215),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_218),
.B(n_193),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

OA21x2_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_246),
.B(n_202),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_251),
.B(n_261),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_246),
.C(n_11),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_10),
.B(n_11),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_266),
.B(n_268),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_260),
.A3(n_263),
.B1(n_13),
.B2(n_14),
.C1(n_10),
.C2(n_12),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_13),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_270),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_269),
.B1(n_13),
.B2(n_14),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_272),
.Y(n_273)
);


endmodule