module fake_jpeg_2243_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_66),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_48),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_85),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_84),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_51),
.B1(n_63),
.B2(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_51),
.B1(n_63),
.B2(n_62),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_71),
.B1(n_69),
.B2(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_94),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_48),
.B1(n_67),
.B2(n_59),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_25),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_78),
.A3(n_58),
.B1(n_56),
.B2(n_5),
.Y(n_116)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_89),
.B(n_96),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_21),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_98),
.B1(n_87),
.B2(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_78),
.B1(n_56),
.B2(n_27),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_78),
.C(n_56),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_113),
.Y(n_135)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_2),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_20),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_35),
.B1(n_42),
.B2(n_41),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_23),
.B(n_47),
.C(n_46),
.D(n_45),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_112),
.B(n_34),
.Y(n_146)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_78),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_137),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_109),
.B(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_104),
.B(n_12),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_31),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_122),
.B1(n_120),
.B2(n_119),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_123),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_154),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_33),
.Y(n_154)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_126),
.A3(n_36),
.B1(n_29),
.B2(n_43),
.C1(n_39),
.C2(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_147),
.B1(n_143),
.B2(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_38),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_125),
.B1(n_141),
.B2(n_124),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_153),
.B1(n_148),
.B2(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_167),
.B(n_171),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_169),
.B1(n_161),
.B2(n_159),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_165),
.C(n_154),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.C(n_168),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_170),
.B(n_160),
.C(n_169),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_166),
.B(n_37),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_30),
.B1(n_15),
.B2(n_16),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_14),
.C(n_17),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_18),
.C(n_14),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_17),
.Y(n_184)
);


endmodule