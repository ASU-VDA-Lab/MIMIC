module real_aes_14593_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_898;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_633;
wire n_926;
wire n_679;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g687 ( .A(n_0), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_1), .Y(n_576) );
INVx1_ASAP7_75t_L g132 ( .A(n_2), .Y(n_132) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_2), .A2(n_50), .B(n_134), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_3), .B(n_245), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_4), .B(n_241), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_5), .B(n_200), .Y(n_199) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_6), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g667 ( .A(n_7), .B(n_228), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_8), .A2(n_93), .B1(n_922), .B2(n_923), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_8), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_9), .B(n_259), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_10), .B(n_148), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_11), .B(n_173), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_12), .Y(n_129) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_13), .B(n_227), .Y(n_644) );
BUFx3_ASAP7_75t_L g150 ( .A(n_14), .Y(n_150) );
INVx1_ASAP7_75t_L g167 ( .A(n_14), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_15), .A2(n_181), .B(n_182), .C(n_184), .Y(n_180) );
BUFx10_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_17), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_18), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_112) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_18), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_19), .B(n_259), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_20), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_21), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_22), .B(n_247), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_23), .A2(n_164), .B(n_168), .C(n_171), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_24), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_25), .B(n_269), .C(n_700), .Y(n_702) );
AND2x2_ASAP7_75t_L g237 ( .A(n_26), .B(n_236), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_27), .A2(n_919), .B1(n_925), .B2(n_926), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_27), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_28), .B(n_200), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_29), .B(n_227), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_30), .A2(n_75), .B1(n_151), .B2(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
INVx1_ASAP7_75t_L g204 ( .A(n_32), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_33), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_34), .B(n_151), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_35), .A2(n_105), .B1(n_935), .B2(n_946), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_36), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_37), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g532 ( .A(n_38), .Y(n_532) );
AND3x2_ASAP7_75t_L g933 ( .A(n_38), .B(n_550), .C(n_551), .Y(n_933) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_39), .B(n_165), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_40), .B(n_181), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_41), .B(n_227), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_42), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_43), .B(n_189), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_44), .Y(n_183) );
AND2x4_ASAP7_75t_L g139 ( .A(n_45), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_46), .B(n_227), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_47), .B(n_236), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_48), .B(n_227), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_49), .A2(n_87), .B1(n_148), .B2(n_151), .Y(n_147) );
INVx1_ASAP7_75t_L g131 ( .A(n_50), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_51), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_52), .A2(n_662), .B(n_686), .C(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g134 ( .A(n_53), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_54), .B(n_227), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_55), .A2(n_920), .B1(n_921), .B2(n_924), .Y(n_919) );
INVxp67_ASAP7_75t_SL g924 ( .A(n_55), .Y(n_924) );
AND2x4_ASAP7_75t_L g944 ( .A(n_56), .B(n_945), .Y(n_944) );
OAI22xp33_ASAP7_75t_L g118 ( .A1(n_57), .A2(n_100), .B1(n_119), .B2(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_57), .Y(n_120) );
INVx3_ASAP7_75t_L g628 ( .A(n_58), .Y(n_628) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_59), .B(n_77), .Y(n_533) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_59), .Y(n_939) );
AND2x2_ASAP7_75t_L g311 ( .A(n_60), .B(n_228), .Y(n_311) );
INVx1_ASAP7_75t_L g945 ( .A(n_61), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_62), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_63), .B(n_604), .Y(n_609) );
NAND2x1_ASAP7_75t_L g274 ( .A(n_64), .B(n_181), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_65), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g640 ( .A(n_66), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_67), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_68), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g530 ( .A(n_69), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_70), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_71), .B(n_148), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_72), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_73), .B(n_269), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_74), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_76), .B(n_165), .Y(n_310) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_77), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_78), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_79), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_80), .B(n_259), .Y(n_270) );
NAND2xp33_ASAP7_75t_SL g197 ( .A(n_81), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_82), .B(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g680 ( .A(n_83), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_84), .B(n_192), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_85), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_86), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
BUFx3_ASAP7_75t_L g173 ( .A(n_88), .Y(n_173) );
INVx1_ASAP7_75t_L g195 ( .A(n_88), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_89), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_90), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_91), .B(n_148), .Y(n_574) );
INVx1_ASAP7_75t_L g626 ( .A(n_92), .Y(n_626) );
INVx1_ASAP7_75t_L g923 ( .A(n_93), .Y(n_923) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_94), .B(n_257), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_95), .B(n_228), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g218 ( .A(n_96), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_97), .B(n_608), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_98), .Y(n_622) );
INVx1_ASAP7_75t_L g618 ( .A(n_99), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_100), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_101), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_102), .B(n_189), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_103), .B(n_604), .Y(n_603) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_545), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx3_ASAP7_75t_L g552 ( .A(n_109), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_109), .B(n_933), .Y(n_932) );
OAI21xp5_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_116), .B(n_534), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_112), .B(n_536), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_113), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_525), .Y(n_116) );
INVx1_ASAP7_75t_L g540 ( .A(n_117), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
AOI22x1_ASAP7_75t_L g555 ( .A1(n_121), .A2(n_556), .B1(n_561), .B2(n_915), .Y(n_555) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_429), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_338), .C(n_402), .Y(n_122) );
OAI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_230), .B1(n_277), .B2(n_288), .C(n_293), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_158), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g350 ( .A(n_126), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g365 ( .A(n_126), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g438 ( .A(n_126), .B(n_185), .Y(n_438) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g285 ( .A(n_127), .Y(n_285) );
INVx1_ASAP7_75t_L g317 ( .A(n_127), .Y(n_317) );
AND2x2_ASAP7_75t_L g336 ( .A(n_127), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g363 ( .A(n_127), .B(n_353), .Y(n_363) );
INVxp67_ASAP7_75t_L g378 ( .A(n_127), .Y(n_378) );
AND2x2_ASAP7_75t_L g401 ( .A(n_127), .B(n_212), .Y(n_401) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_127), .Y(n_428) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_135), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_130), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_133), .Y(n_130) );
AOI21x1_ASAP7_75t_L g146 ( .A1(n_131), .A2(n_132), .B(n_133), .Y(n_146) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_147), .B1(n_153), .B2(n_155), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .C(n_145), .Y(n_136) );
NAND3xp33_ASAP7_75t_L g153 ( .A(n_137), .B(n_145), .C(n_154), .Y(n_153) );
BUFx2_ASAP7_75t_L g666 ( .A(n_137), .Y(n_666) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_138), .A2(n_178), .B(n_684), .Y(n_689) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
BUFx6f_ASAP7_75t_SL g210 ( .A(n_139), .Y(n_210) );
INVx1_ASAP7_75t_L g301 ( .A(n_139), .Y(n_301) );
INVx3_ASAP7_75t_L g620 ( .A(n_139), .Y(n_620) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_142), .B(n_620), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_142), .B(n_620), .C(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_145), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_145), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
INVx2_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
INVx2_ASAP7_75t_L g247 ( .A(n_149), .Y(n_247) );
INVx2_ASAP7_75t_L g578 ( .A(n_149), .Y(n_578) );
INVx3_ASAP7_75t_L g654 ( .A(n_149), .Y(n_654) );
INVx3_ASAP7_75t_L g679 ( .A(n_149), .Y(n_679) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g152 ( .A(n_150), .Y(n_152) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_151), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g269 ( .A(n_152), .Y(n_269) );
O2A1O1Ixp5_ASAP7_75t_L g271 ( .A1(n_154), .A2(n_272), .B(n_273), .C(n_274), .Y(n_271) );
INVx2_ASAP7_75t_L g305 ( .A(n_154), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_154), .A2(n_588), .B(n_589), .Y(n_587) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
INVx2_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
INVx2_ASAP7_75t_L g309 ( .A(n_157), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_158), .A2(n_407), .B(n_411), .Y(n_406) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_185), .Y(n_158) );
AND2x2_ASAP7_75t_L g508 ( .A(n_159), .B(n_401), .Y(n_508) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g281 ( .A(n_161), .Y(n_281) );
INVx1_ASAP7_75t_L g319 ( .A(n_161), .Y(n_319) );
AND2x2_ASAP7_75t_L g347 ( .A(n_161), .B(n_284), .Y(n_347) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_161), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_162), .B(n_179), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_162), .B(n_179), .Y(n_337) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_174), .B(n_177), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_164), .A2(n_604), .B1(n_625), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_165), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g593 ( .A(n_165), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_165), .B(n_618), .Y(n_617) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g170 ( .A(n_166), .Y(n_170) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_167), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx2_ASAP7_75t_L g181 ( .A(n_170), .Y(n_181) );
INVx2_ASAP7_75t_L g241 ( .A(n_170), .Y(n_241) );
INVx2_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_170), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_171), .A2(n_222), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_172), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
AOI211x1_ASAP7_75t_L g238 ( .A1(n_173), .A2(n_237), .B(n_239), .C(n_243), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_173), .B(n_620), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_173), .B(n_620), .C(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g179 ( .A(n_174), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g611 ( .A(n_175), .Y(n_611) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
INVx1_ASAP7_75t_L g580 ( .A(n_176), .Y(n_580) );
INVxp67_ASAP7_75t_L g665 ( .A(n_178), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_184), .A2(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g664 ( .A(n_184), .Y(n_664) );
AND2x2_ASAP7_75t_L g335 ( .A(n_185), .B(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g524 ( .A(n_185), .Y(n_524) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_211), .Y(n_185) );
INVx2_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
AND2x2_ASAP7_75t_L g318 ( .A(n_186), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g329 ( .A(n_186), .Y(n_329) );
OR2x2_ASAP7_75t_L g367 ( .A(n_186), .B(n_337), .Y(n_367) );
AND2x2_ASAP7_75t_L g379 ( .A(n_186), .B(n_337), .Y(n_379) );
AND2x2_ASAP7_75t_L g449 ( .A(n_186), .B(n_212), .Y(n_449) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_196), .A3(n_202), .B(n_207), .Y(n_186) );
AO21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B(n_193), .Y(n_187) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g198 ( .A(n_190), .Y(n_198) );
INVx1_ASAP7_75t_L g219 ( .A(n_190), .Y(n_219) );
INVx2_ASAP7_75t_L g245 ( .A(n_190), .Y(n_245) );
INVx2_ASAP7_75t_L g273 ( .A(n_192), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_193), .A2(n_244), .B(n_246), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_193), .A2(n_256), .B(n_258), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_193), .A2(n_268), .B(n_270), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_193), .A2(n_573), .B(n_574), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_193), .A2(n_591), .B(n_592), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_193), .A2(n_642), .B(n_643), .Y(n_641) );
BUFx10_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g700 ( .A(n_194), .Y(n_700) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx3_ASAP7_75t_L g658 ( .A(n_195), .Y(n_658) );
AO21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_199), .B(n_201), .Y(n_196) );
INVx2_ASAP7_75t_L g259 ( .A(n_198), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_201), .A2(n_253), .B(n_254), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_201), .A2(n_576), .B(n_577), .C(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_203), .A2(n_208), .B(n_210), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVxp33_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx2_ASAP7_75t_L g209 ( .A(n_206), .Y(n_209) );
INVx1_ASAP7_75t_L g229 ( .A(n_206), .Y(n_229) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_206), .Y(n_236) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx3_ASAP7_75t_L g213 ( .A(n_209), .Y(n_213) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_210), .A2(n_215), .B(n_221), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_210), .A2(n_235), .B(n_237), .Y(n_234) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_210), .A2(n_252), .B(n_255), .Y(n_251) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_210), .A2(n_587), .B(n_590), .Y(n_586) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_210), .A2(n_635), .B(n_641), .Y(n_634) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g287 ( .A(n_212), .Y(n_287) );
INVx1_ASAP7_75t_L g353 ( .A(n_212), .Y(n_353) );
AND2x2_ASAP7_75t_L g375 ( .A(n_212), .B(n_285), .Y(n_375) );
AND2x2_ASAP7_75t_L g458 ( .A(n_212), .B(n_352), .Y(n_458) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_226), .Y(n_212) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_213), .A2(n_571), .B(n_581), .Y(n_570) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_213), .A2(n_634), .B(n_644), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_218), .B(n_220), .Y(n_215) );
INVx2_ASAP7_75t_L g604 ( .A(n_217), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_217), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g608 ( .A(n_219), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_220), .A2(n_308), .B(n_310), .Y(n_307) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_227), .Y(n_693) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_248), .Y(n_230) );
AND2x2_ASAP7_75t_L g381 ( .A(n_231), .B(n_372), .Y(n_381) );
OR2x2_ASAP7_75t_L g397 ( .A(n_231), .B(n_332), .Y(n_397) );
INVx2_ASAP7_75t_L g409 ( .A(n_231), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_231), .B(n_345), .Y(n_412) );
AND2x2_ASAP7_75t_L g509 ( .A(n_231), .B(n_424), .Y(n_509) );
BUFx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g289 ( .A(n_232), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g419 ( .A(n_232), .B(n_324), .Y(n_419) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g312 ( .A(n_233), .B(n_250), .Y(n_312) );
INVx2_ASAP7_75t_L g343 ( .A(n_233), .Y(n_343) );
BUFx2_ASAP7_75t_L g370 ( .A(n_233), .Y(n_370) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_233), .Y(n_387) );
INVx1_ASAP7_75t_L g394 ( .A(n_233), .Y(n_394) );
AND2x2_ASAP7_75t_L g453 ( .A(n_233), .B(n_396), .Y(n_453) );
INVx1_ASAP7_75t_L g514 ( .A(n_233), .Y(n_514) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_238), .Y(n_233) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
NOR2xp67_ASAP7_75t_SL g300 ( .A(n_236), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g738 ( .A(n_236), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_242), .Y(n_239) );
INVx2_ASAP7_75t_L g662 ( .A(n_245), .Y(n_662) );
INVxp67_ASAP7_75t_L g636 ( .A(n_247), .Y(n_636) );
INVxp67_ASAP7_75t_L g660 ( .A(n_247), .Y(n_660) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_263), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_249), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g323 ( .A(n_250), .B(n_324), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_260), .B(n_262), .Y(n_250) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_251), .A2(n_260), .B(n_262), .Y(n_292) );
INVx2_ASAP7_75t_L g656 ( .A(n_257), .Y(n_656) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_260), .A2(n_266), .B(n_276), .Y(n_265) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_260), .A2(n_586), .B(n_594), .Y(n_585) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_260), .A2(n_651), .B(n_723), .Y(n_722) );
OAI21x1_ASAP7_75t_L g728 ( .A1(n_260), .A2(n_586), .B(n_594), .Y(n_728) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2x1_ASAP7_75t_SL g610 ( .A(n_261), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g479 ( .A(n_263), .Y(n_479) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g396 ( .A(n_264), .Y(n_396) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
INVx1_ASAP7_75t_L g359 ( .A(n_265), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_271), .B(n_275), .Y(n_266) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_277), .A2(n_403), .B(n_406), .C(n_413), .Y(n_402) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_281), .Y(n_326) );
AND2x2_ASAP7_75t_L g445 ( .A(n_281), .B(n_375), .Y(n_445) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
AND2x2_ASAP7_75t_L g355 ( .A(n_283), .B(n_351), .Y(n_355) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g416 ( .A(n_284), .Y(n_416) );
INVx2_ASAP7_75t_L g389 ( .A(n_286), .Y(n_389) );
BUFx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_287), .B(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_287), .Y(n_491) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g345 ( .A(n_290), .B(n_322), .Y(n_345) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g358 ( .A(n_291), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g372 ( .A(n_291), .B(n_298), .Y(n_372) );
AND2x2_ASAP7_75t_L g495 ( .A(n_291), .B(n_322), .Y(n_495) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_298), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_313), .B1(n_320), .B2(n_325), .C(n_330), .Y(n_293) );
AOI222xp33_ASAP7_75t_L g487 ( .A1(n_294), .A2(n_425), .B1(n_488), .B2(n_493), .C1(n_496), .C2(n_497), .Y(n_487) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_312), .Y(n_295) );
INVx4_ASAP7_75t_R g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_297), .B(n_388), .Y(n_405) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_298), .B(n_322), .Y(n_332) );
AND2x4_ASAP7_75t_L g393 ( .A(n_298), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_306), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_300), .A2(n_307), .B(n_311), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_305), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_305), .A2(n_607), .B(n_609), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_309), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_315), .B(n_501), .C(n_504), .Y(n_500) );
OR2x2_ASAP7_75t_L g516 ( .A(n_315), .B(n_504), .Y(n_516) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_316), .A2(n_386), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g450 ( .A(n_317), .B(n_337), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_318), .B(n_401), .Y(n_421) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
OR2x2_ASAP7_75t_L g464 ( .A(n_321), .B(n_333), .Y(n_464) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g442 ( .A(n_323), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_323), .B(n_369), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_323), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_323), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_323), .B(n_479), .Y(n_507) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_324), .B(n_343), .Y(n_342) );
NOR2x1p5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_329), .B(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_334), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g424 ( .A(n_333), .Y(n_424) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_333), .B(n_513), .Y(n_521) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g456 ( .A(n_336), .B(n_449), .Y(n_456) );
INVx2_ASAP7_75t_L g352 ( .A(n_337), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_339), .B(n_382), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_360), .C(n_373), .Y(n_339) );
OAI322xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .A3(n_346), .B1(n_348), .B2(n_349), .C1(n_354), .C2(n_356), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g480 ( .A(n_342), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_344), .A2(n_455), .B1(n_457), .B2(n_459), .Y(n_454) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_345), .B(n_393), .Y(n_498) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_SL g362 ( .A(n_347), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g443 ( .A(n_347), .B(n_401), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_347), .B(n_378), .Y(n_519) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g475 ( .A(n_350), .B(n_416), .Y(n_475) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_356), .A2(n_393), .A3(n_414), .B1(n_417), .B2(n_420), .C1(n_422), .C2(n_425), .Y(n_413) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp33_ASAP7_75t_L g418 ( .A(n_357), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g410 ( .A(n_358), .Y(n_410) );
OR2x2_ASAP7_75t_L g433 ( .A(n_358), .B(n_419), .Y(n_433) );
BUFx2_ASAP7_75t_L g388 ( .A(n_359), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_368), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_391), .B1(n_397), .B2(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g483 ( .A(n_363), .Y(n_483) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g386 ( .A(n_367), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g426 ( .A(n_367), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g466 ( .A(n_367), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g482 ( .A(n_367), .B(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_370), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g441 ( .A(n_370), .Y(n_441) );
OR2x2_ASAP7_75t_L g459 ( .A(n_371), .B(n_395), .Y(n_459) );
OR2x2_ASAP7_75t_L g485 ( .A(n_371), .B(n_479), .Y(n_485) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B(n_380), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_375), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g504 ( .A(n_379), .Y(n_504) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_389), .B(n_390), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_393), .B(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_394), .Y(n_470) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g513 ( .A(n_396), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_398), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_401), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g467 ( .A(n_401), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_403), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g486 ( .A(n_409), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_409), .B(n_424), .C(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g523 ( .A(n_427), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR3xp33_ASAP7_75t_SL g429 ( .A(n_430), .B(n_471), .C(n_499), .Y(n_429) );
NAND3xp33_ASAP7_75t_SL g430 ( .A(n_431), .B(n_444), .C(n_460), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_439), .B2(n_443), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_438), .A2(n_506), .B1(n_508), .B2(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_448), .B2(n_451), .C(n_454), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g462 ( .A(n_448), .Y(n_462) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g492 ( .A(n_450), .Y(n_492) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp33_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B1(n_465), .B2(n_468), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI211xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_474), .B(n_476), .C(n_487), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_475), .A2(n_477), .B1(n_481), .B2(n_484), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g503 ( .A(n_479), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_490), .Y(n_496) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .C(n_510), .D(n_517), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx12f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g539 ( .A(n_528), .Y(n_539) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_528), .Y(n_544) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g551 ( .A(n_530), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
BUFx2_ASAP7_75t_L g560 ( .A(n_532), .Y(n_560) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_533), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_540), .B(n_541), .Y(n_534) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_L g934 ( .A(n_541), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_934), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_553), .B(n_927), .Y(n_546) );
CKINVDCx6p67_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_551), .B(n_941), .Y(n_940) );
OAI22xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_917), .B2(n_918), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx8_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
CKINVDCx10_ASAP7_75t_R g916 ( .A(n_558), .Y(n_916) );
BUFx6f_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g941 ( .A(n_560), .B(n_942), .Y(n_941) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_841), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_776), .C(n_802), .Y(n_562) );
NAND4xp25_ASAP7_75t_SL g563 ( .A(n_564), .B(n_645), .C(n_732), .D(n_756), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_582), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g904 ( .A(n_566), .Y(n_904) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_567), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g647 ( .A(n_568), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g809 ( .A(n_568), .B(n_718), .Y(n_809) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g715 ( .A(n_569), .B(n_716), .Y(n_715) );
INVx3_ASAP7_75t_L g724 ( .A(n_569), .Y(n_724) );
AND2x2_ASAP7_75t_L g833 ( .A(n_569), .B(n_722), .Y(n_833) );
INVx2_ASAP7_75t_L g880 ( .A(n_569), .Y(n_880) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .B(n_580), .Y(n_571) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI21x1_ASAP7_75t_L g694 ( .A1(n_580), .A2(n_695), .B(n_698), .Y(n_694) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_595), .Y(n_582) );
OR2x2_ASAP7_75t_L g849 ( .A(n_583), .B(n_674), .Y(n_849) );
AND2x2_ASAP7_75t_L g861 ( .A(n_583), .B(n_862), .Y(n_861) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g746 ( .A(n_584), .Y(n_746) );
AND2x2_ASAP7_75t_L g800 ( .A(n_584), .B(n_729), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_584), .B(n_818), .Y(n_817) );
AND2x4_ASAP7_75t_L g903 ( .A(n_584), .B(n_785), .Y(n_903) );
AND2x2_ASAP7_75t_L g910 ( .A(n_584), .B(n_597), .Y(n_910) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_585), .Y(n_897) );
INVxp67_ASAP7_75t_L g701 ( .A(n_593), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g843 ( .A1(n_595), .A2(n_789), .B(n_844), .C(n_845), .Y(n_843) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_612), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_596), .B(n_814), .Y(n_825) );
OR2x2_ASAP7_75t_L g840 ( .A(n_596), .B(n_817), .Y(n_840) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_596), .Y(n_852) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g788 ( .A(n_597), .Y(n_788) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g673 ( .A(n_598), .Y(n_673) );
BUFx2_ASAP7_75t_L g706 ( .A(n_598), .Y(n_706) );
OR2x2_ASAP7_75t_L g730 ( .A(n_598), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g735 ( .A(n_598), .B(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g835 ( .A(n_598), .B(n_755), .Y(n_835) );
INVx1_ASAP7_75t_L g892 ( .A(n_598), .Y(n_892) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI21x1_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_606), .B(n_610), .Y(n_601) );
AND2x2_ASAP7_75t_L g707 ( .A(n_612), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g801 ( .A(n_612), .B(n_794), .Y(n_801) );
AND2x2_ASAP7_75t_L g832 ( .A(n_612), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g866 ( .A(n_612), .Y(n_866) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_631), .Y(n_612) );
INVx1_ASAP7_75t_L g716 ( .A(n_613), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_613), .B(n_878), .Y(n_877) );
AO21x1_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_629), .Y(n_613) );
AO21x2_ASAP7_75t_L g720 ( .A1(n_614), .A2(n_615), .B(n_629), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_624), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_621), .B2(n_623), .Y(n_616) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g670 ( .A(n_632), .Y(n_670) );
AND2x2_ASAP7_75t_L g743 ( .A(n_632), .B(n_720), .Y(n_743) );
INVx1_ASAP7_75t_L g752 ( .A(n_632), .Y(n_752) );
INVx1_ASAP7_75t_L g758 ( .A(n_632), .Y(n_758) );
AND2x2_ASAP7_75t_L g770 ( .A(n_632), .B(n_719), .Y(n_770) );
AND2x2_ASAP7_75t_L g805 ( .A(n_632), .B(n_722), .Y(n_805) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_632), .Y(n_824) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_638), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_671), .B1(n_704), .B2(n_707), .C(n_711), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_668), .Y(n_646) );
AND2x2_ASAP7_75t_L g757 ( .A(n_647), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g774 ( .A(n_649), .B(n_724), .Y(n_774) );
OR2x2_ASAP7_75t_L g791 ( .A(n_649), .B(n_670), .Y(n_791) );
AO31x2_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_665), .A3(n_666), .B(n_667), .Y(n_649) );
AO31x2_ASAP7_75t_L g710 ( .A1(n_650), .A2(n_665), .A3(n_666), .B(n_667), .Y(n_710) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22x1_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_658), .B1(n_659), .B2(n_664), .Y(n_651) );
OAI22x1_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g688 ( .A(n_658), .Y(n_688) );
AOI21x1_ASAP7_75t_L g695 ( .A1(n_658), .A2(n_696), .B(n_697), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_659) );
AOI21x1_ASAP7_75t_SL g677 ( .A1(n_664), .A2(n_678), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g723 ( .A(n_667), .Y(n_723) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g839 ( .A(n_669), .B(n_821), .Y(n_839) );
NOR2xp67_ASAP7_75t_L g879 ( .A(n_669), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g768 ( .A1(n_672), .A2(n_769), .B1(n_771), .B2(n_775), .Y(n_768) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_673), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g760 ( .A(n_673), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_673), .B(n_764), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_673), .B(n_797), .Y(n_796) );
NOR2xp67_ASAP7_75t_R g863 ( .A(n_673), .B(n_864), .Y(n_863) );
OR2x2_ASAP7_75t_L g705 ( .A(n_674), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g745 ( .A(n_674), .B(n_746), .Y(n_745) );
OR2x6_ASAP7_75t_L g674 ( .A(n_675), .B(n_690), .Y(n_674) );
INVx2_ASAP7_75t_L g785 ( .A(n_675), .Y(n_785) );
OR2x2_ASAP7_75t_SL g815 ( .A(n_675), .B(n_736), .Y(n_815) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g729 ( .A(n_676), .Y(n_729) );
OAI21x1_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_683), .B(n_689), .Y(n_676) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AND2x2_ASAP7_75t_L g763 ( .A(n_690), .B(n_728), .Y(n_763) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_691), .Y(n_731) );
INVx2_ASAP7_75t_L g755 ( .A(n_691), .Y(n_755) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI21x1_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_703), .Y(n_692) );
OA21x2_ASAP7_75t_L g736 ( .A1(n_694), .A2(n_703), .B(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_702), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g893 ( .A1(n_704), .A2(n_894), .B(n_898), .Y(n_893) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g838 ( .A(n_706), .B(n_800), .Y(n_838) );
OR2x2_ASAP7_75t_L g868 ( .A(n_706), .B(n_754), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_706), .B(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g740 ( .A(n_709), .B(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g750 ( .A(n_709), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g844 ( .A(n_709), .Y(n_844) );
BUFx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g714 ( .A(n_710), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_717), .B(n_725), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_712), .A2(n_748), .B1(n_750), .B2(n_753), .Y(n_747) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g742 ( .A(n_714), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_714), .B(n_770), .Y(n_769) );
OR2x6_ASAP7_75t_L g779 ( .A(n_714), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g794 ( .A(n_714), .Y(n_794) );
INVx1_ASAP7_75t_L g780 ( .A(n_715), .Y(n_780) );
INVx1_ASAP7_75t_L g821 ( .A(n_715), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g855 ( .A(n_718), .Y(n_855) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_719), .B(n_724), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_719), .B(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g830 ( .A(n_719), .Y(n_830) );
INVx3_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_721), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g829 ( .A(n_721), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g867 ( .A(n_721), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_721), .B(n_743), .Y(n_869) );
AND2x2_ASAP7_75t_L g906 ( .A(n_721), .B(n_907), .Y(n_906) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g878 ( .A(n_722), .Y(n_878) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_730), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_727), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g857 ( .A(n_727), .B(n_788), .Y(n_857) );
INVx1_ASAP7_75t_L g873 ( .A(n_727), .Y(n_873) );
AOI322xp5_ASAP7_75t_L g905 ( .A1(n_727), .A2(n_906), .A3(n_908), .B1(n_910), .B2(n_911), .C1(n_913), .C2(n_914), .Y(n_905) );
AND2x4_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AND2x4_ASAP7_75t_L g784 ( .A(n_728), .B(n_785), .Y(n_784) );
AND2x4_ASAP7_75t_L g834 ( .A(n_728), .B(n_835), .Y(n_834) );
OR2x2_ASAP7_75t_L g846 ( .A(n_728), .B(n_815), .Y(n_846) );
AND2x2_ASAP7_75t_L g749 ( .A(n_729), .B(n_736), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_729), .B(n_755), .Y(n_754) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_729), .Y(n_764) );
INVx1_ASAP7_75t_L g798 ( .A(n_729), .Y(n_798) );
INVx2_ASAP7_75t_L g909 ( .A(n_730), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_739), .B1(n_742), .B2(n_744), .C(n_747), .Y(n_732) );
OR2x2_ASAP7_75t_L g895 ( .A(n_734), .B(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g799 ( .A(n_735), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g902 ( .A(n_735), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g790 ( .A(n_741), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g806 ( .A(n_741), .Y(n_806) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_743), .Y(n_767) );
AND2x2_ASAP7_75t_L g898 ( .A(n_743), .B(n_833), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_744), .A2(n_781), .B1(n_901), .B2(n_902), .Y(n_900) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g753 ( .A(n_746), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g811 ( .A(n_748), .Y(n_811) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_751), .Y(n_907) );
INVx2_ASAP7_75t_L g761 ( .A(n_754), .Y(n_761) );
INVx1_ASAP7_75t_L g818 ( .A(n_755), .Y(n_818) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_755), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B1(n_762), .B2(n_765), .C(n_768), .Y(n_756) );
INVx2_ASAP7_75t_L g773 ( .A(n_758), .Y(n_773) );
AND2x4_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_760), .B(n_784), .Y(n_783) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_761), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_762), .B(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
AND2x2_ASAP7_75t_L g797 ( .A(n_763), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g871 ( .A(n_767), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_770), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_770), .B(n_794), .Y(n_912) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_772), .B(n_855), .Y(n_854) );
NOR2x1p5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g781 ( .A(n_773), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_777), .B(n_792), .Y(n_776) );
AOI32xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_781), .A3(n_782), .B1(n_786), .B2(n_789), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g913 ( .A(n_779), .Y(n_913) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g888 ( .A(n_785), .Y(n_888) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_SL g810 ( .A(n_791), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B1(n_799), .B2(n_801), .Y(n_792) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g864 ( .A(n_798), .Y(n_864) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_800), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_800), .B(n_835), .Y(n_872) );
INVx1_ASAP7_75t_L g889 ( .A(n_801), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_826), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_808), .B2(n_811), .C(n_812), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g820 ( .A(n_805), .Y(n_820) );
AND2x4_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_819), .B1(n_822), .B2(n_825), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
AND2x2_ASAP7_75t_L g914 ( .A(n_814), .B(n_910), .Y(n_914) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OR2x2_ASAP7_75t_L g890 ( .A(n_815), .B(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
OR2x2_ASAP7_75t_L g882 ( .A(n_823), .B(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_834), .B(n_836), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_831), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_828), .A2(n_837), .B1(n_839), .B2(n_840), .Y(n_836) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_SL g858 ( .A(n_839), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_881), .C(n_899), .Y(n_841) );
NAND3xp33_ASAP7_75t_SL g842 ( .A(n_843), .B(n_847), .C(n_856), .Y(n_842) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OAI31xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_850), .A3(n_851), .B(n_853), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g901 ( .A(n_855), .Y(n_901) );
AOI211xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B(n_859), .C(n_870), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_865), .B1(n_868), .B2(n_869), .Y(n_859) );
NOR2xp33_ASAP7_75t_SL g860 ( .A(n_861), .B(n_863), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_861), .B(n_886), .Y(n_885) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_876), .B(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g884 ( .A(n_880), .Y(n_884) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_885), .B1(n_889), .B2(n_890), .C(n_893), .Y(n_881) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_904), .B(n_905), .Y(n_899) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_SL g915 ( .A(n_916), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g926 ( .A(n_919), .Y(n_926) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
BUFx3_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx3_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx3_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
CKINVDCx6p67_ASAP7_75t_R g947 ( .A(n_936), .Y(n_947) );
OR2x6_ASAP7_75t_L g936 ( .A(n_937), .B(n_940), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_947), .Y(n_946) );
endmodule