module real_jpeg_1625_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_60),
.B1(n_64),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_79),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_60),
.B1(n_64),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_3),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_4),
.A2(n_35),
.B(n_49),
.C(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_4),
.B(n_35),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_50)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_4),
.A2(n_9),
.B(n_35),
.C(n_136),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_47),
.B1(n_60),
.B2(n_64),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_9),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_50),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_37),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_60),
.C(n_63),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_82),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_9),
.B(n_117),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_60),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_11),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_60),
.B1(n_64),
.B2(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_14),
.A2(n_27),
.B1(n_51),
.B2(n_52),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_35),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_27),
.B1(n_60),
.B2(n_64),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_123),
.B1(n_200),
.B2(n_201),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_18),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_97),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_86),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_21),
.B(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_45),
.C(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_36)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_32),
.A3(n_35),
.B1(n_39),
.B2(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_28),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_28)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_29),
.B(n_33),
.Y(n_75)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_37),
.A2(n_51),
.B(n_54),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_37),
.A2(n_119),
.B(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_41),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_50),
.B2(n_55),
.Y(n_45)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_91),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_52),
.B(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_65),
.B(n_68),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_59),
.A2(n_68),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_59),
.A2(n_131),
.B1(n_149),
.B2(n_161),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_60),
.B(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_69),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_117),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_86),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_80),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_80),
.A2(n_81),
.B1(n_153),
.B2(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_96),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_81),
.B(n_140),
.Y(n_155)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_84),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_82),
.A2(n_139),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_95),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_102),
.A2(n_104),
.B(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_143),
.B(n_199),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_141),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_141),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_134),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_126),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_129),
.B(n_134),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_161),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_137),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_194),
.B(n_198),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_163),
.B(n_193),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_156),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_152),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_175),
.B(n_192),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_186),
.B(n_191),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_185),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_184),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_197),
.Y(n_198)
);


endmodule