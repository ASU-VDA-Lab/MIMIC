module fake_jpeg_31752_n_71 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_37),
.B(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_11),
.B1(n_23),
.B2(n_21),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_28),
.B1(n_2),
.B2(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_26),
.B1(n_32),
.B2(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_26),
.B1(n_25),
.B2(n_38),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_32),
.B(n_14),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_48),
.B(n_33),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_8),
.B(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_51),
.B1(n_57),
.B2(n_5),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_44),
.B1(n_42),
.B2(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_54),
.B1(n_57),
.B2(n_52),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_30),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

OAI22x1_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_15),
.B1(n_16),
.B2(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_5),
.C(n_6),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_58),
.C(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_64),
.B1(n_58),
.B2(n_59),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_65),
.Y(n_71)
);


endmodule