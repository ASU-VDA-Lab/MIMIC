module fake_jpeg_6179_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_20),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_1),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_2),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_36),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_39),
.CON(n_45),
.SN(n_45)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_19),
.B1(n_18),
.B2(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_19),
.B1(n_18),
.B2(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_21),
.B(n_25),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_26),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_26),
.B(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_50),
.B1(n_56),
.B2(n_45),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_45),
.B(n_44),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_42),
.B(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_32),
.B1(n_33),
.B2(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_10),
.B1(n_16),
.B2(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_64),
.A3(n_60),
.B1(n_63),
.B2(n_57),
.C1(n_65),
.C2(n_16),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_57),
.B(n_10),
.C(n_4),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_70),
.Y(n_72)
);


endmodule