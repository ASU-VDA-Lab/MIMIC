module real_aes_18125_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_559;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_0), .A2(n_76), .B1(n_1077), .B2(n_1082), .Y(n_1081) );
INVxp33_ASAP7_75t_SL g1113 ( .A(n_0), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_1), .A2(n_82), .B1(n_514), .B2(n_555), .Y(n_980) );
OAI22xp33_ASAP7_75t_SL g999 ( .A1(n_1), .A2(n_240), .B1(n_483), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g628 ( .A(n_2), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_3), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_4), .A2(n_197), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g752 ( .A(n_4), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_5), .A2(n_119), .B1(n_569), .B2(n_1375), .Y(n_1374) );
AOI22xp33_ASAP7_75t_SL g1395 ( .A1(n_5), .A2(n_123), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx1_ASAP7_75t_L g1015 ( .A(n_6), .Y(n_1015) );
OAI221xp5_ASAP7_75t_SL g1046 ( .A1(n_6), .A2(n_91), .B1(n_336), .B2(n_542), .C(n_549), .Y(n_1046) );
INVx1_ASAP7_75t_L g687 ( .A(n_7), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_7), .A2(n_136), .B1(n_750), .B2(n_755), .C(n_756), .Y(n_754) );
AOI22xp5_ASAP7_75t_SL g1190 ( .A1(n_8), .A2(n_233), .B1(n_1183), .B2(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g972 ( .A(n_9), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_10), .A2(n_18), .B1(n_399), .B2(n_403), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_10), .A2(n_18), .B1(n_438), .B2(n_441), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_11), .A2(n_185), .B1(n_685), .B2(n_1444), .C(n_1445), .Y(n_1443) );
INVx1_ASAP7_75t_L g1472 ( .A(n_11), .Y(n_1472) );
INVx1_ASAP7_75t_L g262 ( .A(n_12), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_12), .B(n_272), .Y(n_343) );
AND2x2_ASAP7_75t_L g458 ( .A(n_12), .B(n_402), .Y(n_458) );
AND2x2_ASAP7_75t_L g481 ( .A(n_12), .B(n_211), .Y(n_481) );
INVx1_ASAP7_75t_L g334 ( .A(n_13), .Y(n_334) );
INVx1_ASAP7_75t_L g852 ( .A(n_14), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_14), .A2(n_33), .B1(n_873), .B2(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g909 ( .A(n_15), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_15), .A2(n_230), .B1(n_708), .B2(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_SL g1373 ( .A1(n_16), .A2(n_147), .B1(n_522), .B2(n_563), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_16), .A2(n_19), .B1(n_987), .B2(n_1389), .C(n_1391), .Y(n_1388) );
INVx2_ASAP7_75t_L g1178 ( .A(n_17), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_17), .B(n_1179), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_17), .B(n_107), .Y(n_1186) );
AOI22xp33_ASAP7_75t_SL g1378 ( .A1(n_19), .A2(n_30), .B1(n_575), .B2(n_1076), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_20), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_20), .A2(n_161), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g1371 ( .A(n_21), .Y(n_1371) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_22), .A2(n_204), .B1(n_953), .B2(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1402 ( .A(n_22), .Y(n_1402) );
AOI22xp5_ASAP7_75t_SL g1205 ( .A1(n_23), .A2(n_127), .B1(n_1183), .B2(n_1191), .Y(n_1205) );
XNOR2x2_ASAP7_75t_L g673 ( .A(n_24), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_SL g1195 ( .A1(n_25), .A2(n_224), .B1(n_1180), .B2(n_1185), .Y(n_1195) );
INVx1_ASAP7_75t_L g802 ( .A(n_26), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_27), .A2(n_81), .B1(n_786), .B2(n_931), .C(n_1085), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_27), .A2(n_28), .B1(n_876), .B2(n_907), .Y(n_1120) );
AOI22xp33_ASAP7_75t_SL g1073 ( .A1(n_28), .A2(n_126), .B1(n_1074), .B2(n_1077), .Y(n_1073) );
XOR2x2_ASAP7_75t_L g450 ( .A(n_29), .B(n_451), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g1405 ( .A1(n_30), .A2(n_614), .B(n_1406), .C(n_1413), .Y(n_1405) );
INVx1_ASAP7_75t_L g894 ( .A(n_31), .Y(n_894) );
INVx1_ASAP7_75t_L g1088 ( .A(n_32), .Y(n_1088) );
OA222x2_ASAP7_75t_L g1102 ( .A1(n_32), .A2(n_153), .B1(n_245), .B2(n_897), .C1(n_1103), .C2(n_1104), .Y(n_1102) );
INVx1_ASAP7_75t_L g862 ( .A(n_33), .Y(n_862) );
OAI22xp5_ASAP7_75t_SL g947 ( .A1(n_34), .A2(n_948), .B1(n_949), .B2(n_1002), .Y(n_947) );
INVx1_ASAP7_75t_L g1002 ( .A(n_34), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_34), .A2(n_948), .B1(n_949), .B2(n_1002), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_34), .A2(n_164), .B1(n_1175), .B2(n_1180), .Y(n_1174) );
INVx1_ASAP7_75t_L g688 ( .A(n_35), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_35), .A2(n_79), .B1(n_746), .B2(n_748), .C(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g859 ( .A(n_36), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_36), .A2(n_165), .B1(n_755), .B2(n_873), .Y(n_879) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_37), .A2(n_237), .B1(n_599), .B2(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_37), .A2(n_237), .B1(n_664), .B2(n_666), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g1078 ( .A1(n_38), .A2(n_196), .B1(n_796), .B2(n_1079), .C(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g1117 ( .A(n_38), .Y(n_1117) );
AOI211xp5_ASAP7_75t_L g1434 ( .A1(n_39), .A2(n_931), .B(n_1435), .C(n_1437), .Y(n_1434) );
INVx1_ASAP7_75t_L g1467 ( .A(n_39), .Y(n_1467) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_40), .A2(n_68), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_707) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_40), .Y(n_737) );
INVx1_ASAP7_75t_L g883 ( .A(n_41), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_42), .A2(n_102), .B1(n_1183), .B2(n_1201), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_43), .A2(n_65), .B1(n_514), .B2(n_555), .Y(n_1384) );
OAI211xp5_ASAP7_75t_L g1386 ( .A1(n_43), .A2(n_483), .B(n_1387), .C(n_1398), .Y(n_1386) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_44), .A2(n_897), .B(n_899), .Y(n_896) );
OAI221xp5_ASAP7_75t_L g938 ( .A1(n_44), .A2(n_55), .B1(n_939), .B2(n_940), .C(n_941), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_45), .A2(n_156), .B1(n_708), .B2(n_710), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_45), .A2(n_84), .B1(n_830), .B2(n_832), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_46), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_46), .A2(n_51), .B1(n_562), .B2(n_563), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_47), .A2(n_167), .B1(n_1183), .B2(n_1185), .Y(n_1182) );
INVx1_ASAP7_75t_L g631 ( .A(n_48), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g1213 ( .A1(n_49), .A2(n_89), .B1(n_1175), .B2(n_1183), .Y(n_1213) );
XNOR2x2_ASAP7_75t_L g1365 ( .A(n_49), .B(n_1366), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_49), .A2(n_1423), .B1(n_1474), .B2(n_1476), .Y(n_1422) );
INVx1_ASAP7_75t_L g298 ( .A(n_50), .Y(n_298) );
INVx1_ASAP7_75t_L g304 ( .A(n_50), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_51), .A2(n_161), .B1(n_489), .B2(n_490), .C(n_494), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_52), .A2(n_144), .B1(n_729), .B2(n_876), .Y(n_1032) );
INVx1_ASAP7_75t_L g1049 ( .A(n_52), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1431 ( .A1(n_53), .A2(n_222), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_53), .A2(n_120), .B1(n_515), .B2(n_732), .Y(n_1456) );
INVx1_ASAP7_75t_L g910 ( .A(n_54), .Y(n_910) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_55), .Y(n_944) );
INVx1_ASAP7_75t_L g791 ( .A(n_56), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_57), .A2(n_158), .B1(n_576), .B2(n_955), .C(n_957), .Y(n_954) );
OAI211xp5_ASAP7_75t_L g982 ( .A1(n_57), .A2(n_983), .B(n_984), .C(n_988), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_58), .A2(n_109), .B1(n_702), .B2(n_705), .C(n_841), .Y(n_840) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_58), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g1217 ( .A1(n_59), .A2(n_242), .B1(n_1175), .B2(n_1180), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_60), .A2(n_123), .B1(n_566), .B2(n_569), .Y(n_1376) );
AOI221xp5_ASAP7_75t_L g1407 ( .A1(n_60), .A2(n_119), .B1(n_1408), .B2(n_1409), .C(n_1410), .Y(n_1407) );
INVx1_ASAP7_75t_L g388 ( .A(n_61), .Y(n_388) );
INVx1_ASAP7_75t_L g255 ( .A(n_62), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_63), .A2(n_203), .B1(n_702), .B2(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g744 ( .A(n_63), .Y(n_744) );
INVx2_ASAP7_75t_L g289 ( .A(n_64), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_66), .A2(n_178), .B1(n_678), .B2(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g739 ( .A(n_66), .Y(n_739) );
INVx1_ASAP7_75t_L g622 ( .A(n_67), .Y(n_622) );
INVx1_ASAP7_75t_L g767 ( .A(n_68), .Y(n_767) );
INVx1_ASAP7_75t_L g1138 ( .A(n_69), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_69), .A2(n_210), .B1(n_729), .B2(n_876), .Y(n_1160) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_70), .A2(n_77), .B1(n_1175), .B2(n_1183), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1148 ( .A(n_71), .Y(n_1148) );
INVx1_ASAP7_75t_L g299 ( .A(n_72), .Y(n_299) );
INVx1_ASAP7_75t_L g321 ( .A(n_73), .Y(n_321) );
INVx1_ASAP7_75t_L g291 ( .A(n_74), .Y(n_291) );
AOI21xp33_ASAP7_75t_L g795 ( .A1(n_75), .A2(n_568), .B(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g820 ( .A(n_75), .Y(n_820) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_76), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_78), .A2(n_381), .B(n_382), .C(n_387), .Y(n_380) );
INVx1_ASAP7_75t_L g436 ( .A(n_78), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_79), .A2(n_198), .B1(n_685), .B2(n_691), .C(n_693), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_80), .A2(n_169), .B1(n_490), .B2(n_494), .C(n_1031), .Y(n_1033) );
INVx1_ASAP7_75t_L g1050 ( .A(n_80), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_81), .A2(n_196), .B1(n_1031), .B2(n_1110), .C(n_1111), .Y(n_1109) );
INVx1_ASAP7_75t_L g623 ( .A(n_83), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_84), .A2(n_155), .B1(n_1145), .B2(n_1146), .C(n_1147), .Y(n_1144) );
INVx1_ASAP7_75t_L g1096 ( .A(n_85), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1100 ( .A(n_85), .B(n_809), .Y(n_1100) );
INVx1_ASAP7_75t_L g307 ( .A(n_86), .Y(n_307) );
INVx1_ASAP7_75t_L g860 ( .A(n_87), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_87), .A2(n_212), .B1(n_729), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g1212 ( .A1(n_88), .A2(n_177), .B1(n_1180), .B2(n_1191), .Y(n_1212) );
INVx1_ASAP7_75t_L g612 ( .A(n_90), .Y(n_612) );
INVx1_ASAP7_75t_L g1026 ( .A(n_91), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_92), .Y(n_847) );
INVx1_ASAP7_75t_L g510 ( .A(n_93), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_94), .A2(n_170), .B1(n_678), .B2(n_681), .Y(n_803) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_94), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1442 ( .A1(n_95), .A2(n_120), .B1(n_678), .B2(n_681), .Y(n_1442) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_95), .A2(n_809), .B(n_1450), .C(n_1453), .Y(n_1449) );
INVx1_ASAP7_75t_L g1097 ( .A(n_96), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_96), .A2(n_174), .B1(n_515), .B2(n_732), .Y(n_1121) );
OAI221xp5_ASAP7_75t_L g1011 ( .A1(n_97), .A2(n_247), .B1(n_995), .B2(n_1012), .C(n_1013), .Y(n_1011) );
INVx1_ASAP7_75t_L g1038 ( .A(n_97), .Y(n_1038) );
INVx1_ASAP7_75t_L g1441 ( .A(n_98), .Y(n_1441) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_99), .Y(n_257) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_99), .B(n_255), .Y(n_1176) );
INVx1_ASAP7_75t_L g324 ( .A(n_100), .Y(n_324) );
OA22x2_ASAP7_75t_L g581 ( .A1(n_101), .A2(n_582), .B1(n_670), .B2(n_671), .Y(n_581) );
INVxp67_ASAP7_75t_L g671 ( .A(n_101), .Y(n_671) );
INVx1_ASAP7_75t_L g1447 ( .A(n_103), .Y(n_1447) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_104), .A2(n_148), .B1(n_1175), .B2(n_1180), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1424 ( .A1(n_105), .A2(n_1425), .B1(n_1426), .B2(n_1473), .Y(n_1424) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_105), .Y(n_1425) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_106), .A2(n_173), .B1(n_492), .B2(n_755), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_106), .A2(n_159), .B1(n_566), .B2(n_796), .C(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g1179 ( .A(n_107), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_107), .B(n_1178), .Y(n_1184) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_108), .A2(n_175), .B1(n_1175), .B2(n_1180), .Y(n_1192) );
INVx1_ASAP7_75t_L g882 ( .A(n_109), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_110), .Y(n_536) );
INVx1_ASAP7_75t_L g1446 ( .A(n_111), .Y(n_1446) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_112), .A2(n_238), .B1(n_496), .B2(n_500), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_112), .A2(n_145), .B1(n_566), .B2(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g607 ( .A(n_113), .Y(n_607) );
INVx1_ASAP7_75t_L g1021 ( .A(n_114), .Y(n_1021) );
OAI21xp33_ASAP7_75t_L g1044 ( .A1(n_114), .A2(n_532), .B(n_1045), .Y(n_1044) );
INVx2_ASAP7_75t_L g288 ( .A(n_115), .Y(n_288) );
INVx1_ASAP7_75t_L g332 ( .A(n_115), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_115), .B(n_289), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_116), .A2(n_248), .B1(n_587), .B2(n_589), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_116), .A2(n_248), .B1(n_264), .B2(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g793 ( .A(n_117), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g1133 ( .A(n_118), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_121), .A2(n_232), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_121), .A2(n_202), .B1(n_562), .B2(n_786), .C(n_931), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_122), .A2(n_1006), .B1(n_1007), .B2(n_1008), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_122), .Y(n_1006) );
INVx1_ASAP7_75t_L g863 ( .A(n_124), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_124), .A2(n_179), .B1(n_501), .B2(n_881), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_125), .A2(n_168), .B1(n_407), .B2(n_408), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_125), .A2(n_168), .B1(n_418), .B2(n_419), .Y(n_417) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_126), .Y(n_1112) );
INVx1_ASAP7_75t_L g699 ( .A(n_128), .Y(n_699) );
INVx1_ASAP7_75t_L g313 ( .A(n_129), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_130), .A2(n_181), .B1(n_906), .B2(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1058 ( .A(n_130), .Y(n_1058) );
INVx1_ASAP7_75t_L g620 ( .A(n_131), .Y(n_620) );
INVx1_ASAP7_75t_L g1271 ( .A(n_132), .Y(n_1271) );
XOR2x2_ASAP7_75t_L g774 ( .A(n_133), .B(n_775), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_134), .A2(n_705), .B1(n_1136), .B2(n_1139), .Y(n_1135) );
INVx1_ASAP7_75t_L g1154 ( .A(n_134), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1432 ( .A1(n_135), .A2(n_139), .B1(n_702), .B2(n_705), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1454 ( .A(n_135), .Y(n_1454) );
INVx1_ASAP7_75t_L g694 ( .A(n_136), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_137), .A2(n_201), .B1(n_906), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_137), .A2(n_232), .B1(n_562), .B2(n_929), .Y(n_928) );
AOI221xp5_ASAP7_75t_SL g1030 ( .A1(n_138), .A2(n_160), .B1(n_490), .B2(n_998), .C(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1052 ( .A(n_138), .Y(n_1052) );
INVxp67_ASAP7_75t_SL g1451 ( .A(n_139), .Y(n_1451) );
INVx1_ASAP7_75t_L g463 ( .A(n_140), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_140), .A2(n_238), .B1(n_569), .B2(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_141), .A2(n_172), .B1(n_1183), .B2(n_1201), .Y(n_1200) );
BUFx3_ASAP7_75t_L g296 ( .A(n_142), .Y(n_296) );
INVx1_ASAP7_75t_L g965 ( .A(n_143), .Y(n_965) );
INVx1_ASAP7_75t_L g1060 ( .A(n_144), .Y(n_1060) );
INVx1_ASAP7_75t_L g465 ( .A(n_145), .Y(n_465) );
INVx1_ASAP7_75t_L g778 ( .A(n_146), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_147), .B(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1436 ( .A(n_149), .Y(n_1436) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_150), .A2(n_205), .B1(n_1183), .B2(n_1191), .Y(n_1218) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_151), .Y(n_269) );
INVx1_ASAP7_75t_L g900 ( .A(n_152), .Y(n_900) );
INVx1_ASAP7_75t_L g1099 ( .A(n_153), .Y(n_1099) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_154), .A2(n_514), .B(n_520), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g1152 ( .A1(n_155), .A2(n_720), .B(n_1153), .C(n_1156), .Y(n_1152) );
INVx1_ASAP7_75t_L g1155 ( .A(n_156), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g1132 ( .A(n_157), .Y(n_1132) );
OAI221xp5_ASAP7_75t_SL g989 ( .A1(n_158), .A2(n_190), .B1(n_477), .B2(n_990), .C(n_992), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_159), .A2(n_202), .B1(n_916), .B2(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g1057 ( .A(n_160), .Y(n_1057) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_162), .A2(n_562), .B(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_162), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_163), .Y(n_1028) );
INVx1_ASAP7_75t_L g850 ( .A(n_165), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_166), .A2(n_225), .B1(n_684), .B2(n_974), .Y(n_973) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_166), .Y(n_996) );
INVx1_ASAP7_75t_L g1061 ( .A(n_169), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_170), .A2(n_199), .B1(n_769), .B2(n_830), .C(n_832), .Y(n_829) );
INVx1_ASAP7_75t_L g1141 ( .A(n_171), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_171), .A2(n_183), .B1(n_485), .B2(n_876), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_173), .A2(n_201), .B1(n_929), .B2(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g1087 ( .A(n_174), .Y(n_1087) );
OAI211xp5_ASAP7_75t_SL g590 ( .A1(n_176), .A2(n_423), .B(n_591), .C(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g660 ( .A(n_176), .Y(n_660) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_178), .Y(n_762) );
INVx1_ASAP7_75t_L g856 ( .A(n_179), .Y(n_856) );
INVx1_ASAP7_75t_L g596 ( .A(n_180), .Y(n_596) );
INVx1_ASAP7_75t_L g1055 ( .A(n_181), .Y(n_1055) );
INVx1_ASAP7_75t_L g801 ( .A(n_182), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_183), .A2(n_210), .B1(n_798), .B2(n_929), .C(n_1131), .Y(n_1130) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_184), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_184), .A2(n_216), .B1(n_750), .B2(n_986), .C(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1460 ( .A(n_185), .Y(n_1460) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_186), .Y(n_268) );
OAI222xp33_ASAP7_75t_L g453 ( .A1(n_187), .A2(n_236), .B1(n_454), .B2(n_459), .C1(n_469), .C2(n_477), .Y(n_453) );
INVx1_ASAP7_75t_L g539 ( .A(n_187), .Y(n_539) );
INVx1_ASAP7_75t_L g788 ( .A(n_188), .Y(n_788) );
INVx1_ASAP7_75t_L g843 ( .A(n_189), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_189), .A2(n_191), .B1(n_515), .B2(n_732), .Y(n_870) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_190), .Y(n_951) );
INVx1_ASAP7_75t_L g846 ( .A(n_191), .Y(n_846) );
INVx1_ASAP7_75t_L g1439 ( .A(n_192), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g1137 ( .A(n_193), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_194), .Y(n_1383) );
INVx1_ASAP7_75t_L g597 ( .A(n_195), .Y(n_597) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_195), .A2(n_382), .B(n_656), .C(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g757 ( .A(n_197), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_198), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g779 ( .A1(n_199), .A2(n_214), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_779) );
INVx1_ASAP7_75t_L g506 ( .A(n_200), .Y(n_506) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_203), .Y(n_718) );
INVx1_ASAP7_75t_L g1399 ( .A(n_204), .Y(n_1399) );
INVx1_ASAP7_75t_L g1370 ( .A(n_206), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_207), .A2(n_556), .B(n_712), .C(n_845), .Y(n_844) );
INVxp33_ASAP7_75t_SL g869 ( .A(n_207), .Y(n_869) );
INVx1_ASAP7_75t_L g1430 ( .A(n_208), .Y(n_1430) );
INVx1_ASAP7_75t_L g966 ( .A(n_209), .Y(n_966) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_209), .A2(n_225), .B1(n_873), .B2(n_986), .C(n_987), .Y(n_985) );
BUFx3_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
INVx1_ASAP7_75t_L g402 ( .A(n_211), .Y(n_402) );
INVx1_ASAP7_75t_L g854 ( .A(n_212), .Y(n_854) );
INVx1_ASAP7_75t_L g1122 ( .A(n_213), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_214), .Y(n_834) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_215), .A2(n_483), .B(n_487), .C(n_503), .Y(n_482) );
INVx1_ASAP7_75t_L g553 ( .A(n_215), .Y(n_553) );
INVx1_ASAP7_75t_L g968 ( .A(n_216), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_217), .A2(n_245), .B1(n_971), .B2(n_1093), .C(n_1095), .Y(n_1092) );
INVxp67_ASAP7_75t_SL g1106 ( .A(n_217), .Y(n_1106) );
INVx1_ASAP7_75t_L g286 ( .A(n_218), .Y(n_286) );
INVx1_ASAP7_75t_L g331 ( .A(n_218), .Y(n_331) );
INVx2_ASAP7_75t_L g342 ( .A(n_218), .Y(n_342) );
XOR2x2_ASAP7_75t_L g278 ( .A(n_219), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g695 ( .A(n_220), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_221), .A2(n_229), .B1(n_570), .B2(n_798), .Y(n_797) );
INVxp67_ASAP7_75t_SL g826 ( .A(n_221), .Y(n_826) );
INVxp67_ASAP7_75t_SL g1452 ( .A(n_222), .Y(n_1452) );
INVx1_ASAP7_75t_L g1126 ( .A(n_223), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_223), .A2(n_246), .B1(n_1175), .B2(n_1180), .Y(n_1204) );
INVx1_ASAP7_75t_L g979 ( .A(n_226), .Y(n_979) );
INVx1_ASAP7_75t_L g1143 ( .A(n_227), .Y(n_1143) );
INVx1_ASAP7_75t_L g782 ( .A(n_228), .Y(n_782) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_229), .Y(n_815) );
INVx1_ASAP7_75t_L g901 ( .A(n_230), .Y(n_901) );
INVx1_ASAP7_75t_L g1269 ( .A(n_231), .Y(n_1269) );
OAI21xp33_ASAP7_75t_SL g838 ( .A1(n_234), .A2(n_809), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g842 ( .A(n_234), .Y(n_842) );
INVx1_ASAP7_75t_L g337 ( .A(n_235), .Y(n_337) );
INVx1_ASAP7_75t_L g546 ( .A(n_236), .Y(n_546) );
INVx1_ASAP7_75t_L g963 ( .A(n_239), .Y(n_963) );
OAI322xp33_ASAP7_75t_SL g958 ( .A1(n_240), .A2(n_325), .A3(n_633), .B1(n_959), .B2(n_964), .C1(n_967), .C2(n_975), .Y(n_958) );
INVx1_ASAP7_75t_L g392 ( .A(n_241), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_241), .A2(n_335), .B(n_423), .C(n_427), .Y(n_422) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_242), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g1014 ( .A(n_243), .Y(n_1014) );
INVx1_ASAP7_75t_L g616 ( .A(n_244), .Y(n_616) );
INVx1_ASAP7_75t_L g1040 ( .A(n_247), .Y(n_1040) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_273), .B(n_1166), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_258), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1421 ( .A(n_252), .B(n_261), .Y(n_1421) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g1475 ( .A(n_254), .B(n_257), .Y(n_1475) );
INVx1_ASAP7_75t_L g1477 ( .A(n_254), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g1479 ( .A(n_257), .B(n_1477), .Y(n_1479) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g413 ( .A(n_261), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g375 ( .A(n_262), .B(n_272), .Y(n_375) );
AND2x4_ASAP7_75t_L g468 ( .A(n_262), .B(n_271), .Y(n_468) );
INVx1_ASAP7_75t_L g407 ( .A(n_263), .Y(n_407) );
AND2x4_ASAP7_75t_SL g1420 ( .A(n_263), .B(n_1421), .Y(n_1420) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_270), .Y(n_264) );
OR2x6_ASAP7_75t_L g400 ( .A(n_265), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g611 ( .A(n_265), .Y(n_611) );
INVxp67_ASAP7_75t_L g1412 ( .A(n_265), .Y(n_1412) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g348 ( .A(n_266), .Y(n_348) );
BUFx4f_ASAP7_75t_L g627 ( .A(n_266), .Y(n_627) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g354 ( .A(n_268), .Y(n_354) );
INVx2_ASAP7_75t_L g359 ( .A(n_268), .Y(n_359) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_268), .B(n_269), .Y(n_364) );
AND2x2_ASAP7_75t_L g386 ( .A(n_268), .B(n_269), .Y(n_386) );
INVx1_ASAP7_75t_L g397 ( .A(n_268), .Y(n_397) );
AND2x2_ASAP7_75t_L g410 ( .A(n_268), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_269), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g358 ( .A(n_269), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g391 ( .A(n_269), .Y(n_391) );
INVx2_ASAP7_75t_L g411 ( .A(n_269), .Y(n_411) );
AND2x2_ASAP7_75t_L g486 ( .A(n_269), .B(n_354), .Y(n_486) );
INVx1_ASAP7_75t_L g499 ( .A(n_269), .Y(n_499) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g384 ( .A(n_271), .Y(n_384) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g390 ( .A(n_272), .Y(n_390) );
AND2x4_ASAP7_75t_L g395 ( .A(n_272), .B(n_396), .Y(n_395) );
XNOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_885), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_772), .B2(n_884), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AO22x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_578), .B1(n_579), .B2(n_771), .Y(n_276) );
INVx1_ASAP7_75t_L g771 ( .A(n_277), .Y(n_771) );
XNOR2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_450), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_379), .C(n_416), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_338), .Y(n_280) );
OAI33xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_290), .A3(n_306), .B1(n_318), .B2(n_325), .B3(n_333), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx4f_ASAP7_75t_L g634 ( .A(n_283), .Y(n_634) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx1_ASAP7_75t_L g374 ( .A(n_284), .Y(n_374) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_284), .Y(n_449) );
OR2x2_ASAP7_75t_L g518 ( .A(n_284), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g828 ( .A(n_284), .B(n_375), .Y(n_828) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g415 ( .A(n_285), .Y(n_415) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g796 ( .A(n_287), .Y(n_796) );
NAND2xp33_ASAP7_75t_SL g287 ( .A(n_288), .B(n_289), .Y(n_287) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_288), .Y(n_447) );
INVx1_ASAP7_75t_L g545 ( .A(n_288), .Y(n_545) );
AND3x4_ASAP7_75t_L g560 ( .A(n_288), .B(n_431), .C(n_512), .Y(n_560) );
AND2x2_ASAP7_75t_L g689 ( .A(n_288), .B(n_431), .Y(n_689) );
INVx3_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
BUFx3_ASAP7_75t_L g431 ( .A(n_289), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B1(n_299), .B2(n_300), .Y(n_290) );
OAI22xp5_ASAP7_75t_SL g344 ( .A1(n_291), .A2(n_334), .B1(n_345), .B2(n_349), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_292), .A2(n_334), .B1(n_335), .B2(n_337), .Y(n_333) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_294), .A2(n_336), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_294), .A2(n_300), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_294), .A2(n_336), .B1(n_1060), .B2(n_1061), .Y(n_1059) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_294), .A2(n_593), .B1(n_696), .B2(n_1137), .C(n_1138), .Y(n_1136) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x4_ASAP7_75t_L g418 ( .A(n_295), .B(n_329), .Y(n_418) );
OR2x4_ASAP7_75t_L g440 ( .A(n_295), .B(n_421), .Y(n_440) );
BUFx3_ASAP7_75t_L g638 ( .A(n_295), .Y(n_638) );
INVx2_ASAP7_75t_L g651 ( .A(n_295), .Y(n_651) );
BUFx3_ASAP7_75t_L g1438 ( .A(n_295), .Y(n_1438) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_296), .Y(n_305) );
INVx2_ASAP7_75t_L g312 ( .A(n_296), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_296), .B(n_304), .Y(n_317) );
AND2x4_ASAP7_75t_L g425 ( .A(n_296), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g525 ( .A(n_297), .Y(n_525) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_299), .A2(n_337), .B1(n_366), .B2(n_369), .Y(n_365) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_300), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_300), .A2(n_689), .B1(n_850), .B2(n_851), .C(n_852), .Y(n_849) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g517 ( .A(n_301), .B(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g653 ( .A(n_301), .Y(n_653) );
INVx4_ASAP7_75t_L g784 ( .A(n_301), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g1131 ( .A1(n_301), .A2(n_689), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_1131) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
BUFx2_ASAP7_75t_L g593 ( .A(n_302), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
BUFx2_ASAP7_75t_L g435 ( .A(n_303), .Y(n_435) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
BUFx2_ASAP7_75t_L g432 ( .A(n_305), .Y(n_432) );
INVx2_ASAP7_75t_L g542 ( .A(n_305), .Y(n_542) );
AND2x4_ASAP7_75t_L g570 ( .A(n_305), .B(n_551), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_313), .B2(n_314), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_307), .A2(n_321), .B1(n_356), .B2(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g1444 ( .A(n_308), .Y(n_1444) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g420 ( .A(n_309), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g939 ( .A(n_309), .Y(n_939) );
INVx2_ASAP7_75t_L g1134 ( .A(n_309), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g320 ( .A(n_310), .Y(n_320) );
BUFx8_ASAP7_75t_L g528 ( .A(n_310), .Y(n_528) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_310), .Y(n_568) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x4_ASAP7_75t_L g524 ( .A(n_312), .B(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_313), .A2(n_324), .B1(n_345), .B2(n_377), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_314), .A2(n_971), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g642 ( .A(n_315), .Y(n_642) );
INVx3_ASAP7_75t_L g857 ( .A(n_315), .Y(n_857) );
CKINVDCx8_ASAP7_75t_R g940 ( .A(n_315), .Y(n_940) );
INVx1_ASAP7_75t_L g1440 ( .A(n_315), .Y(n_1440) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g323 ( .A(n_316), .Y(n_323) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g443 ( .A(n_317), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B1(n_322), .B2(n_324), .Y(n_318) );
INVx2_ASAP7_75t_L g1375 ( .A(n_319), .Y(n_1375) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g645 ( .A(n_320), .Y(n_645) );
OR2x6_ASAP7_75t_SL g702 ( .A(n_320), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g962 ( .A(n_320), .Y(n_962) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g532 ( .A(n_323), .B(n_518), .Y(n_532) );
INVx1_ASAP7_75t_L g790 ( .A(n_323), .Y(n_790) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI33xp33_ASAP7_75t_L g558 ( .A1(n_326), .A2(n_559), .A3(n_561), .B1(n_565), .B2(n_571), .B3(n_573), .Y(n_558) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g1377 ( .A(n_327), .Y(n_1377) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx3_ASAP7_75t_L g648 ( .A(n_328), .Y(n_648) );
NAND3x1_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .C(n_332), .Y(n_328) );
INVx1_ASAP7_75t_L g421 ( .A(n_329), .Y(n_421) );
AND2x4_ASAP7_75t_L g424 ( .A(n_329), .B(n_425), .Y(n_424) );
OR2x6_ASAP7_75t_L g442 ( .A(n_329), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g544 ( .A(n_329), .B(n_545), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_329), .B(n_332), .Y(n_697) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g534 ( .A(n_331), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_331), .B(n_458), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_335), .A2(n_636), .B1(n_965), .B2(n_966), .Y(n_964) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_336), .A2(n_641), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g1445 ( .A1(n_336), .A2(n_638), .B1(n_696), .B2(n_1446), .C(n_1447), .Y(n_1445) );
OAI33xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_344), .A3(n_355), .B1(n_365), .B2(n_370), .B3(n_376), .Y(n_338) );
OAI33xp33_ASAP7_75t_L g1457 ( .A1(n_339), .A2(n_1458), .A3(n_1461), .B1(n_1464), .B2(n_1469), .B3(n_1470), .Y(n_1457) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g605 ( .A(n_340), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g740 ( .A1(n_340), .A2(n_741), .B1(n_744), .B2(n_745), .C1(n_754), .C2(n_760), .Y(n_740) );
INVx2_ASAP7_75t_L g813 ( .A(n_340), .Y(n_813) );
INVx4_ASAP7_75t_L g878 ( .A(n_340), .Y(n_878) );
AOI31xp33_ASAP7_75t_L g903 ( .A1(n_340), .A2(n_768), .A3(n_904), .B(n_905), .Y(n_903) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g716 ( .A(n_341), .Y(n_716) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_341), .B(n_697), .Y(n_1062) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g512 ( .A(n_342), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_342), .B(n_481), .Y(n_734) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g472 ( .A(n_348), .Y(n_472) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_348), .Y(n_816) );
BUFx3_ASAP7_75t_L g1471 ( .A(n_348), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_350), .A2(n_695), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx4_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g475 ( .A(n_351), .Y(n_475) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_351), .Y(n_614) );
INVx1_ASAP7_75t_L g630 ( .A(n_351), .Y(n_630) );
INVx2_ASAP7_75t_SL g759 ( .A(n_351), .Y(n_759) );
INVx2_ASAP7_75t_L g1463 ( .A(n_351), .Y(n_1463) );
INVx8_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g405 ( .A(n_352), .B(n_390), .Y(n_405) );
BUFx2_ASAP7_75t_L g818 ( .A(n_352), .Y(n_818) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g464 ( .A(n_357), .Y(n_464) );
BUFx2_ASAP7_75t_L g1466 ( .A(n_357), .Y(n_1466) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g368 ( .A(n_358), .Y(n_368) );
BUFx2_ASAP7_75t_L g619 ( .A(n_358), .Y(n_619) );
INVx1_ASAP7_75t_L g822 ( .A(n_358), .Y(n_822) );
BUFx2_ASAP7_75t_L g824 ( .A(n_358), .Y(n_824) );
AND2x2_ASAP7_75t_L g498 ( .A(n_359), .B(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g1118 ( .A(n_362), .Y(n_1118) );
INVx1_ASAP7_75t_L g1468 ( .A(n_362), .Y(n_1468) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_L g369 ( .A(n_363), .Y(n_369) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_363), .Y(n_381) );
OR2x6_ASAP7_75t_L g769 ( .A(n_363), .B(n_770), .Y(n_769) );
BUFx4f_ASAP7_75t_L g1159 ( .A(n_363), .Y(n_1159) );
BUFx4f_ASAP7_75t_L g1459 ( .A(n_363), .Y(n_1459) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g462 ( .A(n_364), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_366), .A2(n_1117), .B1(n_1118), .B2(n_1119), .C(n_1120), .Y(n_1116) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g1158 ( .A1(n_368), .A2(n_1133), .B1(n_1140), .B2(n_1159), .C(n_1160), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g603 ( .A1(n_370), .A2(n_604), .A3(n_606), .B1(n_615), .B2(n_621), .B3(n_624), .Y(n_603) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_SL g1157 ( .A1(n_372), .A2(n_813), .B1(n_1158), .B2(n_1161), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
AND2x4_ASAP7_75t_L g760 ( .A(n_373), .B(n_375), .Y(n_760) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx4_ASAP7_75t_L g494 ( .A(n_375), .Y(n_494) );
INVx4_ASAP7_75t_L g987 ( .A(n_375), .Y(n_987) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_377), .A2(n_471), .B1(n_963), .B2(n_972), .C(n_985), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_377), .A2(n_965), .B1(n_993), .B2(n_996), .C(n_997), .Y(n_992) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI31xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_398), .A3(n_406), .B(n_412), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_381), .A2(n_616), .B1(n_617), .B2(n_620), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_381), .A2(n_782), .B1(n_793), .B2(n_824), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_381), .A2(n_464), .B1(n_1132), .B2(n_1137), .C(n_1162), .Y(n_1161) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_385), .B(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g489 ( .A(n_385), .Y(n_489) );
AND2x6_ASAP7_75t_L g502 ( .A(n_385), .B(n_481), .Y(n_502) );
INVx1_ASAP7_75t_L g747 ( .A(n_385), .Y(n_747) );
BUFx3_ASAP7_75t_L g755 ( .A(n_385), .Y(n_755) );
BUFx3_ASAP7_75t_L g874 ( .A(n_385), .Y(n_874) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_385), .Y(n_1031) );
BUFx6f_ASAP7_75t_L g1390 ( .A(n_385), .Y(n_1390) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g919 ( .A(n_386), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_392), .B2(n_393), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_428), .B1(n_433), .B2(n_436), .Y(n_427) );
BUFx3_ASAP7_75t_L g659 ( .A(n_389), .Y(n_659) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g479 ( .A(n_391), .Y(n_479) );
INVx1_ASAP7_75t_L g736 ( .A(n_391), .Y(n_736) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_391), .Y(n_1025) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g662 ( .A(n_395), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_396), .B(n_481), .Y(n_516) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g665 ( .A(n_400), .Y(n_665) );
AND2x4_ASAP7_75t_L g409 ( .A(n_401), .B(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g667 ( .A(n_405), .Y(n_667) );
INVx3_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g669 ( .A(n_409), .Y(n_669) );
INVx2_ASAP7_75t_L g493 ( .A(n_410), .Y(n_493) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_410), .Y(n_509) );
BUFx3_ASAP7_75t_L g750 ( .A(n_410), .Y(n_750) );
OAI31xp33_ASAP7_75t_L g654 ( .A1(n_412), .A2(n_655), .A3(n_663), .B(n_668), .Y(n_654) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g515 ( .A(n_415), .B(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g557 ( .A(n_415), .Y(n_557) );
INVx1_ASAP7_75t_L g722 ( .A(n_415), .Y(n_722) );
OR2x2_ASAP7_75t_L g832 ( .A(n_415), .B(n_516), .Y(n_832) );
OAI31xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_422), .A3(n_437), .B(n_444), .Y(n_416) );
INVx2_ASAP7_75t_SL g588 ( .A(n_418), .Y(n_588) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g589 ( .A(n_420), .Y(n_589) );
CKINVDCx8_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g564 ( .A(n_425), .Y(n_564) );
BUFx2_ASAP7_75t_L g575 ( .A(n_425), .Y(n_575) );
AND2x2_ASAP7_75t_L g682 ( .A(n_425), .B(n_680), .Y(n_682) );
BUFx3_ASAP7_75t_L g931 ( .A(n_425), .Y(n_931) );
BUFx2_ASAP7_75t_L g974 ( .A(n_425), .Y(n_974) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_425), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_425), .Y(n_1098) );
INVx1_ASAP7_75t_L g551 ( .A(n_426), .Y(n_551) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g595 ( .A(n_429), .Y(n_595) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
AND2x4_ASAP7_75t_L g434 ( .A(n_430), .B(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_433), .A2(n_595), .B1(n_596), .B2(n_597), .Y(n_594) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g599 ( .A(n_440), .Y(n_599) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g601 ( .A(n_442), .Y(n_601) );
BUFx3_ASAP7_75t_L g646 ( .A(n_443), .Y(n_646) );
INVx1_ASAP7_75t_L g1054 ( .A(n_443), .Y(n_1054) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_448), .Y(n_445) );
AND2x4_ASAP7_75t_L g584 ( .A(n_446), .B(n_448), .Y(n_584) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_529), .C(n_537), .Y(n_451) );
O2A1O1Ixp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_482), .B(n_511), .C(n_513), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g983 ( .A(n_455), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_455), .A2(n_478), .B1(n_1370), .B2(n_1371), .Y(n_1413) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g484 ( .A(n_458), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g505 ( .A(n_458), .B(n_498), .Y(n_505) );
AND2x4_ASAP7_75t_L g508 ( .A(n_458), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g723 ( .A(n_458), .B(n_509), .Y(n_723) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_458), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_464), .B2(n_465), .C(n_466), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_460), .A2(n_617), .B1(n_622), .B2(n_623), .Y(n_621) );
INVx5_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g657 ( .A(n_462), .Y(n_657) );
OR2x2_ASAP7_75t_L g766 ( .A(n_462), .B(n_728), .Y(n_766) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_462), .B(n_728), .Y(n_1104) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g998 ( .A(n_468), .Y(n_998) );
INVx2_ASAP7_75t_L g1410 ( .A(n_468), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_473), .B2(n_476), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_471), .A2(n_791), .B1(n_818), .B2(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g1022 ( .A(n_480), .Y(n_1022) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_481), .B(n_498), .Y(n_535) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_481), .B(n_1025), .Y(n_1024) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g914 ( .A(n_485), .Y(n_914) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_485), .Y(n_1035) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g501 ( .A(n_486), .Y(n_501) );
INVx2_ASAP7_75t_L g730 ( .A(n_486), .Y(n_730) );
BUFx3_ASAP7_75t_L g907 ( .A(n_486), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_495), .B(n_502), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_489), .A2(n_501), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
A2O1A1Ixp33_ASAP7_75t_L g1018 ( .A1(n_489), .A2(n_1019), .B(n_1021), .C(n_1022), .Y(n_1018) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g916 ( .A(n_491), .Y(n_916) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_492), .Y(n_1409) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g1110 ( .A(n_493), .Y(n_1110) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g881 ( .A(n_497), .Y(n_881) );
INVx2_ASAP7_75t_L g1396 ( .A(n_497), .Y(n_1396) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_498), .Y(n_876) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g1397 ( .A(n_501), .Y(n_1397) );
INVx1_ASAP7_75t_L g988 ( .A(n_502), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g1387 ( .A1(n_502), .A2(n_1388), .B(n_1395), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_506), .B1(n_507), .B2(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g1000 ( .A(n_504), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g763 ( .A(n_505), .B(n_722), .Y(n_763) );
INVx1_ASAP7_75t_L g1401 ( .A(n_505), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_506), .A2(n_510), .B1(n_521), .B2(n_527), .Y(n_520) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_508), .Y(n_991) );
INVx1_ASAP7_75t_L g1404 ( .A(n_508), .Y(n_1404) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_509), .Y(n_873) );
INVx2_ASAP7_75t_L g1394 ( .A(n_509), .Y(n_1394) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g805 ( .A(n_512), .Y(n_805) );
OAI31xp33_ASAP7_75t_SL g839 ( .A1(n_512), .A2(n_840), .A3(n_844), .B(n_848), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_512), .A2(n_719), .B1(n_921), .B2(n_944), .Y(n_920) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
INVx2_ASAP7_75t_SL g738 ( .A(n_515), .Y(n_738) );
INVx1_ASAP7_75t_L g1027 ( .A(n_516), .Y(n_1027) );
INVx2_ASAP7_75t_L g1042 ( .A(n_517), .Y(n_1042) );
INVx1_ASAP7_75t_L g526 ( .A(n_518), .Y(n_526) );
INVx1_ASAP7_75t_L g977 ( .A(n_518), .Y(n_977) );
INVx1_ASAP7_75t_L g680 ( .A(n_519), .Y(n_680) );
INVx1_ASAP7_75t_L g704 ( .A(n_519), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_521), .B(n_1038), .Y(n_1037) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx8_ASAP7_75t_L g562 ( .A(n_523), .Y(n_562) );
INVx3_ASAP7_75t_L g574 ( .A(n_523), .Y(n_574) );
INVx2_ASAP7_75t_L g684 ( .A(n_523), .Y(n_684) );
INVx8_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_524), .B(n_544), .Y(n_556) );
AND2x2_ASAP7_75t_L g679 ( .A(n_524), .B(n_680), .Y(n_679) );
BUFx3_ASAP7_75t_L g798 ( .A(n_524), .Y(n_798) );
BUFx3_ASAP7_75t_L g1076 ( .A(n_524), .Y(n_1076) );
AND2x4_ASAP7_75t_L g527 ( .A(n_526), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g953 ( .A(n_527), .Y(n_953) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_528), .Y(n_572) );
INVx2_ASAP7_75t_SL g692 ( .A(n_528), .Y(n_692) );
INVx3_ASAP7_75t_L g851 ( .A(n_528), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_530), .A2(n_979), .B(n_980), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g1382 ( .A1(n_530), .A2(n_1383), .B(n_1384), .Y(n_1382) );
INVx8_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g898 ( .A(n_533), .Y(n_898) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x4_ASAP7_75t_L g543 ( .A(n_534), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g742 ( .A(n_534), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_535), .Y(n_743) );
AND4x1_ASAP7_75t_SL g537 ( .A(n_538), .B(n_552), .C(n_558), .D(n_576), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_546), .B2(n_547), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_540), .A2(n_547), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x6_ASAP7_75t_L g709 ( .A(n_541), .B(n_544), .Y(n_709) );
AND2x2_ASAP7_75t_L g956 ( .A(n_541), .B(n_543), .Y(n_956) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g547 ( .A(n_543), .B(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g577 ( .A(n_543), .B(n_564), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g1045 ( .A1(n_543), .A2(n_562), .B(n_1014), .C(n_1046), .Y(n_1045) );
AND2x2_ASAP7_75t_L g711 ( .A(n_544), .B(n_550), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_544), .Y(n_713) );
INVx1_ASAP7_75t_L g957 ( .A(n_547), .Y(n_957) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g700 ( .A(n_556), .Y(n_700) );
AOI33xp33_ASAP7_75t_L g1372 ( .A1(n_559), .A2(n_1373), .A3(n_1374), .B1(n_1376), .B2(n_1377), .B3(n_1378), .Y(n_1372) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_564), .A2(n_574), .B1(n_894), .B2(n_910), .Y(n_941) );
INVx8_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_567), .A2(n_1052), .B1(n_1053), .B2(n_1055), .Y(n_1051) );
INVx5_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g641 ( .A(n_568), .Y(n_641) );
INVx3_ASAP7_75t_L g971 ( .A(n_568), .Y(n_971) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_568), .Y(n_1083) );
BUFx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g685 ( .A(n_570), .Y(n_685) );
AND2x4_ASAP7_75t_L g706 ( .A(n_570), .B(n_704), .Y(n_706) );
BUFx12f_ASAP7_75t_L g929 ( .A(n_570), .Y(n_929) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_570), .Y(n_1077) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_577), .Y(n_1381) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_672), .B2(n_673), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g670 ( .A(n_582), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_602), .C(n_654), .Y(n_582) );
CKINVDCx14_ASAP7_75t_R g583 ( .A(n_584), .Y(n_583) );
NOR3xp33_ASAP7_75t_SL g585 ( .A(n_586), .B(n_590), .C(n_598), .Y(n_585) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x6_ASAP7_75t_L g712 ( .A(n_593), .B(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_596), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_632), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g1115 ( .A1(n_604), .A2(n_769), .B(n_1116), .Y(n_1115) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_612), .B2(n_613), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_607), .A2(n_622), .B1(n_636), .B2(n_639), .Y(n_635) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_610), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_612), .A2(n_623), .B1(n_650), .B2(n_652), .Y(n_649) );
INVx5_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx6_ASAP7_75t_L g1114 ( .A(n_614), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_616), .A2(n_628), .B1(n_641), .B2(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g1012 ( .A(n_618), .Y(n_1012) );
INVx4_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_620), .A2(n_631), .B1(n_644), .B2(n_646), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B1(n_629), .B2(n_631), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g1462 ( .A(n_626), .Y(n_1462) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx4_ASAP7_75t_L g753 ( .A(n_627), .Y(n_753) );
INVx3_ASAP7_75t_L g995 ( .A(n_627), .Y(n_995) );
BUFx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI33xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .A3(n_640), .B1(n_643), .B2(n_647), .B3(n_649), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI33xp33_ASAP7_75t_L g1047 ( .A1(n_634), .A2(n_1048), .A3(n_1051), .B1(n_1056), .B2(n_1059), .B3(n_1062), .Y(n_1047) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_638), .A2(n_696), .B1(n_783), .B2(n_859), .C(n_860), .Y(n_858) );
INVx2_ASAP7_75t_L g1080 ( .A(n_641), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_644), .A2(n_1053), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_645), .B(n_977), .Y(n_1041) );
INVx2_ASAP7_75t_L g1145 ( .A(n_645), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_646), .A2(n_960), .B1(n_961), .B2(n_963), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_646), .A2(n_968), .B1(n_969), .B2(n_972), .C(n_973), .Y(n_967) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g975 ( .A(n_650), .B(n_976), .Y(n_975) );
OR2x6_ASAP7_75t_L g1380 ( .A(n_650), .B(n_976), .Y(n_1380) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g855 ( .A(n_651), .Y(n_855) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g794 ( .A(n_653), .Y(n_794) );
INVx2_ASAP7_75t_L g1146 ( .A(n_653), .Y(n_1146) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_657), .A2(n_788), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_724), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_698), .B(n_714), .C(n_717), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_683), .C(n_690), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_679), .A2(n_682), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_684), .A2(n_1096), .B1(n_1097), .B2(n_1098), .Y(n_1095) );
OAI21xp33_ASAP7_75t_L g1435 ( .A1(n_689), .A2(n_851), .B(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_692), .A2(n_788), .B1(n_789), .B2(n_791), .Y(n_787) );
INVx3_ASAP7_75t_L g786 ( .A(n_696), .Y(n_786) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_700), .B(n_701), .C(n_707), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g725 ( .A1(n_699), .A2(n_726), .B1(n_731), .B2(n_737), .C1(n_738), .C2(n_739), .Y(n_725) );
AOI211xp5_ASAP7_75t_L g777 ( .A1(n_700), .A2(n_778), .B(n_779), .C(n_780), .Y(n_777) );
INVx2_ASAP7_75t_L g943 ( .A(n_700), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_700), .A2(n_1090), .B1(n_1092), .B2(n_1099), .Y(n_1089) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_700), .A2(n_936), .B1(n_1143), .B2(n_1144), .C(n_1149), .Y(n_1142) );
AOI211xp5_ASAP7_75t_L g1429 ( .A1(n_700), .A2(n_1430), .B(n_1431), .C(n_1432), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_702), .Y(n_800) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_704), .Y(n_937) );
INVx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g799 ( .A1(n_706), .A2(n_800), .B1(n_801), .B2(n_802), .C(n_803), .Y(n_799) );
INVx4_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_709), .A2(n_711), .B1(n_846), .B2(n_847), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_709), .A2(n_711), .B1(n_926), .B2(n_1087), .C(n_1088), .Y(n_1086) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_711), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_712), .Y(n_926) );
INVx1_ASAP7_75t_L g1448 ( .A(n_714), .Y(n_1448) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1001 ( .A(n_715), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1070 ( .A1(n_715), .A2(n_1071), .B(n_1100), .Y(n_1070) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI21xp5_ASAP7_75t_SL g1009 ( .A1(n_716), .A2(n_1010), .B(n_1029), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_721), .B(n_801), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_721), .B(n_867), .Y(n_866) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_721), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_721), .B(n_1454), .Y(n_1453) );
AND2x4_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_740), .C(n_761), .D(n_764), .Y(n_724) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_726), .A2(n_741), .B1(n_765), .B2(n_778), .C1(n_802), .C2(n_834), .Y(n_833) );
AOI21xp33_ASAP7_75t_L g868 ( .A1(n_726), .A2(n_869), .B(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_726), .A2(n_765), .B1(n_900), .B2(n_901), .Y(n_899) );
INVxp67_ASAP7_75t_L g1103 ( .A(n_726), .Y(n_1103) );
AOI222xp33_ASAP7_75t_L g1450 ( .A1(n_726), .A2(n_741), .B1(n_765), .B2(n_1430), .C1(n_1451), .C2(n_1452), .Y(n_1450) );
AND2x4_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
AOI332xp33_ASAP7_75t_L g1153 ( .A1(n_727), .A2(n_729), .A3(n_742), .B1(n_743), .B2(n_765), .B3(n_1143), .C1(n_1154), .C2(n_1155), .Y(n_1153) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_731), .A2(n_738), .B1(n_909), .B2(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_SL g831 ( .A(n_732), .Y(n_831) );
NAND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g770 ( .A(n_733), .Y(n_770) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
AOI332xp33_ASAP7_75t_L g871 ( .A1(n_741), .A2(n_760), .A3(n_872), .B1(n_875), .B2(n_877), .B3(n_879), .C1(n_880), .C2(n_882), .Y(n_871) );
AND2x4_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g986 ( .A(n_747), .Y(n_986) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_759), .A2(n_1441), .B1(n_1471), .B2(n_1472), .Y(n_1470) );
NAND3xp33_ASAP7_75t_L g911 ( .A(n_760), .B(n_912), .C(n_915), .Y(n_911) );
AOI211xp5_ASAP7_75t_L g1108 ( .A1(n_760), .A2(n_1109), .B(n_1115), .C(n_1121), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx3_ASAP7_75t_L g809 ( .A(n_763), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_763), .B(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_763), .B(n_1148), .Y(n_1151) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B(n_768), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_765), .A2(n_768), .B(n_847), .Y(n_865) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g1156 ( .A(n_768), .B(n_1157), .C(n_1163), .Y(n_1156) );
OR3x1_ASAP7_75t_L g1455 ( .A(n_768), .B(n_1456), .C(n_1457), .Y(n_1455) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g884 ( .A(n_772), .Y(n_884) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_836), .Y(n_773) );
OR2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_810), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_799), .B(n_804), .C(n_806), .Y(n_776) );
OAI21xp33_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_787), .B(n_792), .Y(n_780) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B(n_785), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_789), .A2(n_851), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI211xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B(n_795), .C(n_797), .Y(n_792) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_798), .Y(n_1085) );
INVx1_ASAP7_75t_L g1415 ( .A(n_804), .Y(n_1415) );
BUFx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_805), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_833), .C(n_835), .Y(n_810) );
NOR2xp33_ASAP7_75t_SL g811 ( .A(n_812), .B(n_829), .Y(n_811) );
OAI33xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .A3(n_819), .B1(n_823), .B2(n_825), .B3(n_827), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_814) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g1469 ( .A(n_828), .Y(n_1469) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_883), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_864), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_853), .B1(n_858), .B2(n_861), .Y(n_848) );
INVx1_ASAP7_75t_L g934 ( .A(n_851), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_853) );
NAND4xp25_ASAP7_75t_SL g864 ( .A(n_865), .B(n_866), .C(n_868), .D(n_871), .Y(n_864) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_876), .Y(n_906) );
INVx3_ASAP7_75t_L g1020 ( .A(n_876), .Y(n_1020) );
INVx2_ASAP7_75t_SL g877 ( .A(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_1064), .B1(n_1065), .B2(n_1165), .Y(n_885) );
INVx1_ASAP7_75t_L g1165 ( .A(n_886), .Y(n_1165) );
XNOR2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_946), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI21x1_ASAP7_75t_SL g889 ( .A1(n_890), .A2(n_891), .B(n_945), .Y(n_889) );
NAND4xp25_ASAP7_75t_L g945 ( .A(n_890), .B(n_893), .C(n_895), .D(n_920), .Y(n_945) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_895), .C(n_920), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_902), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_900), .A2(n_936), .B1(n_938), .B2(n_942), .Y(n_935) );
NAND3xp33_ASAP7_75t_SL g902 ( .A(n_903), .B(n_908), .C(n_911), .Y(n_902) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g1408 ( .A(n_918), .Y(n_1408) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_927), .C(n_935), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_926), .Y(n_922) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NOR3xp33_ASAP7_75t_L g1129 ( .A(n_926), .B(n_1130), .C(n_1135), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_930), .B1(n_932), .B2(n_933), .Y(n_927) );
BUFx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1091 ( .A(n_937), .Y(n_1091) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_1003), .B1(n_1004), .B2(n_1063), .Y(n_946) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
AND3x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_978), .C(n_981), .Y(n_949) );
AOI211xp5_ASAP7_75t_SL g950 ( .A1(n_951), .A2(n_952), .B(n_954), .C(n_958), .Y(n_950) );
INVxp67_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVxp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI31xp33_ASAP7_75t_L g981 ( .A1(n_982), .A2(n_989), .A3(n_999), .B(n_1001), .Y(n_981) );
INVxp67_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx2_ASAP7_75t_SL g994 ( .A(n_995), .Y(n_994) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_995), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1036), .Y(n_1008) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1016), .B(n_1017), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_1012), .A2(n_1436), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1023), .Y(n_1017) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_1024), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_1028), .A2(n_1040), .B1(n_1041), .B2(n_1042), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1032), .B1(n_1033), .B2(n_1034), .Y(n_1029) );
NAND3xp33_ASAP7_75t_SL g1036 ( .A(n_1037), .B(n_1039), .C(n_1043), .Y(n_1036) );
NOR2xp33_ASAP7_75t_SL g1043 ( .A(n_1044), .B(n_1047), .Y(n_1043) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_1054), .Y(n_1094) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B1(n_1124), .B2(n_1164), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
BUFx2_ASAP7_75t_SL g1067 ( .A(n_1068), .Y(n_1067) );
AOI21xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1122), .B(n_1123), .Y(n_1068) );
AND3x1_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1101), .C(n_1108), .Y(n_1069) );
AOI31xp33_ASAP7_75t_L g1123 ( .A1(n_1070), .A2(n_1101), .A3(n_1108), .B(n_1122), .Y(n_1123) );
NAND3xp33_ASAP7_75t_SL g1071 ( .A(n_1072), .B(n_1086), .C(n_1089), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1078), .B1(n_1081), .B2(n_1084), .Y(n_1072) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1076), .B(n_1148), .Y(n_1147) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx3_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1124), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
XNOR2x1_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1152), .Y(n_1127) );
A2O1A1Ixp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1142), .B(n_1150), .C(n_1151), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1361), .B1(n_1364), .B2(n_1416), .C(n_1422), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1303), .Y(n_1167) );
OAI32xp33_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1232), .A3(n_1264), .B1(n_1278), .B2(n_1293), .Y(n_1168) );
OAI311xp33_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1197), .A3(n_1202), .B1(n_1206), .C1(n_1225), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1187), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1171), .B(n_1288), .Y(n_1287) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_1172), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1172), .B(n_1239), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1172), .B(n_1224), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1172), .B(n_1259), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1172), .B(n_1241), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1344 ( .A(n_1172), .B(n_1255), .Y(n_1344) );
INVx4_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1209 ( .A(n_1173), .B(n_1210), .Y(n_1209) );
INVx4_ASAP7_75t_L g1229 ( .A(n_1173), .Y(n_1229) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1173), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1173), .B(n_1243), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1173), .B(n_1235), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1173), .B(n_1231), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_1173), .A2(n_1229), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1173), .B(n_1236), .Y(n_1320) );
NAND2xp5_ASAP7_75t_SL g1329 ( .A(n_1173), .B(n_1231), .Y(n_1329) );
AND2x4_ASAP7_75t_SL g1173 ( .A(n_1174), .B(n_1182), .Y(n_1173) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
AND2x6_ASAP7_75t_L g1180 ( .A(n_1176), .B(n_1181), .Y(n_1180) );
AND2x6_ASAP7_75t_L g1183 ( .A(n_1176), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1176), .B(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1176), .B(n_1186), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1176), .B(n_1186), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1176), .B(n_1177), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1180), .Y(n_1270) );
INVx2_ASAP7_75t_L g1363 ( .A(n_1183), .Y(n_1363) );
OAI21xp5_ASAP7_75t_L g1476 ( .A1(n_1184), .A2(n_1477), .B(n_1478), .Y(n_1476) );
AOI222xp33_ASAP7_75t_L g1284 ( .A1(n_1187), .A2(n_1285), .B1(n_1286), .B2(n_1289), .C1(n_1290), .C2(n_1291), .Y(n_1284) );
O2A1O1Ixp33_ASAP7_75t_SL g1323 ( .A1(n_1187), .A2(n_1320), .B(n_1324), .C(n_1330), .Y(n_1323) );
O2A1O1Ixp33_ASAP7_75t_L g1345 ( .A1(n_1187), .A2(n_1346), .B(n_1347), .C(n_1348), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_1188), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1188), .B(n_1223), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1193), .Y(n_1188) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1189), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1192), .Y(n_1189) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1193), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1193), .B(n_1237), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1193), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1194), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1194), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1197), .B(n_1253), .Y(n_1252) );
OAI211xp5_ASAP7_75t_L g1304 ( .A1(n_1197), .A2(n_1305), .B(n_1313), .C(n_1323), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1197), .B(n_1236), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1197), .B(n_1311), .Y(n_1355) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx3_ASAP7_75t_L g1223 ( .A(n_1198), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1198), .B(n_1237), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1198), .B(n_1285), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1198), .B(n_1237), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1200), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1202), .B(n_1211), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1202), .B(n_1230), .Y(n_1241) );
OAI21xp33_ASAP7_75t_L g1257 ( .A1(n_1202), .A2(n_1258), .B(n_1259), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1202), .B(n_1231), .Y(n_1279) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1203), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1203), .B(n_1211), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1203), .B(n_1261), .Y(n_1260) );
NAND2x1p5_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1205), .Y(n_1203) );
OAI21xp5_ASAP7_75t_SL g1206 ( .A1(n_1207), .A2(n_1214), .B(n_1221), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
NAND3xp33_ASAP7_75t_SL g1342 ( .A(n_1208), .B(n_1338), .C(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1209), .B(n_1216), .Y(n_1337) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1210), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1210), .B(n_1296), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1210), .B(n_1230), .Y(n_1325) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1211), .Y(n_1256) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1211), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1211), .B(n_1231), .Y(n_1288) );
OAI32xp33_ASAP7_75t_L g1353 ( .A1(n_1211), .A2(n_1240), .A3(n_1287), .B1(n_1292), .B2(n_1354), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1213), .Y(n_1211) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1215), .B(n_1280), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1219), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1216), .B(n_1260), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1216), .B(n_1235), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1217), .B(n_1218), .Y(n_1231) );
NOR2x1_ASAP7_75t_L g1228 ( .A(n_1219), .B(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1220), .B(n_1295), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1220), .B(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
CKINVDCx14_ASAP7_75t_R g1245 ( .A(n_1223), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1223), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1223), .B(n_1237), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1223), .B(n_1249), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1223), .B(n_1244), .Y(n_1358) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1224), .Y(n_1226) );
O2A1O1Ixp33_ASAP7_75t_L g1293 ( .A1(n_1224), .A2(n_1294), .B(n_1297), .C(n_1301), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
OAI21xp5_ASAP7_75t_L g1349 ( .A1(n_1227), .A2(n_1245), .B(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1230), .Y(n_1227) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1229), .B(n_1285), .Y(n_1309) );
CKINVDCx5p33_ASAP7_75t_R g1311 ( .A(n_1229), .Y(n_1311) );
O2A1O1Ixp33_ASAP7_75t_SL g1336 ( .A1(n_1229), .A2(n_1279), .B(n_1337), .C(n_1338), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1229), .B(n_1267), .Y(n_1360) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_1230), .A2(n_1233), .B1(n_1245), .B2(n_1246), .C(n_1250), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1230), .B(n_1235), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1230), .B(n_1260), .Y(n_1300) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1231), .B(n_1256), .Y(n_1255) );
AOI22xp5_ASAP7_75t_SL g1233 ( .A1(n_1234), .A2(n_1236), .B1(n_1238), .B2(n_1242), .Y(n_1233) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1234), .Y(n_1322) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1235), .Y(n_1308) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1236), .Y(n_1262) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1237), .Y(n_1277) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1237), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1237), .B(n_1244), .Y(n_1312) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_SL g1281 ( .A(n_1243), .B(n_1282), .Y(n_1281) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1244), .B(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1356 ( .A1(n_1247), .A2(n_1290), .B1(n_1298), .B2(n_1357), .Y(n_1356) );
O2A1O1Ixp33_ASAP7_75t_L g1352 ( .A1(n_1248), .A2(n_1298), .B(n_1315), .C(n_1353), .Y(n_1352) );
CKINVDCx5p33_ASAP7_75t_R g1248 ( .A(n_1249), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1254), .B1(n_1257), .B2(n_1262), .C(n_1263), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1253), .Y(n_1332) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_1256), .A2(n_1306), .B1(n_1309), .B2(n_1310), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1260), .B(n_1308), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1262), .B(n_1355), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1273), .Y(n_1263) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1264), .Y(n_1333) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .B1(n_1270), .B2(n_1271), .C(n_1272), .Y(n_1267) );
NAND3xp33_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1276), .C(n_1277), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1276), .B(n_1328), .Y(n_1347) );
OAI211xp5_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1280), .B(n_1281), .C(n_1284), .Y(n_1278) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1288), .Y(n_1290) );
CKINVDCx14_ASAP7_75t_R g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
AOI21xp5_ASAP7_75t_L g1330 ( .A1(n_1300), .A2(n_1331), .B(n_1332), .Y(n_1330) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1304), .A2(n_1333), .B(n_1334), .Y(n_1303) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1312), .Y(n_1310) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1312), .Y(n_1359) );
AOI211xp5_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1315), .B(n_1316), .C(n_1318), .Y(n_1313) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1314), .Y(n_1321) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1317), .Y(n_1346) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_1319), .A2(n_1321), .B(n_1322), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1326), .Y(n_1324) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NAND5xp2_ASAP7_75t_SL g1334 ( .A(n_1335), .B(n_1345), .C(n_1349), .D(n_1352), .E(n_1356), .Y(n_1334) );
OAI21xp5_ASAP7_75t_SL g1335 ( .A1(n_1336), .A2(n_1340), .B(n_1342), .Y(n_1335) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVxp67_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1347), .Y(n_1351) );
AOI21xp33_ASAP7_75t_L g1357 ( .A1(n_1358), .A2(n_1359), .B(n_1360), .Y(n_1357) );
CKINVDCx20_ASAP7_75t_R g1361 ( .A(n_1362), .Y(n_1361) );
CKINVDCx20_ASAP7_75t_R g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1382), .C(n_1385), .Y(n_1366) );
NOR3xp33_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1379), .C(n_1381), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1372), .Y(n_1368) );
OAI21xp5_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1405), .B(n_1414), .Y(n_1385) );
BUFx2_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .B1(n_1402), .B2(n_1403), .Y(n_1398) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1411), .Y(n_1406) );
INVx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
CKINVDCx20_ASAP7_75t_R g1416 ( .A(n_1417), .Y(n_1416) );
CKINVDCx20_ASAP7_75t_R g1417 ( .A(n_1418), .Y(n_1417) );
INVx3_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
BUFx3_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVxp33_ASAP7_75t_SL g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1426), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
AOI211x1_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1448), .B(n_1449), .C(n_1455), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1433), .Y(n_1428) );
NOR3xp33_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1442), .C(n_1443), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1437 ( .A1(n_1438), .A2(n_1439), .B1(n_1440), .B2(n_1441), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g1461 ( .A1(n_1439), .A2(n_1447), .B1(n_1462), .B2(n_1463), .Y(n_1461) );
OAI22xp5_ASAP7_75t_L g1464 ( .A1(n_1446), .A2(n_1465), .B1(n_1467), .B2(n_1468), .Y(n_1464) );
INVx4_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
endmodule