module fake_jpeg_3059_n_107 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_33),
.B1(n_30),
.B2(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_42),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_36),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_41),
.C(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_31),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_58),
.Y(n_69)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_52),
.B(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_42),
.B1(n_50),
.B2(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_53),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_49),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_50),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_15),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_31),
.B(n_29),
.C(n_34),
.D(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_29),
.B(n_38),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_1),
.B(n_3),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_16),
.B(n_28),
.C(n_25),
.D(n_23),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_32),
.C(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_49),
.B1(n_12),
.B2(n_13),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_82),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_1),
.B(n_3),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_4),
.B(n_6),
.Y(n_90)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_73),
.B1(n_81),
.B2(n_80),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_88),
.C(n_73),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_87),
.B(n_90),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_91),
.C(n_9),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_97),
.C(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_93),
.C(n_18),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_17),
.C(n_21),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_11),
.B(n_19),
.C(n_20),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_22),
.A3(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_10),
.Y(n_107)
);


endmodule