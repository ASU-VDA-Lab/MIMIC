module fake_ariane_273_n_3945 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_3945);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_3945;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2680;
wire n_2334;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_690;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_524;
wire n_2731;
wire n_3703;
wire n_634;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_520;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2663;
wire n_559;
wire n_2233;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2391;
wire n_2332;
wire n_3828;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3883;
wire n_1013;
wire n_3571;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_533;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_440;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_3739;
wire n_512;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_490;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_575;
wire n_546;
wire n_3472;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2326;
wire n_2145;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_3234;
wire n_3280;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_1179;
wire n_468;
wire n_3284;
wire n_3909;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_3678;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_3937;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_615;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_3891;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3724;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_3257;
wire n_477;
wire n_650;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3912;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2695;
wire n_2557;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3727;
wire n_3700;
wire n_712;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_489;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_3884;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_479;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3179;
wire n_2262;
wire n_3031;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_706;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_441;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3876;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_487;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_502;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_3599;
wire n_3618;
wire n_604;
wire n_439;
wire n_677;
wire n_3705;
wire n_3022;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_681;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_707;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_699;
wire n_1726;
wire n_2075;
wire n_3263;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3835;
wire n_3837;
wire n_3569;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_3819;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_887;
wire n_729;
wire n_3403;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_527;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2949;
wire n_2300;
wire n_2894;
wire n_3896;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_551;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3924;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_2893;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3617;
wire n_3459;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_3340;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2468;
wire n_2171;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3836;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_3097;
wire n_624;
wire n_3507;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_3864;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_480;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_730;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2723;
wire n_3925;
wire n_2928;
wire n_1118;
wire n_943;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2353;
wire n_2064;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_686;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_3718;
wire n_756;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2890;
wire n_515;
wire n_3381;
wire n_807;
wire n_3455;
wire n_3736;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3605;
wire n_3345;
wire n_2170;
wire n_3560;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_3809;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_2044;
wire n_928;
wire n_3886;
wire n_1153;
wire n_465;
wire n_3769;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_689;
wire n_1116;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_467;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3731;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2431;
wire n_2110;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3322;
wire n_2666;
wire n_3289;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2935;
wire n_2401;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_617;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_543;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_3790;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_3288;
wire n_3251;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_2371;
wire n_1978;
wire n_571;
wire n_3880;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_532;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_2315;
wire n_1857;
wire n_3926;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3807;
wire n_580;
wire n_3664;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_923;
wire n_1645;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_1564;
wire n_2010;
wire n_3677;
wire n_1054;
wire n_508;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_2425;
wire n_1952;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3576;
wire n_3558;
wire n_3782;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_679;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_443;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_761;
wire n_733;
wire n_2212;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_2897;
wire n_816;
wire n_1322;
wire n_3273;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_2580;
wire n_485;
wire n_1792;
wire n_504;
wire n_3351;
wire n_2062;
wire n_483;
wire n_435;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_3933;
wire n_778;
wire n_1619;
wire n_2351;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_3232;
wire n_3001;
wire n_3188;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2447;
wire n_1845;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_671;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1409;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_488;
wire n_3018;
wire n_904;
wire n_505;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_498;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_3874;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_459;
wire n_1136;
wire n_2515;
wire n_3845;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_448;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_450;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_3918;
wire n_716;
wire n_1571;
wire n_1698;
wire n_3902;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_656;
wire n_492;
wire n_574;
wire n_3593;
wire n_2673;
wire n_664;
wire n_2585;
wire n_1591;
wire n_2995;
wire n_3293;
wire n_3361;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2485;
wire n_2052;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_537;
wire n_1063;
wire n_3934;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_1581;
wire n_3849;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3592;
wire n_3725;
wire n_3557;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3075;
wire n_3030;
wire n_3505;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_3771;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_548;
wire n_3427;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_457;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_3041;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2423;
wire n_2689;
wire n_2208;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_796;
wire n_573;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_76),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_38),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_212),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_45),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_175),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_148),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_283),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_147),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_14),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_21),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_97),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_272),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_87),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_303),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_89),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_366),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_92),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_284),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_338),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_289),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_107),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_424),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_206),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_35),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_2),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_22),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_101),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_129),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_60),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_165),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_211),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_96),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_341),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_21),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_175),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_141),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_351),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_297),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_405),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_6),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_232),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_153),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_120),
.Y(n_481)
);

BUFx8_ASAP7_75t_SL g482 ( 
.A(n_234),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_365),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_59),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_411),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_99),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_332),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_336),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_157),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_325),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_54),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_310),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_209),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_38),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_308),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_213),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_0),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_222),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_81),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_348),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_147),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_378),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_322),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_250),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_134),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_350),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_211),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_339),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_307),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_287),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_131),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_91),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_232),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_62),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_181),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_68),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_359),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_237),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_26),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_188),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_357),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_304),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_214),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_166),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_145),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_180),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_394),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_174),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_179),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_73),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_407),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_104),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_216),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_160),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_306),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_395),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_10),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_295),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_401),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_387),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_126),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_62),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_115),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_10),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_103),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_337),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_314),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_404),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_247),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_227),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_2),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_108),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_0),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_116),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_47),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_61),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_305),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_301),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_421),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_419),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_431),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_225),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_75),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_121),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_191),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_317),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_98),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_224),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_209),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_326),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_290),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_271),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_37),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_137),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_330),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_110),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_358),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_275),
.Y(n_580)
);

BUFx5_ASAP7_75t_L g581 ( 
.A(n_106),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_364),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_418),
.Y(n_583)
);

BUFx5_ASAP7_75t_L g584 ( 
.A(n_73),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_68),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_114),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_52),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_67),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_155),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_381),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_128),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_300),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_344),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_334),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_375),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_195),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_374),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_66),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_76),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_53),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_118),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_247),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_225),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_296),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_414),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_131),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_320),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_353),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_346),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_19),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_113),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_91),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_288),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_183),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_64),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_133),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_134),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_177),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_161),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_328),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_390),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_221),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_93),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_208),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_135),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_192),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_24),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_195),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_158),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_420),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_273),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_258),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_57),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_252),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_61),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_210),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_367),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_1),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_51),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_377),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_302),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_48),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_389),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_283),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_272),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_368),
.Y(n_646)
);

BUFx2_ASAP7_75t_SL g647 ( 
.A(n_132),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_202),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_142),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_107),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_169),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_114),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_7),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_159),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_3),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_149),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_16),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_396),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_267),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_224),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_34),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_28),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_39),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_160),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_15),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_220),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_355),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_423),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_82),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_201),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_333),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_120),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_78),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_267),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_33),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_415),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_260),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_53),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_281),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_196),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_356),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_388),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_244),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_417),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_110),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_383),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_371),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_117),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_20),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_309),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_122),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_240),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_241),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_203),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_379),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_60),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_369),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_98),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_429),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_130),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_240),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_56),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_88),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_170),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_65),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_362),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_158),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_163),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_352),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_292),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_79),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_312),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_163),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_342),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_127),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_249),
.Y(n_716)
);

BUFx2_ASAP7_75t_SL g717 ( 
.A(n_165),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_86),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_5),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_74),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_422),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_208),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_201),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_96),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_79),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_174),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_277),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_210),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_360),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_139),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_194),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_159),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_103),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_188),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_48),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_261),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_218),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_428),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_275),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_59),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_241),
.Y(n_741)
);

BUFx5_ASAP7_75t_L g742 ( 
.A(n_324),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_8),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_81),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_70),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_363),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_287),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_581),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_468),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_569),
.Y(n_752)
);

INVxp67_ASAP7_75t_SL g753 ( 
.A(n_552),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_482),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_558),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_581),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_581),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_450),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_452),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_581),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_495),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_538),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_597),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_604),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_605),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_581),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_681),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_439),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_466),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_584),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_584),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_439),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_625),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_491),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_584),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_584),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_625),
.Y(n_779)
);

INVxp33_ASAP7_75t_SL g780 ( 
.A(n_574),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_584),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_544),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_434),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_584),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_584),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_435),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_551),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_584),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_507),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_450),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_438),
.Y(n_791)
);

CKINVDCx14_ASAP7_75t_R g792 ( 
.A(n_540),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_734),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_564),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_564),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_447),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_509),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_448),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_453),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_458),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_540),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_584),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_552),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_436),
.B(n_1),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_747),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_444),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_444),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_457),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_457),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_459),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_459),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_478),
.Y(n_813)
);

CKINVDCx16_ASAP7_75t_R g814 ( 
.A(n_507),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_462),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_464),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_478),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_507),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_487),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_465),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_467),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_461),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_469),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_487),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_521),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_471),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_521),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_534),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_473),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_534),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_537),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_608),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_537),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_559),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_559),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_563),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_563),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_583),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_583),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_480),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_608),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_450),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_590),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_590),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_461),
.Y(n_846)
);

INVxp33_ASAP7_75t_L g847 ( 
.A(n_440),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_461),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_592),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_592),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_451),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_595),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_595),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_494),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_461),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_637),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_489),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_607),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_607),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_613),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_613),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_499),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_556),
.Y(n_863)
);

BUFx10_ASAP7_75t_L g864 ( 
.A(n_461),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_637),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_501),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_630),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_637),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_630),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_450),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_504),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_640),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_647),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_505),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_507),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_640),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_511),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_516),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_519),
.Y(n_879)
);

INVxp33_ASAP7_75t_L g880 ( 
.A(n_440),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_641),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_524),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_526),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_531),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_488),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_727),
.Y(n_886)
);

CKINVDCx14_ASAP7_75t_R g887 ( 
.A(n_488),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_641),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_643),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_643),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_717),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_533),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_658),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_535),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_658),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_667),
.Y(n_896)
);

BUFx10_ASAP7_75t_L g897 ( 
.A(n_461),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_667),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_682),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_536),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_539),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_543),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_488),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_727),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_682),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_697),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_697),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_545),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_699),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_699),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_709),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_709),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_547),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_712),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_554),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_555),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_712),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_474),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_437),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_437),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_488),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_474),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_565),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_437),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_493),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_566),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_493),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_575),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_578),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_474),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_493),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_738),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_497),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_497),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_727),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_497),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_580),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_510),
.Y(n_938)
);

CKINVDCx14_ASAP7_75t_R g939 ( 
.A(n_738),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_738),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_510),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_585),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_510),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_621),
.B(n_3),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_496),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_586),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_525),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_738),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_525),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_587),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_450),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_589),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_485),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_525),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_527),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_527),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_591),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_599),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_717),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_527),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_600),
.Y(n_961)
);

CKINVDCx14_ASAP7_75t_R g962 ( 
.A(n_746),
.Y(n_962)
);

CKINVDCx14_ASAP7_75t_R g963 ( 
.A(n_443),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_530),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_530),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_601),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_530),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_496),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_606),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_603),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_606),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_606),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_619),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_619),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_610),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_612),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_485),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_614),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_615),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_619),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_622),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_645),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_645),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_485),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_623),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_645),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_523),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_496),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_496),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_496),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_496),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_661),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_669),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_669),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_624),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_669),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_669),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_669),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_450),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_441),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_669),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_719),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_719),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_719),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_627),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_628),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_523),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_719),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_629),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_631),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_632),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_719),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_719),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_436),
.B(n_4),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_523),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_745),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_441),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_633),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_634),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_572),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_442),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_445),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_635),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_445),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_636),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_446),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_446),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_638),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_639),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_454),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_644),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_572),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_648),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_454),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_460),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_649),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_460),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_572),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_650),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_472),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_651),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_652),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_472),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_479),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_479),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_654),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_655),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_656),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_659),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_660),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_481),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_481),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_664),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_498),
.Y(n_1054)
);

CKINVDCx14_ASAP7_75t_R g1055 ( 
.A(n_449),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_665),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_498),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_512),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_666),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_512),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_513),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_742),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_670),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_513),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_514),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_673),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_514),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_477),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_742),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_677),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_679),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_518),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_518),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_520),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_477),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_520),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_680),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_621),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_553),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_553),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_486),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_557),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_557),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_683),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_567),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_685),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_742),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_692),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_742),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_695),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_742),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_695),
.B(n_4),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_567),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_689),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_455),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_770),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_776),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1015),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_855),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_787),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_864),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_789),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1015),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_759),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_761),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_918),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_763),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_793),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_764),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_765),
.Y(n_1110)
);

INVxp33_ASAP7_75t_SL g1111 ( 
.A(n_755),
.Y(n_1111)
);

INVxp67_ASAP7_75t_SL g1112 ( 
.A(n_918),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_762),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_767),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_754),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_855),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1020),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_782),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1020),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_L g1120 ( 
.A(n_807),
.B(n_456),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_751),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1032),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_752),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_806),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_885),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1032),
.Y(n_1126)
);

CKINVDCx16_ASAP7_75t_R g1127 ( 
.A(n_814),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_922),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_783),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1032),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_932),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1032),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_786),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_948),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1032),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_922),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_791),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_748),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_887),
.B(n_475),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_978),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_748),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1095),
.B(n_710),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_930),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_985),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_796),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_799),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_800),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1006),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1095),
.B(n_710),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_750),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_750),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_930),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_801),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_1023),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1025),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_815),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_756),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_756),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_816),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_820),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_757),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_757),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_760),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_760),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_821),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_851),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_823),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_826),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_864),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_829),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_841),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_766),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_766),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_768),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_962),
.B(n_562),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_768),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_771),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_857),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_L g1179 ( 
.A(n_862),
.B(n_470),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_771),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_772),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_866),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_871),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_863),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_772),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1036),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_773),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1039),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_874),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_773),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_777),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_877),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_992),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_855),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1084),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_792),
.B(n_847),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_878),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_879),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_880),
.B(n_486),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_777),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1088),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_903),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_939),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_882),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_883),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_884),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_778),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_892),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_778),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_769),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_894),
.B(n_476),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_921),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_784),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_784),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_R g1215 ( 
.A(n_774),
.B(n_691),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_900),
.B(n_483),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_775),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_785),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_785),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_818),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_953),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_788),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_901),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_940),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_788),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_803),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_803),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_856),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_988),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_988),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_902),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_908),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_913),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_915),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_865),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_953),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_989),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_779),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_807),
.B(n_490),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_916),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_963),
.B(n_687),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1013),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_989),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_990),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_875),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_854),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_990),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1055),
.B(n_492),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_991),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_991),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_942),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_957),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_977),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_923),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_842),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_926),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_993),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1022),
.B(n_500),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_928),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_929),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_981),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_993),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_937),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_946),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_950),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_952),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1068),
.B(n_502),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_994),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_864),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_958),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_994),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_996),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1075),
.B(n_503),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_961),
.B(n_506),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_966),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_970),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_996),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_975),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_976),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_979),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_995),
.Y(n_1281)
);

CKINVDCx16_ASAP7_75t_R g1282 ( 
.A(n_802),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1005),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1009),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1010),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_802),
.B(n_832),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1011),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1018),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1019),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_977),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1028),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1029),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_753),
.B(n_508),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1031),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_984),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1013),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1033),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1041),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_997),
.Y(n_1299)
);

INVxp33_ASAP7_75t_SL g1300 ( 
.A(n_1042),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1046),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1047),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1048),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1049),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_897),
.Y(n_1305)
);

INVxp33_ASAP7_75t_SL g1306 ( 
.A(n_1050),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_997),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_998),
.Y(n_1308)
);

INVxp33_ASAP7_75t_SL g1309 ( 
.A(n_1053),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1056),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1059),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_998),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1002),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1063),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1066),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1070),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1071),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1002),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1003),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1013),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1003),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1077),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1086),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_984),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1004),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1004),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1094),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1008),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1008),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1012),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_868),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_832),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_987),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_987),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1013),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1012),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_868),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_797),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_797),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_797),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_749),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_749),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_781),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1024),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_839),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_781),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_873),
.B(n_517),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_919),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_780),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_919),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_891),
.Y(n_1351)
);

CKINVDCx16_ASAP7_75t_R g1352 ( 
.A(n_1024),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1007),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_794),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1078),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1081),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_920),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_920),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1078),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1090),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1007),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1090),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1038),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_804),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_804),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1081),
.Y(n_1366)
);

XOR2xp5_ASAP7_75t_L g1367 ( 
.A(n_944),
.B(n_693),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_935),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_959),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_795),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_798),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_808),
.B(n_522),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1013),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1038),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1092),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_924),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_897),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_925),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_897),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_925),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_886),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_927),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_904),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_927),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1341),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1341),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1355),
.B(n_805),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1383),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1295),
.B(n_808),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1184),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1331),
.B(n_1337),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1201),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1342),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1342),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1139),
.B(n_809),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1166),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1178),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1383),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1196),
.B(n_1000),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1099),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1375),
.A2(n_529),
.B1(n_700),
.B2(n_463),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1193),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1258),
.A2(n_1273),
.B1(n_1267),
.B2(n_1251),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1101),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1343),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1343),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1371),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1101),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1346),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1346),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1099),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1370),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1106),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1199),
.B(n_1017),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1142),
.A2(n_1149),
.B1(n_1286),
.B2(n_1241),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1381),
.B(n_1021),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1295),
.B(n_809),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1112),
.B(n_810),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1169),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1116),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1199),
.B(n_1017),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1128),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1136),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1169),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1229),
.A2(n_1069),
.B(n_1062),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1255),
.A2(n_515),
.B1(n_618),
.B2(n_484),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1102),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1116),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1104),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1143),
.B(n_1152),
.Y(n_1431)
);

NOR2x1_ASAP7_75t_L g1432 ( 
.A(n_1175),
.B(n_812),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1368),
.B(n_810),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1221),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1194),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1366),
.B(n_1026),
.Y(n_1436)
);

AOI22x1_ASAP7_75t_SL g1437 ( 
.A1(n_1144),
.A2(n_515),
.B1(n_618),
.B2(n_484),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1236),
.Y(n_1439)
);

OAI22x1_ASAP7_75t_SL g1440 ( 
.A1(n_1148),
.A2(n_694),
.B1(n_702),
.B2(n_698),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1194),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1138),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_L g1443 ( 
.A(n_1248),
.B(n_811),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1138),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1229),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1141),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1253),
.B(n_1027),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1129),
.B(n_1044),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1141),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1150),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1150),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1151),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1344),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1290),
.B(n_1079),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1344),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1230),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1324),
.B(n_1026),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1230),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1151),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1237),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1237),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1157),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1333),
.B(n_812),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1157),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1158),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1158),
.Y(n_1466)
);

XNOR2xp5_ASAP7_75t_L g1467 ( 
.A(n_1367),
.B(n_1096),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1334),
.B(n_813),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1161),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1161),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1243),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1162),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1293),
.B(n_813),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1362),
.B(n_1030),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1162),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1243),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1352),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1163),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1163),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_SL g1480 ( 
.A(n_1300),
.B(n_1014),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1133),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1164),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1282),
.B(n_817),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1244),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1244),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1164),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1172),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1172),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1353),
.B(n_1030),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1173),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1247),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1173),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1361),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1332),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1363),
.B(n_1034),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1348),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1348),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1174),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1174),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1367),
.A2(n_704),
.B1(n_707),
.B2(n_705),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1269),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1377),
.B(n_817),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1379),
.B(n_819),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1176),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1120),
.B(n_1034),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1154),
.A2(n_708),
.B1(n_715),
.B2(n_711),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1352),
.B(n_1035),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1176),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1269),
.B(n_819),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1177),
.Y(n_1510)
);

BUFx8_ASAP7_75t_L g1511 ( 
.A(n_1140),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1350),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1177),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1356),
.B(n_1035),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1305),
.B(n_824),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1350),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1133),
.B(n_824),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1180),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1356),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1247),
.A2(n_1069),
.B(n_1062),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1249),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1282),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1097),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1305),
.B(n_825),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1246),
.A2(n_713),
.B1(n_723),
.B2(n_720),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1120),
.B(n_1037),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1180),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1133),
.B(n_825),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1239),
.B(n_1037),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1105),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1181),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1357),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1252),
.A2(n_736),
.B1(n_740),
.B2(n_735),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1261),
.A2(n_743),
.B1(n_744),
.B2(n_741),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1249),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1354),
.B(n_1040),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1100),
.Y(n_1537)
);

AND2x2_ASAP7_75t_SL g1538 ( 
.A(n_1102),
.B(n_827),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1181),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1155),
.A2(n_728),
.B1(n_730),
.B2(n_546),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1185),
.Y(n_1541)
);

NOR2x1_ASAP7_75t_L g1542 ( 
.A(n_1179),
.B(n_827),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1357),
.B(n_1040),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1250),
.A2(n_1089),
.B(n_1087),
.Y(n_1544)
);

INVx6_ASAP7_75t_L g1545 ( 
.A(n_1133),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1280),
.B(n_828),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1250),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1239),
.B(n_1043),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1107),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1211),
.B(n_828),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1303),
.B(n_830),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1358),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1349),
.A2(n_831),
.B1(n_833),
.B2(n_830),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1372),
.B(n_1185),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1372),
.B(n_831),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1187),
.B(n_833),
.Y(n_1556)
);

INVx6_ASAP7_75t_L g1557 ( 
.A(n_1127),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1109),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1187),
.B(n_834),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1127),
.B(n_974),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1110),
.Y(n_1561)
);

AND2x6_ASAP7_75t_L g1562 ( 
.A(n_1122),
.B(n_834),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1115),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1374),
.B(n_1043),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1190),
.A2(n_1089),
.B(n_1087),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1140),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1376),
.B(n_1045),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1376),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1378),
.B(n_1045),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1190),
.B(n_835),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1191),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1380),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1191),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1345),
.A2(n_1351),
.B1(n_1369),
.B2(n_1215),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1380),
.B(n_1051),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1200),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1200),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1207),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1207),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1209),
.B(n_836),
.Y(n_1580)
);

CKINVDCx6p67_ASAP7_75t_R g1581 ( 
.A(n_1260),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1257),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1257),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1262),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1186),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1382),
.B(n_1051),
.Y(n_1586)
);

BUFx8_ASAP7_75t_L g1587 ( 
.A(n_1186),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1216),
.B(n_837),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1306),
.A2(n_1309),
.B1(n_1145),
.B2(n_1146),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1209),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1213),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1262),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1304),
.B(n_838),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1263),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1213),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1214),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1214),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1268),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1265),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_L g1600 ( 
.A(n_1218),
.B(n_742),
.Y(n_1600)
);

AND2x6_ASAP7_75t_L g1601 ( 
.A(n_1122),
.B(n_838),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1270),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1114),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1268),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1218),
.Y(n_1605)
);

OAI22x1_ASAP7_75t_R g1606 ( 
.A1(n_1275),
.A2(n_571),
.B1(n_576),
.B2(n_570),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1271),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1271),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1279),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1219),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1272),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1382),
.B(n_1052),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1272),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1219),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1277),
.A2(n_1091),
.B(n_844),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1384),
.B(n_1052),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1384),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1188),
.A2(n_571),
.B1(n_576),
.B2(n_570),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1222),
.A2(n_1091),
.B(n_844),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1222),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1098),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1277),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1225),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1347),
.B(n_1054),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1225),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1226),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1226),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1299),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1227),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1108),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1291),
.B(n_1054),
.Y(n_1631)
);

XNOR2x2_ASAP7_75t_L g1632 ( 
.A(n_1338),
.B(n_588),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1299),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1227),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1307),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1126),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1291),
.B(n_1057),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1126),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1130),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1130),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1203),
.B(n_1057),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1285),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1098),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1297),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1137),
.A2(n_596),
.B1(n_598),
.B2(n_588),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1274),
.B(n_1103),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1308),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1240),
.B(n_840),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1103),
.B(n_840),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1117),
.B(n_845),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1119),
.B(n_845),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1195),
.A2(n_598),
.B1(n_602),
.B2(n_596),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1119),
.B(n_1058),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1278),
.B(n_1060),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1322),
.B(n_1060),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1312),
.A2(n_850),
.B(n_849),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1313),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1313),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1132),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1415),
.A2(n_1339),
.B1(n_1340),
.B2(n_1220),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1480),
.A2(n_1153),
.B1(n_1156),
.B2(n_1147),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1596),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1663)
);

AO22x2_ASAP7_75t_L g1664 ( 
.A1(n_1437),
.A2(n_1235),
.B1(n_1228),
.B2(n_1113),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1557),
.B(n_1238),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1596),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1403),
.A2(n_1160),
.B1(n_1165),
.B2(n_1159),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1390),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1392),
.B(n_1238),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1631),
.B(n_1167),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1405),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1436),
.B(n_1118),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1557),
.B(n_1210),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1436),
.B(n_1124),
.Y(n_1674)
);

AO22x2_ASAP7_75t_L g1675 ( 
.A1(n_1437),
.A2(n_1202),
.B1(n_1224),
.B2(n_1212),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1676)
);

INVx8_ASAP7_75t_L g1677 ( 
.A(n_1481),
.Y(n_1677)
);

OAI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1553),
.A2(n_1170),
.B1(n_1171),
.B2(n_1168),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1500),
.A2(n_1301),
.B1(n_1314),
.B2(n_1298),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1395),
.A2(n_849),
.B1(n_852),
.B2(n_850),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1405),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_R g1683 ( 
.A1(n_1546),
.A2(n_611),
.B1(n_616),
.B2(n_602),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1557),
.B(n_1217),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1397),
.B(n_1430),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1445),
.Y(n_1686)
);

AO22x2_ASAP7_75t_L g1687 ( 
.A1(n_1401),
.A2(n_1645),
.B1(n_1606),
.B2(n_1632),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1445),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1473),
.A2(n_852),
.B1(n_858),
.B2(n_853),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1631),
.A2(n_1637),
.B1(n_1562),
.B2(n_1601),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1402),
.B(n_1220),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1402),
.B(n_1182),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1456),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1456),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1433),
.B(n_1183),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1631),
.A2(n_853),
.B1(n_859),
.B2(n_858),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1458),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1396),
.B(n_1189),
.Y(n_1698)
);

OAI22xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1637),
.A2(n_1197),
.B1(n_1198),
.B2(n_1192),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1637),
.A2(n_1205),
.B1(n_1206),
.B2(n_1204),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1562),
.A2(n_859),
.B1(n_861),
.B2(n_860),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1557),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1523),
.A2(n_1323),
.B1(n_1327),
.B2(n_1317),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1458),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1405),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1399),
.B(n_1208),
.Y(n_1706)
);

AO22x2_ASAP7_75t_L g1707 ( 
.A1(n_1632),
.A2(n_974),
.B1(n_861),
.B2(n_867),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1624),
.A2(n_1223),
.B1(n_1232),
.B2(n_1231),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1399),
.B(n_1233),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1460),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1519),
.B(n_1234),
.Y(n_1711)
);

XNOR2xp5_ASAP7_75t_L g1712 ( 
.A(n_1467),
.B(n_1121),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1564),
.A2(n_1503),
.B1(n_1502),
.B2(n_1654),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1624),
.A2(n_1254),
.B1(n_1259),
.B2(n_1256),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1624),
.A2(n_1264),
.B1(n_1276),
.B2(n_1266),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1564),
.A2(n_1283),
.B1(n_1284),
.B2(n_1281),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1551),
.B(n_1287),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1648),
.A2(n_1288),
.B1(n_1292),
.B2(n_1289),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1405),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1474),
.A2(n_1294),
.B1(n_1310),
.B2(n_1302),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1562),
.A2(n_860),
.B1(n_869),
.B2(n_867),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1399),
.B(n_1311),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1562),
.A2(n_1601),
.B1(n_1538),
.B2(n_1526),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1562),
.A2(n_869),
.B1(n_876),
.B2(n_872),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1562),
.A2(n_872),
.B1(n_881),
.B2(n_876),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1601),
.A2(n_881),
.B1(n_889),
.B2(n_888),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1601),
.A2(n_888),
.B1(n_890),
.B2(n_889),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1405),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1391),
.B(n_1315),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1601),
.A2(n_890),
.B1(n_895),
.B2(n_893),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1564),
.B(n_1316),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1601),
.A2(n_893),
.B1(n_896),
.B2(n_895),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1538),
.A2(n_896),
.B1(n_899),
.B2(n_898),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1461),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1483),
.B(n_1125),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1483),
.B(n_1536),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1589),
.A2(n_906),
.B1(n_907),
.B2(n_905),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1429),
.A2(n_907),
.B1(n_909),
.B2(n_906),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1461),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1569),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1471),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1523),
.A2(n_1123),
.B1(n_1134),
.B2(n_1131),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1505),
.A2(n_909),
.B1(n_911),
.B2(n_910),
.Y(n_1743)
);

AO22x2_ASAP7_75t_L g1744 ( 
.A1(n_1525),
.A2(n_911),
.B1(n_912),
.B2(n_910),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1471),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1429),
.A2(n_914),
.B1(n_917),
.B2(n_912),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1519),
.B(n_1061),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1476),
.Y(n_1748)
);

OAI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1530),
.A2(n_917),
.B1(n_914),
.B2(n_1111),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1476),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1545),
.A2(n_616),
.B1(n_617),
.B2(n_611),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1654),
.A2(n_626),
.B1(n_642),
.B2(n_617),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1505),
.A2(n_646),
.B1(n_1135),
.B2(n_1132),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1536),
.B(n_1245),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1505),
.A2(n_1135),
.B1(n_1319),
.B2(n_1318),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1545),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1618),
.A2(n_657),
.B1(n_662),
.B2(n_653),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1593),
.A2(n_662),
.B1(n_663),
.B2(n_657),
.Y(n_1758)
);

OAI22xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1655),
.A2(n_672),
.B1(n_674),
.B2(n_663),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1549),
.A2(n_674),
.B1(n_678),
.B2(n_672),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1457),
.B(n_1318),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1427),
.B(n_678),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1569),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1526),
.A2(n_1321),
.B1(n_1325),
.B2(n_1319),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1400),
.Y(n_1765)
);

OA22x2_ASAP7_75t_L g1766 ( 
.A1(n_1652),
.A2(n_1016),
.B1(n_1065),
.B2(n_1064),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1526),
.A2(n_1325),
.B1(n_1326),
.B2(n_1321),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1549),
.A2(n_696),
.B1(n_701),
.B2(n_688),
.Y(n_1768)
);

AO22x2_ASAP7_75t_L g1769 ( 
.A1(n_1560),
.A2(n_696),
.B1(n_701),
.B2(n_688),
.Y(n_1769)
);

NAND3x1_ASAP7_75t_L g1770 ( 
.A(n_1574),
.B(n_1438),
.C(n_1641),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1529),
.A2(n_1548),
.B1(n_1655),
.B2(n_1489),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1561),
.A2(n_716),
.B1(n_718),
.B2(n_703),
.Y(n_1772)
);

AO22x2_ASAP7_75t_L g1773 ( 
.A1(n_1467),
.A2(n_1426),
.B1(n_1534),
.B2(n_1533),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1529),
.A2(n_1328),
.B1(n_1329),
.B2(n_1326),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1459),
.A2(n_716),
.B1(n_718),
.B2(n_703),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1529),
.A2(n_1329),
.B1(n_1330),
.B2(n_1328),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1548),
.A2(n_1489),
.B1(n_1457),
.B2(n_1454),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1416),
.B(n_1067),
.Y(n_1778)
);

AO22x2_ASAP7_75t_L g1779 ( 
.A1(n_1414),
.A2(n_724),
.B1(n_725),
.B2(n_722),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1400),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1548),
.A2(n_1336),
.B1(n_1330),
.B2(n_724),
.Y(n_1781)
);

AO22x2_ASAP7_75t_L g1782 ( 
.A1(n_1414),
.A2(n_725),
.B1(n_726),
.B2(n_722),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1441),
.Y(n_1783)
);

AO22x2_ASAP7_75t_L g1784 ( 
.A1(n_1421),
.A2(n_731),
.B1(n_732),
.B2(n_726),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1457),
.A2(n_1336),
.B1(n_732),
.B2(n_733),
.Y(n_1785)
);

AO22x2_ASAP7_75t_L g1786 ( 
.A1(n_1421),
.A2(n_733),
.B1(n_737),
.B2(n_731),
.Y(n_1786)
);

INVx8_ASAP7_75t_L g1787 ( 
.A(n_1481),
.Y(n_1787)
);

AO22x2_ASAP7_75t_L g1788 ( 
.A1(n_1511),
.A2(n_739),
.B1(n_745),
.B2(n_737),
.Y(n_1788)
);

OAI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1517),
.A2(n_739),
.B1(n_1072),
.B2(n_1067),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1453),
.B(n_1072),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1416),
.B(n_1073),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1441),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1416),
.B(n_1438),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_R g1794 ( 
.A1(n_1558),
.A2(n_1074),
.B1(n_1076),
.B2(n_1073),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1522),
.B(n_1074),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1569),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1455),
.B(n_1477),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1489),
.A2(n_1082),
.B1(n_1083),
.B2(n_1080),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1448),
.B(n_1080),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_SL g1800 ( 
.A1(n_1528),
.A2(n_1085),
.B1(n_1093),
.B2(n_1083),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1441),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1411),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1447),
.B(n_1085),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1411),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1447),
.A2(n_1093),
.B1(n_933),
.B2(n_934),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1447),
.A2(n_933),
.B1(n_934),
.B2(n_931),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1420),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1561),
.Y(n_1808)
);

AO22x2_ASAP7_75t_L g1809 ( 
.A1(n_1511),
.A2(n_943),
.B1(n_941),
.B2(n_936),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1454),
.B(n_931),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1575),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1413),
.B(n_528),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1443),
.B(n_532),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1459),
.A2(n_542),
.B1(n_548),
.B2(n_541),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1407),
.B(n_938),
.Y(n_1815)
);

OAI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1555),
.A2(n_947),
.B1(n_949),
.B2(n_938),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1459),
.A2(n_550),
.B1(n_560),
.B2(n_549),
.Y(n_1817)
);

OA22x2_ASAP7_75t_L g1818 ( 
.A1(n_1540),
.A2(n_949),
.B1(n_954),
.B2(n_947),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1511),
.A2(n_955),
.B1(n_956),
.B2(n_954),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1575),
.A2(n_956),
.B1(n_960),
.B2(n_955),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1566),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1575),
.A2(n_964),
.B1(n_965),
.B2(n_960),
.Y(n_1822)
);

AO22x2_ASAP7_75t_L g1823 ( 
.A1(n_1587),
.A2(n_965),
.B1(n_967),
.B2(n_964),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1612),
.A2(n_969),
.B1(n_971),
.B2(n_967),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1484),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1389),
.A2(n_971),
.B1(n_972),
.B2(n_969),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1612),
.A2(n_973),
.B1(n_980),
.B2(n_972),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1420),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1435),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1612),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1484),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1537),
.A2(n_568),
.B1(n_573),
.B2(n_561),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1495),
.B(n_973),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1495),
.B(n_980),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1417),
.A2(n_983),
.B1(n_986),
.B2(n_982),
.Y(n_1835)
);

AO22x2_ASAP7_75t_L g1836 ( 
.A1(n_1587),
.A2(n_983),
.B1(n_986),
.B2(n_982),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1585),
.B(n_822),
.Y(n_1837)
);

OA22x2_ASAP7_75t_L g1838 ( 
.A1(n_1506),
.A2(n_579),
.B1(n_582),
.B2(n_577),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1485),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1422),
.B(n_593),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1432),
.B(n_822),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1428),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1537),
.Y(n_1843)
);

INVxp33_ASAP7_75t_L g1844 ( 
.A(n_1412),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1603),
.B(n_846),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1603),
.B(n_846),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1435),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1462),
.A2(n_609),
.B1(n_620),
.B2(n_594),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1494),
.B(n_1412),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1442),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1462),
.A2(n_671),
.B1(n_676),
.B2(n_668),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1630),
.A2(n_686),
.B1(n_690),
.B2(n_684),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1542),
.B(n_848),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1470),
.A2(n_714),
.B1(n_721),
.B2(n_706),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1470),
.A2(n_729),
.B1(n_968),
.B2(n_945),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1563),
.B(n_945),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1509),
.A2(n_1001),
.B1(n_968),
.B2(n_1242),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1515),
.A2(n_1001),
.B1(n_1296),
.B2(n_1242),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1524),
.A2(n_1463),
.B1(n_1468),
.B2(n_1418),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1470),
.A2(n_1488),
.B1(n_1499),
.B2(n_1478),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1424),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1543),
.B(n_1567),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1630),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1556),
.A2(n_1320),
.B1(n_1335),
.B2(n_1296),
.Y(n_1864)
);

AO22x2_ASAP7_75t_L g1865 ( 
.A1(n_1587),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_SL g1866 ( 
.A1(n_1388),
.A2(n_1335),
.B1(n_1373),
.B2(n_1320),
.Y(n_1866)
);

AO22x2_ASAP7_75t_L g1867 ( 
.A1(n_1440),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1559),
.A2(n_1373),
.B1(n_12),
.B2(n_9),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1442),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1581),
.B(n_11),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1570),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1871)
);

OR2x6_ASAP7_75t_L g1872 ( 
.A(n_1594),
.B(n_758),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1444),
.Y(n_1873)
);

AO22x2_ASAP7_75t_L g1874 ( 
.A1(n_1581),
.A2(n_17),
.B1(n_13),
.B2(n_16),
.Y(n_1874)
);

AND2x2_ASAP7_75t_SL g1875 ( 
.A(n_1594),
.B(n_17),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1609),
.Y(n_1876)
);

XOR2xp5_ASAP7_75t_L g1877 ( 
.A(n_1609),
.B(n_291),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1543),
.B(n_18),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1642),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_1879)
);

AOI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1550),
.A2(n_742),
.B1(n_790),
.B2(n_758),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1398),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1491),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1491),
.Y(n_1883)
);

OAI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1580),
.A2(n_1646),
.B1(n_1554),
.B2(n_1649),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1444),
.Y(n_1885)
);

OAI22xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1387),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1446),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1588),
.A2(n_742),
.B1(n_790),
.B2(n_758),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1446),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1466),
.Y(n_1890)
);

OAI22xp33_ASAP7_75t_R g1891 ( 
.A1(n_1642),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1567),
.A2(n_742),
.B1(n_790),
.B2(n_758),
.Y(n_1892)
);

OAI22xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1423),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_1893)
);

AO22x2_ASAP7_75t_L g1894 ( 
.A1(n_1434),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1478),
.A2(n_1499),
.B1(n_1504),
.B2(n_1488),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1469),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1478),
.A2(n_790),
.B1(n_843),
.B2(n_758),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1521),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1428),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1644),
.B(n_31),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1488),
.A2(n_843),
.B1(n_870),
.B2(n_790),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1469),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1521),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1472),
.Y(n_1904)
);

INVx5_ASAP7_75t_L g1905 ( 
.A(n_1424),
.Y(n_1905)
);

AO22x2_ASAP7_75t_L g1906 ( 
.A1(n_1439),
.A2(n_1493),
.B1(n_1497),
.B2(n_1496),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1499),
.A2(n_870),
.B1(n_951),
.B2(n_843),
.Y(n_1907)
);

OA22x2_ASAP7_75t_L g1908 ( 
.A1(n_1644),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1908)
);

AO22x2_ASAP7_75t_L g1909 ( 
.A1(n_1512),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1650),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1428),
.Y(n_1911)
);

OAI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1651),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1504),
.A2(n_870),
.B1(n_951),
.B2(n_843),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1431),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1914)
);

AOI22x1_ASAP7_75t_SL g1915 ( 
.A1(n_1599),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1504),
.A2(n_870),
.B1(n_951),
.B2(n_843),
.Y(n_1916)
);

AO22x2_ASAP7_75t_L g1917 ( 
.A1(n_1516),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1917)
);

AOI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1579),
.A2(n_951),
.B1(n_870),
.B2(n_999),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1579),
.A2(n_50),
.B1(n_46),
.B2(n_49),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1428),
.Y(n_1920)
);

BUFx10_ASAP7_75t_L g1921 ( 
.A(n_1424),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1475),
.Y(n_1922)
);

OAI22xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1532),
.A2(n_54),
.B1(n_50),
.B2(n_52),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1586),
.B(n_55),
.Y(n_1924)
);

OAI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1552),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1599),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1686),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1862),
.B(n_1616),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_1668),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1861),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1802),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1861),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1804),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1921),
.Y(n_1934)
);

INVx6_ASAP7_75t_L g1935 ( 
.A(n_1921),
.Y(n_1935)
);

AND2x6_ASAP7_75t_L g1936 ( 
.A(n_1690),
.B(n_1579),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1905),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1663),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1665),
.Y(n_1939)
);

AOI21x1_ASAP7_75t_L g1940 ( 
.A1(n_1688),
.A2(n_1406),
.B(n_1386),
.Y(n_1940)
);

INVxp67_ASAP7_75t_SL g1941 ( 
.A(n_1777),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1665),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1693),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1843),
.B(n_1602),
.Y(n_1944)
);

AND3x1_ASAP7_75t_L g1945 ( 
.A(n_1720),
.B(n_1653),
.C(n_1568),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1884),
.A2(n_1859),
.B(n_1864),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1862),
.B(n_1653),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1685),
.B(n_1404),
.Y(n_1948)
);

NAND2xp33_ASAP7_75t_L g1949 ( 
.A(n_1860),
.B(n_1449),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1807),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1677),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1842),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1771),
.B(n_1404),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1694),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1697),
.Y(n_1955)
);

CKINVDCx6p67_ASAP7_75t_R g1956 ( 
.A(n_1677),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1704),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1787),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1905),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1828),
.Y(n_1960)
);

INVx5_ASAP7_75t_L g1961 ( 
.A(n_1756),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1676),
.B(n_1656),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1899),
.Y(n_1963)
);

AND3x2_ASAP7_75t_L g1964 ( 
.A(n_1698),
.B(n_1617),
.C(n_1572),
.Y(n_1964)
);

NAND2xp33_ASAP7_75t_L g1965 ( 
.A(n_1860),
.B(n_1895),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1687),
.A2(n_1393),
.B1(n_1394),
.B2(n_1385),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1710),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1771),
.B(n_1408),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1799),
.B(n_1803),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1829),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1717),
.B(n_1408),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1847),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1777),
.B(n_1408),
.Y(n_1973)
);

INVx5_ASAP7_75t_L g1974 ( 
.A(n_1740),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1734),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1739),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1690),
.B(n_1419),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1741),
.Y(n_1978)
);

NAND2xp33_ASAP7_75t_L g1979 ( 
.A(n_1895),
.B(n_1449),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1740),
.A2(n_1449),
.B1(n_1451),
.B2(n_1450),
.Y(n_1980)
);

AND2x2_ASAP7_75t_SL g1981 ( 
.A(n_1875),
.B(n_1600),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1763),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1745),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1899),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1661),
.B(n_1419),
.Y(n_1985)
);

INVx4_ASAP7_75t_L g1986 ( 
.A(n_1763),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1748),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1750),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1825),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1831),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1687),
.A2(n_1393),
.B1(n_1394),
.B2(n_1385),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1695),
.B(n_1419),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1911),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1850),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1839),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1869),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1873),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1882),
.Y(n_1998)
);

AND2x6_ASAP7_75t_L g1999 ( 
.A(n_1723),
.B(n_1449),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1833),
.B(n_1834),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1911),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1883),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1926),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1729),
.B(n_1501),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_R g2005 ( 
.A(n_1808),
.B(n_1425),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1898),
.Y(n_2006)
);

AND2x6_ASAP7_75t_L g2007 ( 
.A(n_1723),
.B(n_1449),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1680),
.B(n_1656),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1673),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1903),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1906),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1920),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1906),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1798),
.B(n_1501),
.Y(n_2014)
);

OAI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1796),
.A2(n_1450),
.B1(n_1452),
.B2(n_1451),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1885),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1920),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1796),
.B(n_1386),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1787),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1887),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1811),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_1703),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1671),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1889),
.Y(n_2024)
);

INVx4_ASAP7_75t_SL g2025 ( 
.A(n_1673),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1718),
.B(n_1424),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1811),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1890),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1682),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1684),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1736),
.B(n_1656),
.Y(n_2031)
);

INVxp33_ASAP7_75t_SL g2032 ( 
.A(n_1679),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1863),
.B(n_1691),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1705),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1684),
.Y(n_2035)
);

INVxp33_ASAP7_75t_SL g2036 ( 
.A(n_1708),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1707),
.A2(n_1409),
.B1(n_1410),
.B2(n_1406),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1670),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1712),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1896),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1902),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1778),
.B(n_1791),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1830),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1719),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1672),
.B(n_1656),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1681),
.B(n_1621),
.Y(n_2046)
);

INVxp33_ASAP7_75t_L g2047 ( 
.A(n_1669),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1670),
.B(n_1450),
.Y(n_2048)
);

INVx5_ASAP7_75t_L g2049 ( 
.A(n_1662),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1904),
.Y(n_2050)
);

AND2x6_ASAP7_75t_L g2051 ( 
.A(n_1701),
.B(n_1450),
.Y(n_2051)
);

INVx4_ASAP7_75t_L g2052 ( 
.A(n_1662),
.Y(n_2052)
);

INVx1_ASAP7_75t_SL g2053 ( 
.A(n_1692),
.Y(n_2053)
);

BUFx2_ASAP7_75t_L g2054 ( 
.A(n_1849),
.Y(n_2054)
);

NOR2x1p5_ASAP7_75t_L g2055 ( 
.A(n_1711),
.B(n_1643),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1922),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1681),
.B(n_1479),
.Y(n_2057)
);

AND2x2_ASAP7_75t_SL g2058 ( 
.A(n_1733),
.B(n_1600),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1689),
.B(n_1486),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1810),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1742),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1793),
.A2(n_1451),
.B1(n_1452),
.B2(n_1450),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1674),
.B(n_1667),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1696),
.B(n_1486),
.Y(n_2064)
);

BUFx10_ASAP7_75t_L g2065 ( 
.A(n_1702),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1841),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1666),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1678),
.B(n_1451),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1696),
.B(n_1490),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1765),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1764),
.A2(n_1452),
.B1(n_1464),
.B2(n_1451),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1761),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1853),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1701),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_L g2075 ( 
.A(n_1714),
.B(n_1715),
.C(n_1848),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1780),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1783),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1792),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1707),
.A2(n_1410),
.B1(n_1409),
.B2(n_1647),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1728),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1844),
.B(n_1452),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1801),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1853),
.Y(n_2083)
);

AND2x2_ASAP7_75t_SL g2084 ( 
.A(n_1721),
.B(n_1615),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1876),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1837),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_1872),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1749),
.B(n_1452),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_1744),
.A2(n_1773),
.B1(n_1683),
.B2(n_1794),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1770),
.B(n_1492),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1878),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1821),
.B(n_1706),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1709),
.B(n_1722),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_1747),
.B(n_1492),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1924),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1744),
.A2(n_1658),
.B1(n_1647),
.B2(n_1508),
.Y(n_2096)
);

INVx6_ASAP7_75t_L g2097 ( 
.A(n_1872),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1820),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1845),
.B(n_1498),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1897),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1846),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1820),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1743),
.B(n_1508),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1743),
.B(n_1510),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1737),
.A2(n_1465),
.B1(n_1482),
.B2(n_1464),
.Y(n_2105)
);

CKINVDCx6p67_ASAP7_75t_R g2106 ( 
.A(n_1762),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1897),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1713),
.B(n_1464),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1805),
.B(n_1510),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1901),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1738),
.B(n_1465),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1901),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1822),
.Y(n_2113)
);

OAI21xp33_ASAP7_75t_SL g2114 ( 
.A1(n_1721),
.A2(n_1619),
.B(n_1547),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1907),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1856),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1731),
.B(n_1513),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1764),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1767),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1746),
.B(n_1465),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1805),
.B(n_1465),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1907),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1767),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1774),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1806),
.B(n_1615),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1754),
.B(n_1465),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1913),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1913),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1916),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_1795),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1774),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1724),
.B(n_1482),
.Y(n_2132)
);

INVxp67_ASAP7_75t_SL g2133 ( 
.A(n_1724),
.Y(n_2133)
);

BUFx10_ASAP7_75t_L g2134 ( 
.A(n_1812),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1797),
.Y(n_2135)
);

INVx11_ASAP7_75t_L g2136 ( 
.A(n_1877),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1776),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1776),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1755),
.Y(n_2139)
);

AND2x6_ASAP7_75t_L g2140 ( 
.A(n_1725),
.B(n_1482),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1806),
.B(n_1513),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1755),
.B(n_1781),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1916),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1918),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1785),
.B(n_1518),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1918),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1785),
.B(n_1518),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1824),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_L g2149 ( 
.A(n_1813),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1892),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1725),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_1781),
.B(n_1527),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1779),
.B(n_1615),
.Y(n_2153)
);

BUFx3_ASAP7_75t_L g2154 ( 
.A(n_1735),
.Y(n_2154)
);

AOI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_1840),
.A2(n_1487),
.B1(n_1541),
.B2(n_1482),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1726),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1726),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_SL g2158 ( 
.A1(n_1773),
.A2(n_1531),
.B1(n_1539),
.B2(n_1527),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1727),
.B(n_1730),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1751),
.A2(n_1487),
.B1(n_1541),
.B2(n_1482),
.Y(n_2160)
);

BUFx10_ASAP7_75t_L g2161 ( 
.A(n_1832),
.Y(n_2161)
);

AO22x2_ASAP7_75t_L g2162 ( 
.A1(n_1915),
.A2(n_1658),
.B1(n_1539),
.B2(n_1571),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1727),
.Y(n_2163)
);

OR2x6_ASAP7_75t_L g2164 ( 
.A(n_1819),
.B(n_1531),
.Y(n_2164)
);

INVx4_ASAP7_75t_L g2165 ( 
.A(n_1819),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_1790),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1730),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1824),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_SL g2169 ( 
.A1(n_1788),
.A2(n_1590),
.B1(n_1597),
.B2(n_1577),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_1815),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1827),
.B(n_1577),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1732),
.B(n_1487),
.Y(n_2172)
);

NAND2xp33_ASAP7_75t_L g2173 ( 
.A(n_1732),
.B(n_1487),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1766),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1775),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1779),
.B(n_1782),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1816),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1880),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1660),
.B(n_1541),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1826),
.Y(n_2180)
);

INVxp33_ASAP7_75t_L g2181 ( 
.A(n_1852),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1870),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_1900),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1866),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1888),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1835),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1855),
.Y(n_2187)
);

INVx4_ASAP7_75t_L g2188 ( 
.A(n_1935),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_1929),
.Y(n_2189)
);

AO22x2_ASAP7_75t_L g2190 ( 
.A1(n_2165),
.A2(n_1788),
.B1(n_1758),
.B2(n_1823),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1951),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1937),
.Y(n_2192)
);

AND2x6_ASAP7_75t_L g2193 ( 
.A(n_2142),
.B(n_1753),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1947),
.B(n_1753),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1927),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1943),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2118),
.B(n_1597),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2170),
.B(n_1757),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2142),
.A2(n_1891),
.B1(n_1757),
.B2(n_1865),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1957),
.Y(n_2200)
);

INVxp33_ASAP7_75t_L g2201 ( 
.A(n_2092),
.Y(n_2201)
);

AND2x4_ASAP7_75t_SL g2202 ( 
.A(n_1956),
.B(n_1605),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1937),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2118),
.B(n_1605),
.Y(n_2204)
);

INVx2_ASAP7_75t_SL g2205 ( 
.A(n_1951),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_1947),
.B(n_1610),
.Y(n_2206)
);

BUFx4f_ASAP7_75t_L g2207 ( 
.A(n_1956),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1931),
.Y(n_2208)
);

INVxp67_ASAP7_75t_L g2209 ( 
.A(n_2170),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1967),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1937),
.Y(n_2211)
);

AOI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_2142),
.A2(n_1782),
.B1(n_1786),
.B2(n_1784),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_2003),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1931),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1995),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1994),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_1947),
.B(n_1610),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1994),
.Y(n_2218)
);

BUFx4f_ASAP7_75t_L g2219 ( 
.A(n_2106),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2025),
.B(n_1614),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2119),
.B(n_1614),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1933),
.Y(n_2222)
);

INVx4_ASAP7_75t_SL g2223 ( 
.A(n_1999),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2166),
.B(n_1769),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1996),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1998),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2119),
.B(n_2138),
.Y(n_2227)
);

INVx6_ASAP7_75t_L g2228 ( 
.A(n_2025),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1996),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2002),
.Y(n_2230)
);

INVx5_ASAP7_75t_L g2231 ( 
.A(n_1999),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_1935),
.Y(n_2232)
);

INVx4_ASAP7_75t_L g2233 ( 
.A(n_1935),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2006),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2010),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1937),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_2003),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2042),
.B(n_1769),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2042),
.B(n_1784),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1954),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1954),
.Y(n_2241)
);

BUFx4f_ASAP7_75t_L g2242 ( 
.A(n_2106),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1933),
.Y(n_2243)
);

BUFx2_ASAP7_75t_L g2244 ( 
.A(n_2085),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1955),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1950),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1950),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_1944),
.Y(n_2248)
);

AND2x6_ASAP7_75t_L g2249 ( 
.A(n_2123),
.B(n_1573),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1975),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_1937),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_2054),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2058),
.B(n_1573),
.Y(n_2253)
);

AND2x2_ASAP7_75t_SL g2254 ( 
.A(n_2058),
.B(n_1865),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1975),
.Y(n_2255)
);

AND2x6_ASAP7_75t_L g2256 ( 
.A(n_2123),
.B(n_1573),
.Y(n_2256)
);

INVxp67_ASAP7_75t_L g2257 ( 
.A(n_2054),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1976),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1934),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1997),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1976),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1997),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1978),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1978),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1983),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2016),
.Y(n_2266)
);

OR2x2_ASAP7_75t_SL g2267 ( 
.A(n_2075),
.B(n_1675),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1983),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1987),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1987),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2124),
.B(n_1623),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2036),
.B(n_1789),
.Y(n_2272)
);

OAI221xp5_ASAP7_75t_L g2273 ( 
.A1(n_2089),
.A2(n_1879),
.B1(n_1908),
.B2(n_1919),
.C(n_1759),
.Y(n_2273)
);

CKINVDCx14_ASAP7_75t_R g2274 ( 
.A(n_2022),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2025),
.B(n_1623),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2016),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2020),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2131),
.B(n_1576),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1988),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_2047),
.B(n_1800),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1989),
.Y(n_2281)
);

BUFx3_ASAP7_75t_L g2282 ( 
.A(n_1958),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1989),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2025),
.B(n_1627),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2137),
.B(n_1627),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1990),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1928),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1928),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1960),
.Y(n_2289)
);

NAND2x1p5_ASAP7_75t_L g2290 ( 
.A(n_1974),
.B(n_1615),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1934),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2011),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2047),
.B(n_1786),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2063),
.A2(n_1874),
.B1(n_1851),
.B2(n_1854),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_2038),
.B(n_1629),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2053),
.B(n_1752),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_1982),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2137),
.B(n_1629),
.Y(n_2298)
);

NAND2x1p5_ASAP7_75t_L g2299 ( 
.A(n_1974),
.B(n_1657),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2013),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2024),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_1981),
.A2(n_1874),
.B1(n_1854),
.B2(n_1818),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2176),
.B(n_1809),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2138),
.B(n_1634),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_1982),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2086),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2176),
.A2(n_1981),
.B1(n_2164),
.B2(n_2165),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_2038),
.B(n_1634),
.Y(n_2308)
);

AND2x6_ASAP7_75t_L g2309 ( 
.A(n_2139),
.B(n_1576),
.Y(n_2309)
);

BUFx2_ASAP7_75t_L g2310 ( 
.A(n_2085),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2024),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1982),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1941),
.B(n_1969),
.Y(n_2313)
);

AO22x2_ASAP7_75t_L g2314 ( 
.A1(n_2165),
.A2(n_1836),
.B1(n_1823),
.B2(n_1809),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2117),
.B(n_2019),
.Y(n_2315)
);

INVx4_ASAP7_75t_SL g2316 ( 
.A(n_1999),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2028),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2040),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_1945),
.A2(n_1760),
.B1(n_1772),
.B2(n_1768),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_1986),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2117),
.B(n_1657),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2041),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_1938),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2040),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2060),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2093),
.B(n_1836),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_1948),
.B(n_1699),
.Y(n_2327)
);

NAND3x1_ASAP7_75t_L g2328 ( 
.A(n_2032),
.B(n_1867),
.C(n_1675),
.Y(n_2328)
);

AO22x2_ASAP7_75t_L g2329 ( 
.A1(n_2139),
.A2(n_1664),
.B1(n_1917),
.B2(n_1909),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_1934),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2094),
.Y(n_2331)
);

NAND2x1p5_ASAP7_75t_L g2332 ( 
.A(n_1974),
.B(n_1425),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2000),
.B(n_1535),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_1934),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_1934),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_1986),
.Y(n_2336)
);

AND2x6_ASAP7_75t_L g2337 ( 
.A(n_2151),
.B(n_1576),
.Y(n_2337)
);

AO22x2_ASAP7_75t_L g2338 ( 
.A1(n_2159),
.A2(n_1664),
.B1(n_1917),
.B2(n_1909),
.Y(n_2338)
);

BUFx3_ASAP7_75t_L g2339 ( 
.A(n_2035),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_L g2340 ( 
.A(n_2088),
.B(n_1817),
.C(n_1814),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2072),
.B(n_1535),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2117),
.B(n_1547),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1970),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_1939),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2027),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1972),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_1935),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2067),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1972),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2155),
.B(n_1578),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2093),
.B(n_1700),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2093),
.B(n_1716),
.Y(n_2352)
);

INVx8_ASAP7_75t_L g2353 ( 
.A(n_1974),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2009),
.Y(n_2354)
);

CKINVDCx16_ASAP7_75t_R g2355 ( 
.A(n_2022),
.Y(n_2355)
);

NAND2x1p5_ASAP7_75t_L g2356 ( 
.A(n_1974),
.B(n_1425),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2039),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_1942),
.B(n_1582),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2027),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2135),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_R g2361 ( 
.A(n_2061),
.B(n_1578),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2130),
.B(n_1894),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2050),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_1942),
.B(n_1582),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2050),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2130),
.B(n_1894),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2009),
.B(n_2030),
.Y(n_2367)
);

BUFx3_ASAP7_75t_L g2368 ( 
.A(n_2097),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2056),
.Y(n_2369)
);

AND2x6_ASAP7_75t_L g2370 ( 
.A(n_2151),
.B(n_1578),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2126),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2066),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2055),
.B(n_1838),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_2097),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2074),
.A2(n_1925),
.B1(n_1886),
.B2(n_1871),
.Y(n_2375)
);

INVx4_ASAP7_75t_L g2376 ( 
.A(n_2097),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2174),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2181),
.B(n_1855),
.Y(n_2378)
);

BUFx4_ASAP7_75t_L g2379 ( 
.A(n_2032),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2070),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2027),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2076),
.Y(n_2382)
);

OR2x2_ASAP7_75t_SL g2383 ( 
.A(n_1944),
.B(n_1893),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2098),
.B(n_1583),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2102),
.B(n_1583),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2033),
.B(n_2101),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_SL g2387 ( 
.A1(n_2254),
.A2(n_2162),
.B1(n_2133),
.B2(n_2061),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2248),
.B(n_2154),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2361),
.B(n_2134),
.Y(n_2389)
);

INVx2_ASAP7_75t_SL g2390 ( 
.A(n_2207),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2252),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2313),
.B(n_2026),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2294),
.B(n_2134),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2198),
.B(n_2181),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2331),
.B(n_2175),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2252),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_SL g2397 ( 
.A(n_2191),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2201),
.B(n_2101),
.Y(n_2398)
);

AOI22xp33_ASAP7_75t_SL g2399 ( 
.A1(n_2254),
.A2(n_2162),
.B1(n_2164),
.B2(n_2140),
.Y(n_2399)
);

BUFx8_ASAP7_75t_SL g2400 ( 
.A(n_2379),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2195),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2227),
.B(n_2113),
.Y(n_2402)
);

AOI221xp5_ASAP7_75t_SL g2403 ( 
.A1(n_2327),
.A2(n_1910),
.B1(n_1912),
.B2(n_2273),
.C(n_1868),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2386),
.B(n_2148),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2386),
.B(n_2168),
.Y(n_2405)
);

BUFx8_ASAP7_75t_L g2406 ( 
.A(n_2244),
.Y(n_2406)
);

AOI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2319),
.A2(n_2161),
.B1(n_2162),
.B2(n_2183),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2353),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2207),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2201),
.B(n_2101),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_2371),
.B(n_1971),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2212),
.B(n_2081),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2371),
.B(n_1992),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2327),
.B(n_2004),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2196),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2212),
.B(n_2045),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2272),
.B(n_2378),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2200),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2272),
.B(n_2116),
.Y(n_2419)
);

INVxp67_ASAP7_75t_L g2420 ( 
.A(n_2237),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2209),
.B(n_2045),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2210),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2293),
.B(n_2154),
.Y(n_2423)
);

AND3x1_ASAP7_75t_L g2424 ( 
.A(n_2199),
.B(n_2179),
.C(n_2161),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2194),
.B(n_2116),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2228),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2194),
.B(n_2116),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2238),
.B(n_2182),
.Y(n_2428)
);

A2O1A1Ixp33_ASAP7_75t_SL g2429 ( 
.A1(n_2351),
.A2(n_2095),
.B(n_2091),
.C(n_1963),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2239),
.B(n_2095),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2257),
.B(n_2158),
.Y(n_2431)
);

AOI22xp33_ASAP7_75t_L g2432 ( 
.A1(n_2193),
.A2(n_2338),
.B1(n_2190),
.B2(n_2329),
.Y(n_2432)
);

BUFx2_ASAP7_75t_L g2433 ( 
.A(n_2310),
.Y(n_2433)
);

INVx2_ASAP7_75t_SL g2434 ( 
.A(n_2219),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2215),
.Y(n_2435)
);

AOI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2193),
.A2(n_2161),
.B1(n_2162),
.B2(n_1936),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2216),
.Y(n_2437)
);

NAND2xp33_ASAP7_75t_L g2438 ( 
.A(n_2193),
.B(n_1936),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2333),
.B(n_1966),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2226),
.Y(n_2440)
);

O2A1O1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_2273),
.A2(n_1985),
.B(n_1965),
.C(n_2048),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_2237),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2193),
.A2(n_1936),
.B1(n_2152),
.B2(n_2007),
.Y(n_2443)
);

NAND2xp33_ASAP7_75t_L g2444 ( 
.A(n_2193),
.B(n_1936),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2231),
.B(n_2014),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2333),
.B(n_1991),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2189),
.B(n_1964),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2361),
.B(n_2049),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2218),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2189),
.B(n_2152),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2342),
.B(n_2049),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2302),
.B(n_1986),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2368),
.B(n_2090),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2338),
.A2(n_2164),
.B1(n_2090),
.B2(n_2169),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2342),
.B(n_2152),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2225),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2229),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_SL g2458 ( 
.A(n_2357),
.B(n_2087),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2287),
.B(n_2182),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2224),
.B(n_2031),
.Y(n_2460)
);

INVxp67_ASAP7_75t_SL g2461 ( 
.A(n_2197),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2288),
.B(n_2031),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2296),
.B(n_1973),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2338),
.A2(n_1936),
.B1(n_2007),
.B2(n_1999),
.Y(n_2464)
);

BUFx8_ASAP7_75t_L g2465 ( 
.A(n_2213),
.Y(n_2465)
);

AOI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2296),
.A2(n_1936),
.B1(n_2007),
.B2(n_1999),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2321),
.B(n_1953),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2231),
.B(n_2071),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2190),
.A2(n_2164),
.B1(n_2090),
.B2(n_2187),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2231),
.B(n_2099),
.Y(n_2470)
);

OAI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_2340),
.A2(n_2120),
.B(n_2111),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2323),
.B(n_2099),
.Y(n_2472)
);

BUFx2_ASAP7_75t_L g2473 ( 
.A(n_2315),
.Y(n_2473)
);

INVx8_ASAP7_75t_L g2474 ( 
.A(n_2353),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2231),
.B(n_2099),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2190),
.A2(n_2090),
.B1(n_2187),
.B2(n_2157),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2323),
.B(n_2018),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2375),
.A2(n_2046),
.B1(n_2157),
.B2(n_2156),
.Y(n_2478)
);

OR2x2_ASAP7_75t_L g2479 ( 
.A(n_2344),
.B(n_2073),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2230),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2326),
.B(n_2153),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2206),
.B(n_2018),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_2384),
.B(n_2105),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2234),
.Y(n_2484)
);

AOI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_2280),
.A2(n_1999),
.B1(n_2007),
.B2(n_1965),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2280),
.A2(n_2007),
.B1(n_2005),
.B2(n_2051),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2217),
.B(n_2018),
.Y(n_2487)
);

NOR2x2_ASAP7_75t_L g2488 ( 
.A(n_2274),
.B(n_2136),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2329),
.A2(n_2007),
.B1(n_2140),
.B2(n_2051),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2321),
.B(n_2083),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2235),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2329),
.A2(n_2051),
.B1(n_2140),
.B2(n_1968),
.Y(n_2492)
);

BUFx3_ASAP7_75t_L g2493 ( 
.A(n_2191),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2352),
.A2(n_2051),
.B1(n_2140),
.B2(n_2097),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2282),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2306),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2240),
.B(n_1962),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2260),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2242),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2325),
.Y(n_2500)
);

AOI22xp33_ASAP7_75t_L g2501 ( 
.A1(n_2314),
.A2(n_2163),
.B1(n_2167),
.B2(n_2156),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2368),
.B(n_2087),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2262),
.Y(n_2503)
);

AND2x4_ASAP7_75t_L g2504 ( 
.A(n_2374),
.B(n_2087),
.Y(n_2504)
);

NAND4xp25_ASAP7_75t_SL g2505 ( 
.A(n_2307),
.B(n_1923),
.C(n_1914),
.D(n_1881),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_L g2506 ( 
.A(n_2253),
.B(n_2027),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2314),
.A2(n_2303),
.B1(n_2167),
.B2(n_2163),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2266),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2276),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2241),
.B(n_2008),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2384),
.B(n_2108),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2374),
.B(n_2376),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2277),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2245),
.B(n_2008),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2353),
.Y(n_2515)
);

HB1xp67_ASAP7_75t_L g2516 ( 
.A(n_2253),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2314),
.A2(n_2147),
.B1(n_2145),
.B2(n_2051),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2250),
.B(n_2255),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2258),
.B(n_2261),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2360),
.B(n_2064),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2301),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2348),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2383),
.B(n_2043),
.Y(n_2523)
);

INVx8_ASAP7_75t_L g2524 ( 
.A(n_2220),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2351),
.A2(n_2364),
.B1(n_2358),
.B2(n_2373),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2263),
.B(n_2264),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2265),
.B(n_2043),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2376),
.B(n_2043),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2268),
.B(n_2043),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2269),
.B(n_2069),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2242),
.B(n_2049),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2311),
.Y(n_2532)
);

AO22x1_ASAP7_75t_L g2533 ( 
.A1(n_2220),
.A2(n_2140),
.B1(n_2051),
.B2(n_2149),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2228),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2372),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2317),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2341),
.B(n_1977),
.Y(n_2537)
);

BUFx8_ASAP7_75t_L g2538 ( 
.A(n_2205),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2270),
.B(n_2057),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2279),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2362),
.A2(n_2140),
.B1(n_2186),
.B2(n_2180),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2366),
.B(n_2021),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2322),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2281),
.B(n_2059),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2188),
.B(n_2049),
.Y(n_2545)
);

INVx5_ASAP7_75t_L g2546 ( 
.A(n_2228),
.Y(n_2546)
);

A2O1A1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2385),
.A2(n_2068),
.B(n_2173),
.C(n_2062),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2363),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2355),
.B(n_2065),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2401),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2546),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2417),
.B(n_2292),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2424),
.A2(n_2328),
.B1(n_2364),
.B2(n_2358),
.Y(n_2553)
);

INVxp33_ASAP7_75t_L g2554 ( 
.A(n_2388),
.Y(n_2554)
);

NAND3xp33_ASAP7_75t_SL g2555 ( 
.A(n_2407),
.B(n_2385),
.C(n_2341),
.Y(n_2555)
);

BUFx4f_ASAP7_75t_L g2556 ( 
.A(n_2426),
.Y(n_2556)
);

BUFx4f_ASAP7_75t_L g2557 ( 
.A(n_2426),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2415),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2437),
.Y(n_2559)
);

CKINVDCx14_ASAP7_75t_R g2560 ( 
.A(n_2549),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2418),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2422),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2394),
.B(n_2339),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2449),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2538),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2436),
.A2(n_2275),
.B1(n_2284),
.B2(n_2274),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_2392),
.B(n_2223),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2435),
.Y(n_2568)
);

INVx2_ASAP7_75t_SL g2569 ( 
.A(n_2538),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2440),
.Y(n_2570)
);

AND2x6_ASAP7_75t_L g2571 ( 
.A(n_2443),
.B(n_2223),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2463),
.B(n_2283),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_2465),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_2417),
.A2(n_2307),
.B1(n_1946),
.B2(n_2377),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2546),
.B(n_2223),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2463),
.A2(n_2284),
.B1(n_2275),
.B2(n_2249),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2548),
.Y(n_2577)
);

BUFx3_ASAP7_75t_L g2578 ( 
.A(n_2493),
.Y(n_2578)
);

INVxp67_ASAP7_75t_SL g2579 ( 
.A(n_2461),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2546),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2414),
.B(n_2316),
.Y(n_2581)
);

BUFx3_ASAP7_75t_L g2582 ( 
.A(n_2495),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2480),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2484),
.Y(n_2584)
);

AND2x6_ASAP7_75t_SL g2585 ( 
.A(n_2400),
.B(n_2367),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2393),
.B(n_2188),
.Y(n_2586)
);

BUFx2_ASAP7_75t_L g2587 ( 
.A(n_2465),
.Y(n_2587)
);

INVx1_ASAP7_75t_SL g2588 ( 
.A(n_2433),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2491),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2428),
.B(n_2339),
.Y(n_2590)
);

INVx5_ASAP7_75t_L g2591 ( 
.A(n_2546),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2522),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2496),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2474),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2406),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2474),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2516),
.Y(n_2597)
);

INVx5_ASAP7_75t_L g2598 ( 
.A(n_2474),
.Y(n_2598)
);

BUFx4f_ASAP7_75t_L g2599 ( 
.A(n_2426),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2402),
.B(n_2404),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2500),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2405),
.B(n_2286),
.Y(n_2602)
);

INVx3_ASAP7_75t_L g2603 ( 
.A(n_2426),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2524),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2535),
.Y(n_2605)
);

HB1xp67_ASAP7_75t_L g2606 ( 
.A(n_2396),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2540),
.Y(n_2607)
);

INVx5_ASAP7_75t_L g2608 ( 
.A(n_2534),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2387),
.A2(n_1946),
.B1(n_2186),
.B2(n_2295),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_SL g2610 ( 
.A1(n_2419),
.A2(n_2267),
.B1(n_2249),
.B2(n_2256),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2518),
.Y(n_2611)
);

OAI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_2466),
.A2(n_2104),
.B1(n_2103),
.B2(n_2109),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2519),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2534),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2456),
.Y(n_2615)
);

INVx5_ASAP7_75t_L g2616 ( 
.A(n_2534),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2526),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2457),
.Y(n_2618)
);

INVxp67_ASAP7_75t_SL g2619 ( 
.A(n_2461),
.Y(n_2619)
);

INVxp67_ASAP7_75t_L g2620 ( 
.A(n_2419),
.Y(n_2620)
);

BUFx12f_ASAP7_75t_L g2621 ( 
.A(n_2406),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2498),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_2397),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2503),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2508),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2509),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2513),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2393),
.B(n_2232),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2521),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2387),
.A2(n_1946),
.B1(n_2308),
.B2(n_2295),
.Y(n_2630)
);

INVx2_ASAP7_75t_SL g2631 ( 
.A(n_2524),
.Y(n_2631)
);

INVxp67_ASAP7_75t_SL g2632 ( 
.A(n_2438),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_L g2633 ( 
.A(n_2482),
.B(n_2232),
.Y(n_2633)
);

HB1xp67_ASAP7_75t_L g2634 ( 
.A(n_2420),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2532),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2537),
.B(n_2316),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2453),
.B(n_2316),
.Y(n_2637)
);

INVx2_ASAP7_75t_SL g2638 ( 
.A(n_2524),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2536),
.Y(n_2639)
);

AND2x6_ASAP7_75t_L g2640 ( 
.A(n_2489),
.B(n_2345),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2543),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_2397),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2450),
.Y(n_2643)
);

OR2x2_ASAP7_75t_L g2644 ( 
.A(n_2391),
.B(n_2300),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2481),
.B(n_2354),
.Y(n_2645)
);

AOI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_2452),
.A2(n_2256),
.B1(n_2309),
.B2(n_2249),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2527),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2395),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2542),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2529),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2528),
.Y(n_2651)
);

NOR2x1p5_ASAP7_75t_L g2652 ( 
.A(n_2447),
.B(n_2233),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2537),
.B(n_2197),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2453),
.B(n_2233),
.Y(n_2654)
);

NAND3xp33_ASAP7_75t_SL g2655 ( 
.A(n_2458),
.B(n_2096),
.C(n_2347),
.Y(n_2655)
);

NAND2x1p5_ASAP7_75t_L g2656 ( 
.A(n_2448),
.B(n_2345),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2485),
.B(n_2204),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2390),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2539),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2409),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2520),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_R g2662 ( 
.A(n_2444),
.B(n_2347),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2430),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2487),
.B(n_2308),
.Y(n_2664)
);

INVx5_ASAP7_75t_L g2665 ( 
.A(n_2408),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2544),
.Y(n_2666)
);

CKINVDCx6p67_ASAP7_75t_R g2667 ( 
.A(n_2389),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2512),
.Y(n_2668)
);

CKINVDCx16_ASAP7_75t_R g2669 ( 
.A(n_2434),
.Y(n_2669)
);

CKINVDCx20_ASAP7_75t_R g2670 ( 
.A(n_2473),
.Y(n_2670)
);

AND2x6_ASAP7_75t_L g2671 ( 
.A(n_2464),
.B(n_2345),
.Y(n_2671)
);

OR2x6_ASAP7_75t_L g2672 ( 
.A(n_2533),
.B(n_2204),
.Y(n_2672)
);

INVx1_ASAP7_75t_SL g2673 ( 
.A(n_2488),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2420),
.Y(n_2674)
);

BUFx6f_ASAP7_75t_L g2675 ( 
.A(n_2512),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2528),
.Y(n_2676)
);

BUFx2_ASAP7_75t_L g2677 ( 
.A(n_2442),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2442),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2502),
.B(n_2259),
.Y(n_2679)
);

INVx2_ASAP7_75t_SL g2680 ( 
.A(n_2479),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2399),
.A2(n_2084),
.B1(n_2324),
.B2(n_2318),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2502),
.Y(n_2682)
);

CKINVDCx6p67_ASAP7_75t_R g2683 ( 
.A(n_2459),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2411),
.B(n_2221),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2530),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2472),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2504),
.B(n_2259),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2423),
.Y(n_2688)
);

INVx3_ASAP7_75t_L g2689 ( 
.A(n_2408),
.Y(n_2689)
);

AOI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_2452),
.A2(n_2256),
.B1(n_2309),
.B2(n_2249),
.Y(n_2690)
);

NOR3xp33_ASAP7_75t_L g2691 ( 
.A(n_2403),
.B(n_2505),
.C(n_2441),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2504),
.B(n_2259),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2511),
.Y(n_2693)
);

INVx2_ASAP7_75t_SL g2694 ( 
.A(n_2499),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2511),
.Y(n_2695)
);

BUFx12f_ASAP7_75t_SL g2696 ( 
.A(n_2398),
.Y(n_2696)
);

BUFx3_ASAP7_75t_L g2697 ( 
.A(n_2490),
.Y(n_2697)
);

BUFx4f_ASAP7_75t_L g2698 ( 
.A(n_2515),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2477),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2497),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2460),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2510),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_2399),
.A2(n_2084),
.B1(n_2177),
.B2(n_2249),
.Y(n_2703)
);

AOI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2579),
.A2(n_1979),
.B(n_1949),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2579),
.A2(n_1979),
.B(n_1949),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2600),
.B(n_2421),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2618),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2619),
.A2(n_2468),
.B(n_2547),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2668),
.Y(n_2709)
);

O2A1O1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2691),
.A2(n_2429),
.B(n_2413),
.C(n_2478),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2619),
.A2(n_2468),
.B(n_2483),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2622),
.Y(n_2712)
);

OR2x6_ASAP7_75t_SL g2713 ( 
.A(n_2595),
.B(n_2431),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2634),
.Y(n_2714)
);

AOI22x1_ASAP7_75t_L g2715 ( 
.A1(n_2674),
.A2(n_2669),
.B1(n_2678),
.B2(n_2677),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2588),
.B(n_2410),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2560),
.B(n_2523),
.Y(n_2717)
);

O2A1O1Ixp33_ASAP7_75t_SL g2718 ( 
.A1(n_2673),
.A2(n_2429),
.B(n_2531),
.C(n_2523),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2572),
.B(n_2439),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2586),
.B(n_2525),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2626),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2648),
.B(n_2446),
.Y(n_2722)
);

OA22x2_ASAP7_75t_L g2723 ( 
.A1(n_2553),
.A2(n_2486),
.B1(n_2494),
.B2(n_2492),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2691),
.A2(n_2690),
.B1(n_2646),
.B2(n_2703),
.Y(n_2724)
);

AO21x1_ASAP7_75t_L g2725 ( 
.A1(n_2602),
.A2(n_2684),
.B(n_2653),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2703),
.A2(n_2432),
.B1(n_2454),
.B2(n_2541),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2632),
.A2(n_2483),
.B(n_2445),
.Y(n_2727)
);

O2A1O1Ixp5_ASAP7_75t_L g2728 ( 
.A1(n_2657),
.A2(n_2471),
.B(n_2445),
.C(n_2278),
.Y(n_2728)
);

OAI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2620),
.A2(n_2432),
.B1(n_2454),
.B2(n_2541),
.Y(n_2729)
);

OAI21x1_ASAP7_75t_L g2730 ( 
.A1(n_2657),
.A2(n_1940),
.B(n_2567),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_SL g2731 ( 
.A(n_2604),
.B(n_2621),
.Y(n_2731)
);

OAI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2555),
.A2(n_2467),
.B(n_2506),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2551),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2668),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2699),
.B(n_2611),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2613),
.B(n_2617),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2586),
.B(n_2628),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2639),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2569),
.B(n_2578),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2680),
.B(n_2412),
.Y(n_2740)
);

OAI21xp33_ASAP7_75t_L g2741 ( 
.A1(n_2620),
.A2(n_2517),
.B(n_2506),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2641),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2609),
.A2(n_2469),
.B1(n_2517),
.B2(n_2476),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2563),
.B(n_2425),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2649),
.B(n_2501),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_L g2746 ( 
.A(n_2578),
.B(n_2291),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2645),
.B(n_2425),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2606),
.Y(n_2748)
);

OAI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2655),
.A2(n_2467),
.B(n_2309),
.Y(n_2749)
);

AOI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2612),
.A2(n_2672),
.B(n_2114),
.Y(n_2750)
);

O2A1O1Ixp5_ASAP7_75t_L g2751 ( 
.A1(n_2581),
.A2(n_2451),
.B(n_2545),
.C(n_2350),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2582),
.B(n_2291),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2623),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2672),
.A2(n_2015),
.B(n_1980),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2582),
.B(n_2330),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2672),
.A2(n_2514),
.B(n_2285),
.Y(n_2756)
);

AOI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2636),
.A2(n_2285),
.B(n_2271),
.Y(n_2757)
);

AOI22xp33_ASAP7_75t_L g2758 ( 
.A1(n_2609),
.A2(n_2469),
.B1(n_2476),
.B2(n_2416),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2681),
.A2(n_2427),
.B1(n_2507),
.B2(n_2455),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2701),
.B(n_2462),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2607),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_2642),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2636),
.A2(n_2298),
.B(n_2271),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2643),
.B(n_2686),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2551),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2567),
.A2(n_2172),
.B(n_2132),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2661),
.B(n_2507),
.Y(n_2767)
);

A2O1A1Ixp33_ASAP7_75t_L g2768 ( 
.A1(n_2610),
.A2(n_2202),
.B(n_2149),
.C(n_2304),
.Y(n_2768)
);

INVxp67_ASAP7_75t_L g2769 ( 
.A(n_2590),
.Y(n_2769)
);

OAI22x1_ASAP7_75t_L g2770 ( 
.A1(n_2566),
.A2(n_2475),
.B1(n_2470),
.B2(n_2184),
.Y(n_2770)
);

AO21x1_ASAP7_75t_L g2771 ( 
.A1(n_2581),
.A2(n_2475),
.B(n_2470),
.Y(n_2771)
);

AOI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2591),
.A2(n_2121),
.B(n_1961),
.Y(n_2772)
);

BUFx2_ASAP7_75t_L g2773 ( 
.A(n_2696),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2659),
.B(n_2256),
.Y(n_2774)
);

A2O1A1Ixp33_ASAP7_75t_L g2775 ( 
.A1(n_2630),
.A2(n_2202),
.B(n_2149),
.C(n_2141),
.Y(n_2775)
);

CKINVDCx10_ASAP7_75t_R g2776 ( 
.A(n_2585),
.Y(n_2776)
);

AND2x2_ASAP7_75t_SL g2777 ( 
.A(n_2681),
.B(n_2330),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2591),
.A2(n_1961),
.B(n_2171),
.Y(n_2778)
);

AOI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2576),
.A2(n_2309),
.B1(n_2256),
.B2(n_2337),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2550),
.Y(n_2780)
);

OAI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2574),
.A2(n_2160),
.B1(n_2037),
.B2(n_2149),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2574),
.A2(n_2370),
.B1(n_2337),
.B2(n_2149),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2693),
.A2(n_2290),
.B(n_2299),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2630),
.A2(n_2664),
.B(n_2633),
.C(n_2700),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_L g2785 ( 
.A1(n_2693),
.A2(n_2299),
.B(n_2332),
.Y(n_2785)
);

INVxp67_ASAP7_75t_SL g2786 ( 
.A(n_2597),
.Y(n_2786)
);

O2A1O1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2658),
.A2(n_2082),
.B(n_2077),
.C(n_2078),
.Y(n_2787)
);

NOR2x1p5_ASAP7_75t_SL g2788 ( 
.A(n_2695),
.B(n_1940),
.Y(n_2788)
);

OAI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2633),
.A2(n_2370),
.B(n_2337),
.Y(n_2789)
);

A2O1A1Ixp33_ASAP7_75t_L g2790 ( 
.A1(n_2664),
.A2(n_2079),
.B(n_2184),
.C(n_2125),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2558),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2662),
.B(n_2330),
.Y(n_2792)
);

OR2x2_ASAP7_75t_L g2793 ( 
.A(n_2552),
.B(n_2380),
.Y(n_2793)
);

AOI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2571),
.A2(n_2554),
.B1(n_2688),
.B2(n_2671),
.Y(n_2794)
);

OR2x6_ASAP7_75t_SL g2795 ( 
.A(n_2644),
.B(n_2382),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_SL g2796 ( 
.A(n_2654),
.B(n_2334),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_2573),
.Y(n_2797)
);

AO21x1_ASAP7_75t_L g2798 ( 
.A1(n_2561),
.A2(n_2356),
.B(n_2052),
.Y(n_2798)
);

A2O1A1Ixp33_ASAP7_75t_SL g2799 ( 
.A1(n_2689),
.A2(n_2305),
.B(n_2312),
.C(n_2297),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2662),
.B(n_2334),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2665),
.B(n_2551),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2700),
.A2(n_2702),
.B(n_2697),
.C(n_2663),
.Y(n_2802)
);

AOI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2702),
.A2(n_1961),
.B(n_2125),
.Y(n_2803)
);

OAI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2698),
.A2(n_2557),
.B(n_2556),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2587),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2666),
.B(n_2334),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2685),
.B(n_2335),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_2665),
.B(n_2335),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2665),
.B(n_2335),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2685),
.A2(n_2370),
.B(n_2337),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2683),
.A2(n_2370),
.B1(n_2052),
.B2(n_2305),
.Y(n_2811)
);

OAI21x1_ASAP7_75t_L g2812 ( 
.A1(n_2656),
.A2(n_1619),
.B(n_1565),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2565),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2562),
.B(n_2345),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2575),
.A2(n_1932),
.B(n_1930),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2556),
.A2(n_1932),
.B(n_1930),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2559),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2557),
.A2(n_1930),
.B(n_2297),
.Y(n_2818)
);

CKINVDCx11_ASAP7_75t_R g2819 ( 
.A(n_2670),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2551),
.B(n_2192),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2667),
.A2(n_2052),
.B1(n_2320),
.B2(n_2312),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2598),
.A2(n_2336),
.B(n_2320),
.Y(n_2822)
);

O2A1O1Ixp33_ASAP7_75t_L g2823 ( 
.A1(n_2660),
.A2(n_2082),
.B(n_2077),
.C(n_2078),
.Y(n_2823)
);

NAND2xp33_ASAP7_75t_L g2824 ( 
.A(n_2598),
.B(n_2359),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2670),
.B(n_58),
.Y(n_2825)
);

AO22x1_ASAP7_75t_L g2826 ( 
.A1(n_2571),
.A2(n_2369),
.B1(n_2381),
.B2(n_2359),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2599),
.A2(n_2381),
.B(n_2359),
.Y(n_2827)
);

BUFx2_ASAP7_75t_L g2828 ( 
.A(n_2668),
.Y(n_2828)
);

AOI221xp5_ASAP7_75t_L g2829 ( 
.A1(n_2568),
.A2(n_1592),
.B1(n_1604),
.B2(n_1598),
.C(n_1584),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2580),
.B(n_2668),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2675),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2570),
.B(n_2381),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2583),
.B(n_2584),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2554),
.B(n_2651),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2589),
.Y(n_2835)
);

NAND2x1_ASAP7_75t_L g2836 ( 
.A(n_2571),
.B(n_2192),
.Y(n_2836)
);

NOR2x1p5_ASAP7_75t_SL g2837 ( 
.A(n_2592),
.B(n_2076),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2647),
.A2(n_1984),
.B(n_1952),
.Y(n_2838)
);

BUFx6f_ASAP7_75t_L g2839 ( 
.A(n_2580),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2598),
.A2(n_2203),
.B(n_2192),
.Y(n_2840)
);

AOI22x1_ASAP7_75t_L g2841 ( 
.A1(n_2689),
.A2(n_2203),
.B1(n_2211),
.B2(n_2192),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2651),
.B(n_2203),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2656),
.A2(n_2211),
.B(n_2203),
.Y(n_2843)
);

BUFx12f_ASAP7_75t_L g2844 ( 
.A(n_2694),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2647),
.A2(n_2650),
.B(n_2580),
.Y(n_2845)
);

BUFx6f_ASAP7_75t_L g2846 ( 
.A(n_2580),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2676),
.B(n_2211),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2564),
.Y(n_2848)
);

A2O1A1Ixp33_ASAP7_75t_L g2849 ( 
.A1(n_2652),
.A2(n_1959),
.B(n_2082),
.C(n_2029),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2593),
.B(n_2236),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2675),
.B(n_2236),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2601),
.B(n_2236),
.Y(n_2852)
);

A2O1A1Ixp33_ASAP7_75t_L g2853 ( 
.A1(n_2710),
.A2(n_2605),
.B(n_2637),
.C(n_2682),
.Y(n_2853)
);

OAI21xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2724),
.A2(n_2594),
.B(n_2637),
.Y(n_2854)
);

OAI22x1_ASAP7_75t_L g2855 ( 
.A1(n_2715),
.A2(n_2687),
.B1(n_2692),
.B2(n_2679),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2748),
.Y(n_2856)
);

AO21x1_ASAP7_75t_L g2857 ( 
.A1(n_2750),
.A2(n_2687),
.B(n_2679),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2714),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2726),
.A2(n_2571),
.B1(n_2671),
.B2(n_2640),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2704),
.A2(n_2614),
.B(n_2603),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2707),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2769),
.B(n_2675),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2706),
.B(n_2675),
.Y(n_2863)
);

OAI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2750),
.A2(n_2671),
.B(n_2640),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2719),
.B(n_2671),
.Y(n_2865)
);

OAI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2708),
.A2(n_2705),
.B(n_2728),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_SL g2867 ( 
.A(n_2733),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_SL g2868 ( 
.A1(n_2825),
.A2(n_2638),
.B(n_2631),
.Y(n_2868)
);

AOI211x1_ASAP7_75t_L g2869 ( 
.A1(n_2737),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_2869)
);

OAI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2708),
.A2(n_2671),
.B(n_2640),
.Y(n_2870)
);

OAI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2711),
.A2(n_2640),
.B(n_2571),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2733),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2712),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2833),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2716),
.B(n_2577),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2725),
.B(n_2577),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2761),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2740),
.B(n_2760),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2721),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2776),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2780),
.B(n_2615),
.Y(n_2881)
);

NOR4xp25_ASAP7_75t_L g2882 ( 
.A(n_2741),
.B(n_2625),
.C(n_2627),
.D(n_2624),
.Y(n_2882)
);

OAI22x1_ASAP7_75t_L g2883 ( 
.A1(n_2717),
.A2(n_2608),
.B1(n_2616),
.B2(n_2635),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2791),
.B(n_2835),
.Y(n_2884)
);

OAI22x1_ASAP7_75t_L g2885 ( 
.A1(n_2782),
.A2(n_2608),
.B1(n_2616),
.B2(n_2635),
.Y(n_2885)
);

NAND2xp33_ASAP7_75t_L g2886 ( 
.A(n_2813),
.B(n_2251),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2743),
.A2(n_2596),
.B1(n_1984),
.B2(n_2001),
.Y(n_2887)
);

OAI21x1_ASAP7_75t_L g2888 ( 
.A1(n_2754),
.A2(n_2629),
.B(n_1565),
.Y(n_2888)
);

OAI21x1_ASAP7_75t_SL g2889 ( 
.A1(n_2732),
.A2(n_66),
.B(n_67),
.Y(n_2889)
);

AO31x2_ASAP7_75t_L g2890 ( 
.A1(n_2798),
.A2(n_2775),
.A3(n_2770),
.B(n_2810),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2779),
.A2(n_2251),
.B1(n_1993),
.B2(n_2001),
.Y(n_2891)
);

AOI211x1_ASAP7_75t_L g2892 ( 
.A1(n_2720),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2819),
.B(n_69),
.Y(n_2893)
);

A2O1A1Ixp33_ASAP7_75t_L g2894 ( 
.A1(n_2756),
.A2(n_1959),
.B(n_2185),
.C(n_2178),
.Y(n_2894)
);

AO31x2_ASAP7_75t_L g2895 ( 
.A1(n_2810),
.A2(n_2214),
.A3(n_2222),
.B(n_2208),
.Y(n_2895)
);

OAI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2711),
.A2(n_1604),
.B(n_1598),
.Y(n_2896)
);

OAI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2757),
.A2(n_1608),
.B(n_1607),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2736),
.B(n_71),
.Y(n_2898)
);

OAI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2757),
.A2(n_1613),
.B(n_1611),
.Y(n_2899)
);

A2O1A1Ixp33_ASAP7_75t_L g2900 ( 
.A1(n_2768),
.A2(n_2185),
.B(n_2178),
.C(n_2029),
.Y(n_2900)
);

AO31x2_ASAP7_75t_L g2901 ( 
.A1(n_2803),
.A2(n_2243),
.A3(n_2246),
.B(n_2222),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2789),
.A2(n_2012),
.B(n_1952),
.Y(n_2902)
);

INVx5_ASAP7_75t_L g2903 ( 
.A(n_2733),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2795),
.B(n_2735),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2747),
.B(n_72),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2765),
.Y(n_2906)
);

OA21x2_ASAP7_75t_L g2907 ( 
.A1(n_2845),
.A2(n_2289),
.B(n_2247),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2797),
.B(n_72),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2764),
.B(n_74),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2738),
.Y(n_2910)
);

OA22x2_ASAP7_75t_L g2911 ( 
.A1(n_2729),
.A2(n_2365),
.B1(n_2343),
.B2(n_2346),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2824),
.A2(n_2012),
.B(n_1952),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2777),
.A2(n_1993),
.B1(n_2017),
.B2(n_2012),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2727),
.A2(n_2826),
.B(n_2800),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2744),
.B(n_75),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2722),
.B(n_77),
.Y(n_2916)
);

AOI21x1_ASAP7_75t_SL g2917 ( 
.A1(n_2814),
.A2(n_77),
.B(n_80),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2786),
.B(n_80),
.Y(n_2918)
);

OAI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2763),
.A2(n_1613),
.B(n_1611),
.Y(n_2919)
);

INVx5_ASAP7_75t_SL g2920 ( 
.A(n_2765),
.Y(n_2920)
);

OAI21x1_ASAP7_75t_L g2921 ( 
.A1(n_2730),
.A2(n_2365),
.B(n_2349),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2742),
.Y(n_2922)
);

AO22x2_ASAP7_75t_L g2923 ( 
.A1(n_2767),
.A2(n_2349),
.B1(n_2023),
.B2(n_2034),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2834),
.B(n_82),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2773),
.B(n_83),
.Y(n_2925)
);

CKINVDCx10_ASAP7_75t_R g2926 ( 
.A(n_2731),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2828),
.B(n_1993),
.Y(n_2927)
);

O2A1O1Ixp5_ASAP7_75t_L g2928 ( 
.A1(n_2830),
.A2(n_2023),
.B(n_2044),
.C(n_2034),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2793),
.B(n_84),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2765),
.B(n_2065),
.Y(n_2930)
);

AOI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2792),
.A2(n_2017),
.B(n_2100),
.Y(n_2931)
);

OAI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2763),
.A2(n_1628),
.B(n_1622),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2713),
.A2(n_1993),
.B1(n_2044),
.B2(n_2034),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2749),
.A2(n_1628),
.B(n_1622),
.Y(n_2934)
);

BUFx2_ASAP7_75t_L g2935 ( 
.A(n_2844),
.Y(n_2935)
);

AOI21xp5_ASAP7_75t_L g2936 ( 
.A1(n_2778),
.A2(n_2107),
.B(n_2100),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2852),
.B(n_85),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2850),
.B(n_85),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2709),
.Y(n_2939)
);

OAI21x1_ASAP7_75t_SL g2940 ( 
.A1(n_2771),
.A2(n_86),
.B(n_87),
.Y(n_2940)
);

INVx5_ASAP7_75t_L g2941 ( 
.A(n_2839),
.Y(n_2941)
);

BUFx3_ASAP7_75t_L g2942 ( 
.A(n_2805),
.Y(n_2942)
);

BUFx12f_ASAP7_75t_L g2943 ( 
.A(n_2753),
.Y(n_2943)
);

OAI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2766),
.A2(n_1635),
.B(n_1633),
.Y(n_2944)
);

OAI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2781),
.A2(n_1635),
.B(n_1633),
.Y(n_2945)
);

AO31x2_ASAP7_75t_L g2946 ( 
.A1(n_2803),
.A2(n_2112),
.A3(n_2115),
.B(n_2110),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2806),
.B(n_89),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2807),
.B(n_90),
.Y(n_2948)
);

OAI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2758),
.A2(n_1993),
.B1(n_2080),
.B2(n_2110),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2739),
.B(n_90),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2832),
.Y(n_2951)
);

OR2x6_ASAP7_75t_L g2952 ( 
.A(n_2836),
.B(n_2845),
.Y(n_2952)
);

AO31x2_ASAP7_75t_L g2953 ( 
.A1(n_2802),
.A2(n_2112),
.A3(n_2122),
.B(n_2115),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_L g2954 ( 
.A(n_2762),
.B(n_92),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2709),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2784),
.B(n_93),
.Y(n_2956)
);

OR2x2_ASAP7_75t_L g2957 ( 
.A(n_2745),
.B(n_94),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2841),
.A2(n_2127),
.B(n_2122),
.Y(n_2958)
);

CKINVDCx20_ASAP7_75t_R g2959 ( 
.A(n_2746),
.Y(n_2959)
);

OAI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2723),
.A2(n_2128),
.B1(n_2129),
.B2(n_2127),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2759),
.A2(n_2129),
.B1(n_2143),
.B2(n_2128),
.Y(n_2961)
);

INVx4_ASAP7_75t_L g2962 ( 
.A(n_2839),
.Y(n_2962)
);

OAI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2838),
.A2(n_2144),
.B(n_2143),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2723),
.A2(n_2146),
.B1(n_2144),
.B2(n_2150),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2774),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2817),
.Y(n_2966)
);

AOI21x1_ASAP7_75t_SL g2967 ( 
.A1(n_2842),
.A2(n_94),
.B(n_95),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_SL g2968 ( 
.A1(n_2794),
.A2(n_95),
.B(n_97),
.Y(n_2968)
);

NAND3xp33_ASAP7_75t_L g2969 ( 
.A(n_2718),
.B(n_1638),
.C(n_1636),
.Y(n_2969)
);

OAI21x1_ASAP7_75t_L g2970 ( 
.A1(n_2785),
.A2(n_1544),
.B(n_1520),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_SL g2971 ( 
.A1(n_2804),
.A2(n_99),
.B(n_100),
.Y(n_2971)
);

OAI21x1_ASAP7_75t_SL g2972 ( 
.A1(n_2811),
.A2(n_100),
.B(n_101),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2847),
.B(n_102),
.Y(n_2973)
);

NOR2x1_ASAP7_75t_SL g2974 ( 
.A(n_2801),
.B(n_951),
.Y(n_2974)
);

AOI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2816),
.A2(n_1858),
.B(n_1857),
.Y(n_2975)
);

AO31x2_ASAP7_75t_L g2976 ( 
.A1(n_2783),
.A2(n_1520),
.A3(n_1544),
.B(n_1591),
.Y(n_2976)
);

OAI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2751),
.A2(n_1544),
.B(n_1520),
.Y(n_2977)
);

BUFx3_ASAP7_75t_L g2978 ( 
.A(n_2734),
.Y(n_2978)
);

AOI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2816),
.A2(n_1595),
.B(n_1591),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2752),
.B(n_102),
.Y(n_2980)
);

NAND2x1p5_ASAP7_75t_L g2981 ( 
.A(n_2839),
.B(n_1636),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2755),
.B(n_105),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2734),
.B(n_105),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2831),
.B(n_2846),
.Y(n_2984)
);

BUFx10_ASAP7_75t_L g2985 ( 
.A(n_2846),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_SL g2986 ( 
.A1(n_2822),
.A2(n_106),
.B(n_108),
.Y(n_2986)
);

OR2x2_ASAP7_75t_L g2987 ( 
.A(n_2848),
.B(n_109),
.Y(n_2987)
);

BUFx3_ASAP7_75t_L g2988 ( 
.A(n_2846),
.Y(n_2988)
);

OAI21x1_ASAP7_75t_L g2989 ( 
.A1(n_2812),
.A2(n_1595),
.B(n_1591),
.Y(n_2989)
);

BUFx4_ASAP7_75t_SL g2990 ( 
.A(n_2796),
.Y(n_2990)
);

BUFx12f_ASAP7_75t_L g2991 ( 
.A(n_2840),
.Y(n_2991)
);

AO32x2_ASAP7_75t_L g2992 ( 
.A1(n_2821),
.A2(n_109),
.A3(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_2992)
);

AO31x2_ASAP7_75t_L g2993 ( 
.A1(n_2790),
.A2(n_1595),
.A3(n_1625),
.B(n_1620),
.Y(n_2993)
);

OAI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2787),
.A2(n_111),
.B(n_112),
.Y(n_2994)
);

AND2x4_ASAP7_75t_L g2995 ( 
.A(n_2837),
.B(n_115),
.Y(n_2995)
);

BUFx12f_ASAP7_75t_L g2996 ( 
.A(n_2827),
.Y(n_2996)
);

OAI21x1_ASAP7_75t_L g2997 ( 
.A1(n_2772),
.A2(n_1620),
.B(n_1595),
.Y(n_2997)
);

AND2x4_ASAP7_75t_L g2998 ( 
.A(n_2788),
.B(n_116),
.Y(n_2998)
);

INVx5_ASAP7_75t_SL g2999 ( 
.A(n_2851),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2843),
.B(n_117),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2823),
.A2(n_118),
.B(n_119),
.Y(n_3001)
);

OAI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2849),
.A2(n_119),
.B(n_121),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2815),
.A2(n_1625),
.B(n_1620),
.Y(n_3003)
);

OR2x2_ASAP7_75t_L g3004 ( 
.A(n_2820),
.B(n_122),
.Y(n_3004)
);

AO32x2_ASAP7_75t_L g3005 ( 
.A1(n_2799),
.A2(n_123),
.A3(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2827),
.B(n_1636),
.Y(n_3006)
);

OAI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2818),
.A2(n_123),
.B(n_124),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2808),
.B(n_125),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2809),
.B(n_127),
.Y(n_3009)
);

OAI21x1_ASAP7_75t_L g3010 ( 
.A1(n_2815),
.A2(n_1625),
.B(n_1620),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2829),
.Y(n_3011)
);

BUFx4_ASAP7_75t_SL g3012 ( 
.A(n_2880),
.Y(n_3012)
);

A2O1A1Ixp33_ASAP7_75t_L g3013 ( 
.A1(n_2968),
.A2(n_2818),
.B(n_130),
.C(n_128),
.Y(n_3013)
);

AOI21xp5_ASAP7_75t_L g3014 ( 
.A1(n_2864),
.A2(n_1625),
.B(n_1620),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2942),
.Y(n_3015)
);

INVx5_ASAP7_75t_L g3016 ( 
.A(n_2996),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2884),
.Y(n_3017)
);

O2A1O1Ixp33_ASAP7_75t_L g3018 ( 
.A1(n_2956),
.A2(n_133),
.B(n_129),
.C(n_132),
.Y(n_3018)
);

O2A1O1Ixp33_ASAP7_75t_SL g3019 ( 
.A1(n_2868),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_3019)
);

OAI21xp33_ASAP7_75t_SL g3020 ( 
.A1(n_2866),
.A2(n_138),
.B(n_139),
.Y(n_3020)
);

O2A1O1Ixp33_ASAP7_75t_L g3021 ( 
.A1(n_3007),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_3021)
);

OAI21x1_ASAP7_75t_L g3022 ( 
.A1(n_2914),
.A2(n_140),
.B(n_143),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2871),
.A2(n_1626),
.B(n_1625),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2870),
.A2(n_1626),
.B(n_1636),
.Y(n_3024)
);

AOI221x1_ASAP7_75t_L g3025 ( 
.A1(n_2940),
.A2(n_999),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2870),
.A2(n_2969),
.B(n_2896),
.Y(n_3026)
);

OAI21xp33_ASAP7_75t_L g3027 ( 
.A1(n_3007),
.A2(n_144),
.B(n_146),
.Y(n_3027)
);

OAI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2968),
.A2(n_144),
.B(n_149),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2861),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_3011),
.A2(n_1659),
.B1(n_1640),
.B2(n_1639),
.Y(n_3030)
);

AO31x2_ASAP7_75t_L g3031 ( 
.A1(n_2885),
.A2(n_150),
.A3(n_151),
.B(n_152),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2858),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2873),
.Y(n_3033)
);

INVx3_ASAP7_75t_SL g3034 ( 
.A(n_2959),
.Y(n_3034)
);

AOI221x1_ASAP7_75t_L g3035 ( 
.A1(n_2916),
.A2(n_999),
.B1(n_151),
.B2(n_152),
.C(n_153),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2969),
.A2(n_1626),
.B(n_1636),
.Y(n_3036)
);

AOI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2896),
.A2(n_1626),
.B(n_1638),
.Y(n_3037)
);

OAI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_3002),
.A2(n_154),
.B(n_155),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2892),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_3039)
);

AND2x4_ASAP7_75t_SL g3040 ( 
.A(n_2985),
.B(n_999),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2945),
.A2(n_1626),
.B(n_1638),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2978),
.Y(n_3042)
);

BUFx10_ASAP7_75t_L g3043 ( 
.A(n_2980),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2877),
.Y(n_3044)
);

BUFx10_ASAP7_75t_L g3045 ( 
.A(n_2982),
.Y(n_3045)
);

INVx2_ASAP7_75t_SL g3046 ( 
.A(n_2935),
.Y(n_3046)
);

AO21x1_ASAP7_75t_L g3047 ( 
.A1(n_2904),
.A2(n_161),
.B(n_162),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2945),
.A2(n_1639),
.B(n_1638),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2943),
.Y(n_3049)
);

AO31x2_ASAP7_75t_L g3050 ( 
.A1(n_2876),
.A2(n_162),
.A3(n_164),
.B(n_167),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2951),
.B(n_164),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2892),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_3052)
);

O2A1O1Ixp33_ASAP7_75t_L g3053 ( 
.A1(n_3002),
.A2(n_168),
.B(n_170),
.C(n_171),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2874),
.B(n_171),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2879),
.Y(n_3055)
);

OAI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2869),
.A2(n_172),
.B1(n_173),
.B2(n_176),
.Y(n_3056)
);

BUFx8_ASAP7_75t_L g3057 ( 
.A(n_2925),
.Y(n_3057)
);

NOR4xp25_ASAP7_75t_L g3058 ( 
.A(n_2868),
.B(n_172),
.C(n_173),
.D(n_176),
.Y(n_3058)
);

AO32x2_ASAP7_75t_L g3059 ( 
.A1(n_2887),
.A2(n_177),
.A3(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2862),
.B(n_178),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2897),
.A2(n_1640),
.B(n_1639),
.Y(n_3061)
);

A2O1A1Ixp33_ASAP7_75t_L g3062 ( 
.A1(n_2854),
.A2(n_181),
.B(n_182),
.C(n_183),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2856),
.Y(n_3063)
);

O2A1O1Ixp33_ASAP7_75t_L g3064 ( 
.A1(n_2918),
.A2(n_182),
.B(n_184),
.C(n_185),
.Y(n_3064)
);

INVx2_ASAP7_75t_SL g3065 ( 
.A(n_2985),
.Y(n_3065)
);

OAI21x1_ASAP7_75t_L g3066 ( 
.A1(n_2860),
.A2(n_184),
.B(n_185),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2897),
.A2(n_1659),
.B(n_1640),
.Y(n_3067)
);

AOI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2899),
.A2(n_2932),
.B(n_2919),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2881),
.Y(n_3069)
);

BUFx2_ASAP7_75t_R g3070 ( 
.A(n_2988),
.Y(n_3070)
);

INVx5_ASAP7_75t_SL g3071 ( 
.A(n_2872),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2899),
.A2(n_1659),
.B(n_1640),
.Y(n_3072)
);

CKINVDCx20_ASAP7_75t_R g3073 ( 
.A(n_2915),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_2926),
.Y(n_3074)
);

O2A1O1Ixp33_ASAP7_75t_SL g3075 ( 
.A1(n_2893),
.A2(n_186),
.B(n_187),
.C(n_189),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2872),
.Y(n_3076)
);

AOI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2937),
.A2(n_190),
.B(n_191),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2919),
.A2(n_1659),
.B(n_1428),
.Y(n_3078)
);

AND2x4_ASAP7_75t_L g3079 ( 
.A(n_2965),
.B(n_192),
.Y(n_3079)
);

INVx4_ASAP7_75t_L g3080 ( 
.A(n_2872),
.Y(n_3080)
);

OAI21x1_ASAP7_75t_L g3081 ( 
.A1(n_2997),
.A2(n_193),
.B(n_194),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2853),
.A2(n_1659),
.B(n_193),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2878),
.B(n_196),
.Y(n_3083)
);

AO32x2_ASAP7_75t_L g3084 ( 
.A1(n_2887),
.A2(n_197),
.A3(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2926),
.B(n_200),
.Y(n_3085)
);

NOR2xp67_ASAP7_75t_L g3086 ( 
.A(n_2883),
.B(n_2854),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_2984),
.Y(n_3087)
);

AOI21xp5_ASAP7_75t_L g3088 ( 
.A1(n_2886),
.A2(n_202),
.B(n_203),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2859),
.A2(n_204),
.B(n_205),
.C(n_206),
.Y(n_3089)
);

NOR2xp33_ASAP7_75t_L g3090 ( 
.A(n_2954),
.B(n_207),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2979),
.A2(n_213),
.B(n_214),
.Y(n_3091)
);

OAI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_2869),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2875),
.B(n_215),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2921),
.A2(n_219),
.B(n_221),
.Y(n_3094)
);

A2O1A1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2859),
.A2(n_219),
.B(n_222),
.C(n_223),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2994),
.A2(n_223),
.B(n_226),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2863),
.B(n_226),
.Y(n_3097)
);

BUFx2_ASAP7_75t_L g3098 ( 
.A(n_2939),
.Y(n_3098)
);

OAI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_3001),
.A2(n_227),
.B(n_228),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2955),
.B(n_228),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_3001),
.A2(n_229),
.B(n_230),
.Y(n_3101)
);

INVx1_ASAP7_75t_SL g3102 ( 
.A(n_2990),
.Y(n_3102)
);

CKINVDCx11_ASAP7_75t_R g3103 ( 
.A(n_2991),
.Y(n_3103)
);

NAND2x1p5_ASAP7_75t_L g3104 ( 
.A(n_2903),
.B(n_231),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_3006),
.A2(n_231),
.B(n_233),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2957),
.B(n_233),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2962),
.Y(n_3107)
);

OAI21x1_ASAP7_75t_L g3108 ( 
.A1(n_2934),
.A2(n_234),
.B(n_235),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2950),
.A2(n_235),
.B(n_236),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2905),
.B(n_236),
.Y(n_3110)
);

OAI21x1_ASAP7_75t_L g3111 ( 
.A1(n_2934),
.A2(n_237),
.B(n_238),
.Y(n_3111)
);

AO31x2_ASAP7_75t_L g3112 ( 
.A1(n_2857),
.A2(n_238),
.A3(n_239),
.B(n_242),
.Y(n_3112)
);

OAI22xp5_ASAP7_75t_L g3113 ( 
.A1(n_3004),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_3113)
);

AOI21x1_ASAP7_75t_L g3114 ( 
.A1(n_2938),
.A2(n_244),
.B(n_245),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_L g3115 ( 
.A(n_2903),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2865),
.B(n_245),
.Y(n_3116)
);

A2O1A1Ixp33_ASAP7_75t_L g3117 ( 
.A1(n_2908),
.A2(n_246),
.B(n_248),
.C(n_249),
.Y(n_3117)
);

INVx1_ASAP7_75t_SL g3118 ( 
.A(n_2924),
.Y(n_3118)
);

AND2x4_ASAP7_75t_L g3119 ( 
.A(n_2952),
.B(n_246),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2929),
.B(n_250),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2910),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2944),
.A2(n_251),
.B(n_252),
.Y(n_3122)
);

INVx5_ASAP7_75t_L g3123 ( 
.A(n_2952),
.Y(n_3123)
);

CKINVDCx20_ASAP7_75t_R g3124 ( 
.A(n_2973),
.Y(n_3124)
);

AO31x2_ASAP7_75t_L g3125 ( 
.A1(n_2933),
.A2(n_251),
.A3(n_253),
.B(n_254),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2898),
.B(n_253),
.Y(n_3126)
);

O2A1O1Ixp33_ASAP7_75t_L g3127 ( 
.A1(n_2889),
.A2(n_255),
.B(n_256),
.C(n_257),
.Y(n_3127)
);

BUFx6f_ASAP7_75t_L g3128 ( 
.A(n_2903),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2909),
.B(n_256),
.Y(n_3129)
);

A2O1A1Ixp33_ASAP7_75t_L g3130 ( 
.A1(n_2995),
.A2(n_259),
.B(n_260),
.C(n_261),
.Y(n_3130)
);

NOR2x1_ASAP7_75t_SL g3131 ( 
.A(n_2952),
.B(n_259),
.Y(n_3131)
);

AO31x2_ASAP7_75t_L g3132 ( 
.A1(n_2949),
.A2(n_262),
.A3(n_263),
.B(n_264),
.Y(n_3132)
);

O2A1O1Ixp33_ASAP7_75t_SL g3133 ( 
.A1(n_3008),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2894),
.A2(n_265),
.B(n_266),
.Y(n_3134)
);

OAI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_3000),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_3135)
);

BUFx2_ASAP7_75t_R g3136 ( 
.A(n_2906),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2911),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2947),
.B(n_269),
.Y(n_3138)
);

BUFx6f_ASAP7_75t_L g3139 ( 
.A(n_2941),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2948),
.B(n_270),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2966),
.Y(n_3141)
);

NAND3xp33_ASAP7_75t_L g3142 ( 
.A(n_3009),
.B(n_271),
.C(n_273),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2922),
.B(n_274),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3087),
.B(n_2920),
.Y(n_3144)
);

OAI22xp33_ASAP7_75t_L g3145 ( 
.A1(n_3028),
.A2(n_2987),
.B1(n_2855),
.B2(n_2992),
.Y(n_3145)
);

OAI221xp5_ASAP7_75t_L g3146 ( 
.A1(n_3109),
.A2(n_2882),
.B1(n_2964),
.B2(n_2992),
.C(n_2961),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_3038),
.A2(n_2971),
.B1(n_2972),
.B2(n_2995),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_3013),
.A2(n_2998),
.B1(n_2999),
.B2(n_2992),
.Y(n_3148)
);

BUFx2_ASAP7_75t_L g3149 ( 
.A(n_3098),
.Y(n_3149)
);

OAI211xp5_ASAP7_75t_SL g3150 ( 
.A1(n_3090),
.A2(n_2930),
.B(n_2967),
.C(n_2917),
.Y(n_3150)
);

HB1xp67_ASAP7_75t_L g3151 ( 
.A(n_3032),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_3012),
.Y(n_3152)
);

OAI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_3058),
.A2(n_3062),
.B(n_3026),
.Y(n_3153)
);

AOI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_3068),
.A2(n_2928),
.B(n_2975),
.Y(n_3154)
);

BUFx2_ASAP7_75t_L g3155 ( 
.A(n_3034),
.Y(n_3155)
);

OA21x2_ASAP7_75t_L g3156 ( 
.A1(n_3086),
.A2(n_2989),
.B(n_2888),
.Y(n_3156)
);

OAI22x1_ASAP7_75t_L g3157 ( 
.A1(n_3079),
.A2(n_3118),
.B1(n_3119),
.B2(n_3046),
.Y(n_3157)
);

BUFx3_ASAP7_75t_L g3158 ( 
.A(n_3015),
.Y(n_3158)
);

CKINVDCx12_ASAP7_75t_R g3159 ( 
.A(n_3110),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_3027),
.A2(n_2913),
.B1(n_2891),
.B2(n_2923),
.Y(n_3160)
);

INVx1_ASAP7_75t_SL g3161 ( 
.A(n_3074),
.Y(n_3161)
);

BUFx4f_ASAP7_75t_L g3162 ( 
.A(n_3104),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_3023),
.A2(n_3036),
.B(n_3014),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3020),
.A2(n_2983),
.B(n_2902),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_3043),
.B(n_2906),
.Y(n_3165)
);

AND2x4_ASAP7_75t_L g3166 ( 
.A(n_3123),
.B(n_2890),
.Y(n_3166)
);

AO21x2_ASAP7_75t_L g3167 ( 
.A1(n_3116),
.A2(n_2963),
.B(n_2986),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_3024),
.A2(n_2900),
.B(n_2936),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3069),
.Y(n_3169)
);

NAND3xp33_ASAP7_75t_L g3170 ( 
.A(n_3064),
.B(n_2931),
.C(n_2964),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3047),
.A2(n_2960),
.B1(n_2961),
.B2(n_2963),
.Y(n_3171)
);

AND2x4_ASAP7_75t_L g3172 ( 
.A(n_3123),
.B(n_2890),
.Y(n_3172)
);

AND2x2_ASAP7_75t_L g3173 ( 
.A(n_3042),
.B(n_2920),
.Y(n_3173)
);

OA21x2_ASAP7_75t_L g3174 ( 
.A1(n_3063),
.A2(n_3010),
.B(n_3003),
.Y(n_3174)
);

OR2x6_ASAP7_75t_L g3175 ( 
.A(n_3119),
.B(n_2927),
.Y(n_3175)
);

BUFx3_ASAP7_75t_L g3176 ( 
.A(n_3049),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3029),
.Y(n_3177)
);

O2A1O1Ixp33_ASAP7_75t_SL g3178 ( 
.A1(n_3102),
.A2(n_3005),
.B(n_2912),
.C(n_2999),
.Y(n_3178)
);

OA21x2_ASAP7_75t_L g3179 ( 
.A1(n_3051),
.A2(n_3017),
.B(n_3044),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3121),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_3033),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_3043),
.B(n_2941),
.Y(n_3182)
);

NOR2x1_ASAP7_75t_SL g3183 ( 
.A(n_3016),
.B(n_3123),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_3136),
.Y(n_3184)
);

AND2x4_ASAP7_75t_L g3185 ( 
.A(n_3042),
.B(n_2890),
.Y(n_3185)
);

OAI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3107),
.A2(n_2907),
.B(n_2958),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_3099),
.A2(n_3005),
.B1(n_2977),
.B2(n_2867),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3089),
.A2(n_2941),
.B1(n_2981),
.B2(n_2977),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_3050),
.Y(n_3189)
);

AOI221xp5_ASAP7_75t_L g3190 ( 
.A1(n_3075),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.C(n_278),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_3082),
.A2(n_2974),
.B(n_2970),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3055),
.Y(n_3192)
);

NOR2xp67_ASAP7_75t_L g3193 ( 
.A(n_3016),
.B(n_276),
.Y(n_3193)
);

OAI22x1_ASAP7_75t_L g3194 ( 
.A1(n_3079),
.A2(n_2993),
.B1(n_2895),
.B2(n_2946),
.Y(n_3194)
);

AO21x2_ASAP7_75t_L g3195 ( 
.A1(n_3143),
.A2(n_2976),
.B(n_2895),
.Y(n_3195)
);

A2O1A1Ixp33_ASAP7_75t_L g3196 ( 
.A1(n_3053),
.A2(n_2993),
.B(n_279),
.C(n_280),
.Y(n_3196)
);

OR2x6_ASAP7_75t_L g3197 ( 
.A(n_3115),
.B(n_3128),
.Y(n_3197)
);

NAND2x1p5_ASAP7_75t_L g3198 ( 
.A(n_3016),
.B(n_2953),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_SL g3199 ( 
.A(n_3070),
.B(n_2953),
.Y(n_3199)
);

AO31x2_ASAP7_75t_L g3200 ( 
.A1(n_3131),
.A2(n_2901),
.A3(n_2953),
.B(n_2976),
.Y(n_3200)
);

BUFx2_ASAP7_75t_L g3201 ( 
.A(n_3065),
.Y(n_3201)
);

BUFx3_ASAP7_75t_L g3202 ( 
.A(n_3057),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_R g3203 ( 
.A(n_3124),
.B(n_278),
.Y(n_3203)
);

NOR2xp67_ASAP7_75t_L g3204 ( 
.A(n_3142),
.B(n_279),
.Y(n_3204)
);

AO31x2_ASAP7_75t_L g3205 ( 
.A1(n_3039),
.A2(n_2976),
.A3(n_281),
.B(n_282),
.Y(n_3205)
);

BUFx2_ASAP7_75t_R g3206 ( 
.A(n_3106),
.Y(n_3206)
);

BUFx3_ASAP7_75t_L g3207 ( 
.A(n_3057),
.Y(n_3207)
);

OR2x6_ASAP7_75t_SL g3208 ( 
.A(n_3083),
.B(n_280),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_3141),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_3054),
.B(n_3050),
.Y(n_3210)
);

OAI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_3137),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_3211)
);

CKINVDCx20_ASAP7_75t_R g3212 ( 
.A(n_3103),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3050),
.B(n_3093),
.Y(n_3213)
);

NOR2xp67_ASAP7_75t_L g3214 ( 
.A(n_3138),
.B(n_285),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_3045),
.B(n_3140),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3097),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_SL g3217 ( 
.A1(n_3052),
.A2(n_286),
.B1(n_293),
.B2(n_294),
.Y(n_3217)
);

NOR3xp33_ASAP7_75t_L g3218 ( 
.A(n_3117),
.B(n_286),
.C(n_298),
.Y(n_3218)
);

AO31x2_ASAP7_75t_L g3219 ( 
.A1(n_3056),
.A2(n_299),
.A3(n_311),
.B(n_313),
.Y(n_3219)
);

OAI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_3096),
.A2(n_315),
.B(n_316),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3115),
.Y(n_3221)
);

AND2x4_ASAP7_75t_L g3222 ( 
.A(n_3080),
.B(n_318),
.Y(n_3222)
);

OR2x6_ASAP7_75t_L g3223 ( 
.A(n_3115),
.B(n_319),
.Y(n_3223)
);

NOR2x1_ASAP7_75t_SL g3224 ( 
.A(n_3128),
.B(n_321),
.Y(n_3224)
);

AO31x2_ASAP7_75t_L g3225 ( 
.A1(n_3092),
.A2(n_3035),
.A3(n_3025),
.B(n_3101),
.Y(n_3225)
);

BUFx3_ASAP7_75t_L g3226 ( 
.A(n_3073),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3100),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3112),
.B(n_433),
.Y(n_3228)
);

OAI221xp5_ASAP7_75t_L g3229 ( 
.A1(n_3018),
.A2(n_323),
.B1(n_327),
.B2(n_329),
.C(n_331),
.Y(n_3229)
);

O2A1O1Ixp33_ASAP7_75t_L g3230 ( 
.A1(n_3019),
.A2(n_335),
.B(n_340),
.C(n_343),
.Y(n_3230)
);

AOI21xp33_ASAP7_75t_L g3231 ( 
.A1(n_3021),
.A2(n_345),
.B(n_349),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_3045),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3112),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_3060),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_3076),
.Y(n_3235)
);

OA21x2_ASAP7_75t_L g3236 ( 
.A1(n_3066),
.A2(n_354),
.B(n_361),
.Y(n_3236)
);

HB1xp67_ASAP7_75t_L g3237 ( 
.A(n_3112),
.Y(n_3237)
);

OA21x2_ASAP7_75t_L g3238 ( 
.A1(n_3022),
.A2(n_370),
.B(n_372),
.Y(n_3238)
);

AOI22xp33_ASAP7_75t_SL g3239 ( 
.A1(n_3126),
.A2(n_3113),
.B1(n_3135),
.B2(n_3122),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_3129),
.B(n_373),
.Y(n_3240)
);

OAI222xp33_ASAP7_75t_L g3241 ( 
.A1(n_3077),
.A2(n_376),
.B1(n_382),
.B2(n_384),
.C1(n_385),
.C2(n_386),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_3152),
.Y(n_3242)
);

AO31x2_ASAP7_75t_L g3243 ( 
.A1(n_3213),
.A2(n_3095),
.A3(n_3130),
.B(n_3120),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3179),
.B(n_3132),
.Y(n_3244)
);

AOI21x1_ASAP7_75t_L g3245 ( 
.A1(n_3155),
.A2(n_3114),
.B(n_3041),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3151),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3179),
.B(n_3132),
.Y(n_3247)
);

AO21x2_ASAP7_75t_L g3248 ( 
.A1(n_3189),
.A2(n_3134),
.B(n_3088),
.Y(n_3248)
);

CKINVDCx20_ASAP7_75t_R g3249 ( 
.A(n_3212),
.Y(n_3249)
);

OR2x6_ASAP7_75t_L g3250 ( 
.A(n_3198),
.B(n_3139),
.Y(n_3250)
);

OAI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3153),
.A2(n_3127),
.B(n_3091),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3178),
.A2(n_3133),
.B(n_3048),
.Y(n_3252)
);

CKINVDCx6p67_ASAP7_75t_R g3253 ( 
.A(n_3202),
.Y(n_3253)
);

OA21x2_ASAP7_75t_L g3254 ( 
.A1(n_3213),
.A2(n_3094),
.B(n_3081),
.Y(n_3254)
);

OAI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3148),
.A2(n_3105),
.B(n_3085),
.Y(n_3255)
);

CKINVDCx11_ASAP7_75t_R g3256 ( 
.A(n_3208),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3168),
.A2(n_3037),
.B(n_3061),
.Y(n_3257)
);

OA21x2_ASAP7_75t_L g3258 ( 
.A1(n_3210),
.A2(n_3030),
.B(n_3072),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3149),
.B(n_3071),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3173),
.B(n_3071),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3148),
.A2(n_3108),
.B(n_3111),
.Y(n_3261)
);

OA21x2_ASAP7_75t_L g3262 ( 
.A1(n_3210),
.A2(n_3067),
.B(n_3078),
.Y(n_3262)
);

BUFx2_ASAP7_75t_L g3263 ( 
.A(n_3226),
.Y(n_3263)
);

INVx2_ASAP7_75t_SL g3264 ( 
.A(n_3207),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3175),
.B(n_3183),
.Y(n_3265)
);

BUFx3_ASAP7_75t_L g3266 ( 
.A(n_3158),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3169),
.B(n_3125),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3189),
.B(n_3125),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3168),
.A2(n_3163),
.B(n_3154),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3180),
.B(n_3125),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3175),
.B(n_3080),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_3176),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_3175),
.B(n_3139),
.Y(n_3273)
);

AO31x2_ASAP7_75t_L g3274 ( 
.A1(n_3233),
.A2(n_3084),
.A3(n_3059),
.B(n_3031),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3237),
.B(n_3031),
.Y(n_3275)
);

AO21x2_ASAP7_75t_L g3276 ( 
.A1(n_3228),
.A2(n_3084),
.B(n_3059),
.Y(n_3276)
);

OA21x2_ASAP7_75t_L g3277 ( 
.A1(n_3185),
.A2(n_3084),
.B(n_3059),
.Y(n_3277)
);

OAI21x1_ASAP7_75t_L g3278 ( 
.A1(n_3186),
.A2(n_3139),
.B(n_3128),
.Y(n_3278)
);

OAI221xp5_ASAP7_75t_SL g3279 ( 
.A1(n_3239),
.A2(n_3076),
.B1(n_3040),
.B2(n_392),
.C(n_393),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3177),
.Y(n_3280)
);

AOI21xp33_ASAP7_75t_SL g3281 ( 
.A1(n_3157),
.A2(n_3076),
.B(n_391),
.Y(n_3281)
);

AO21x1_ASAP7_75t_L g3282 ( 
.A1(n_3145),
.A2(n_399),
.B(n_402),
.Y(n_3282)
);

OAI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3145),
.A2(n_403),
.B(n_406),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3201),
.B(n_408),
.Y(n_3284)
);

A2O1A1Ixp33_ASAP7_75t_L g3285 ( 
.A1(n_3204),
.A2(n_409),
.B(n_410),
.C(n_412),
.Y(n_3285)
);

CKINVDCx20_ASAP7_75t_R g3286 ( 
.A(n_3159),
.Y(n_3286)
);

BUFx8_ASAP7_75t_L g3287 ( 
.A(n_3222),
.Y(n_3287)
);

INVx1_ASAP7_75t_SL g3288 ( 
.A(n_3206),
.Y(n_3288)
);

OAI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3239),
.A2(n_413),
.B(n_416),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3181),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_3163),
.A2(n_425),
.B(n_427),
.Y(n_3291)
);

AO31x2_ASAP7_75t_L g3292 ( 
.A1(n_3182),
.A2(n_430),
.A3(n_3194),
.B(n_3196),
.Y(n_3292)
);

CKINVDCx20_ASAP7_75t_R g3293 ( 
.A(n_3203),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3154),
.A2(n_3146),
.B(n_3187),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3216),
.B(n_3185),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3232),
.B(n_3215),
.Y(n_3296)
);

OAI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3187),
.A2(n_3218),
.B(n_3146),
.Y(n_3297)
);

INVx2_ASAP7_75t_SL g3298 ( 
.A(n_3144),
.Y(n_3298)
);

OA21x2_ASAP7_75t_L g3299 ( 
.A1(n_3232),
.A2(n_3172),
.B(n_3166),
.Y(n_3299)
);

AOI21xp33_ASAP7_75t_SL g3300 ( 
.A1(n_3215),
.A2(n_3182),
.B(n_3165),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_3197),
.B(n_3234),
.Y(n_3301)
);

A2O1A1Ixp33_ASAP7_75t_L g3302 ( 
.A1(n_3214),
.A2(n_3230),
.B(n_3218),
.C(n_3193),
.Y(n_3302)
);

CKINVDCx14_ASAP7_75t_R g3303 ( 
.A(n_3162),
.Y(n_3303)
);

CKINVDCx20_ASAP7_75t_R g3304 ( 
.A(n_3184),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3192),
.Y(n_3305)
);

AND2x4_ASAP7_75t_L g3306 ( 
.A(n_3197),
.B(n_3221),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3167),
.B(n_3227),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3188),
.A2(n_3230),
.B(n_3229),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3165),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3209),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3167),
.B(n_3205),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3188),
.A2(n_3229),
.B(n_3220),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3205),
.B(n_3195),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3231),
.A2(n_3170),
.B(n_3191),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3205),
.B(n_3195),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3197),
.B(n_3221),
.Y(n_3316)
);

OAI21xp33_ASAP7_75t_SL g3317 ( 
.A1(n_3161),
.A2(n_3235),
.B(n_3164),
.Y(n_3317)
);

AO31x2_ASAP7_75t_L g3318 ( 
.A1(n_3240),
.A2(n_3191),
.A3(n_3224),
.B(n_3206),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3162),
.B(n_3199),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_3156),
.B(n_3174),
.Y(n_3320)
);

BUFx12f_ASAP7_75t_L g3321 ( 
.A(n_3223),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3160),
.B(n_3171),
.Y(n_3322)
);

HB1xp67_ASAP7_75t_L g3323 ( 
.A(n_3200),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3147),
.B(n_3222),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3147),
.B(n_3240),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3225),
.B(n_3219),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3294),
.B(n_3225),
.Y(n_3327)
);

OAI22xp5_ASAP7_75t_L g3328 ( 
.A1(n_3294),
.A2(n_3217),
.B1(n_3190),
.B2(n_3211),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_SL g3329 ( 
.A1(n_3297),
.A2(n_3236),
.B1(n_3238),
.B2(n_3225),
.Y(n_3329)
);

CKINVDCx20_ASAP7_75t_R g3330 ( 
.A(n_3249),
.Y(n_3330)
);

INVx4_ASAP7_75t_L g3331 ( 
.A(n_3253),
.Y(n_3331)
);

OAI22x1_ASAP7_75t_L g3332 ( 
.A1(n_3288),
.A2(n_3238),
.B1(n_3236),
.B2(n_3150),
.Y(n_3332)
);

BUFx4f_ASAP7_75t_SL g3333 ( 
.A(n_3304),
.Y(n_3333)
);

OAI21xp33_ASAP7_75t_L g3334 ( 
.A1(n_3269),
.A2(n_3150),
.B(n_3223),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3282),
.A2(n_3223),
.B1(n_3219),
.B2(n_3225),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_SL g3336 ( 
.A1(n_3322),
.A2(n_3219),
.B1(n_3241),
.B2(n_3326),
.Y(n_3336)
);

CKINVDCx5p33_ASAP7_75t_R g3337 ( 
.A(n_3242),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3312),
.A2(n_3308),
.B1(n_3289),
.B2(n_3248),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3269),
.A2(n_3312),
.B1(n_3308),
.B2(n_3288),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3254),
.Y(n_3340)
);

INVx6_ASAP7_75t_L g3341 ( 
.A(n_3287),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3314),
.B(n_3243),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3314),
.A2(n_3319),
.B(n_3289),
.Y(n_3343)
);

AOI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_3251),
.A2(n_3302),
.B1(n_3325),
.B2(n_3277),
.Y(n_3344)
);

OAI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3252),
.A2(n_3279),
.B1(n_3324),
.B2(n_3255),
.Y(n_3345)
);

BUFx4f_ASAP7_75t_SL g3346 ( 
.A(n_3286),
.Y(n_3346)
);

OAI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3255),
.A2(n_3311),
.B1(n_3321),
.B2(n_3252),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_3279),
.A2(n_3319),
.B1(n_3257),
.B2(n_3261),
.Y(n_3348)
);

NAND2x1_ASAP7_75t_L g3349 ( 
.A(n_3265),
.B(n_3299),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3257),
.A2(n_3261),
.B1(n_3291),
.B2(n_3303),
.Y(n_3350)
);

OAI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3281),
.A2(n_3291),
.B1(n_3244),
.B2(n_3247),
.Y(n_3351)
);

AND2x4_ASAP7_75t_L g3352 ( 
.A(n_3298),
.B(n_3301),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3313),
.A2(n_3315),
.B1(n_3256),
.B2(n_3244),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_3317),
.B(n_3300),
.Y(n_3354)
);

NAND3xp33_ASAP7_75t_L g3355 ( 
.A(n_3268),
.B(n_3275),
.C(n_3307),
.Y(n_3355)
);

BUFx3_ASAP7_75t_L g3356 ( 
.A(n_3272),
.Y(n_3356)
);

BUFx4f_ASAP7_75t_SL g3357 ( 
.A(n_3293),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3296),
.A2(n_3263),
.B1(n_3245),
.B2(n_3309),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_SL g3359 ( 
.A1(n_3258),
.A2(n_3262),
.B1(n_3267),
.B2(n_3270),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3306),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3296),
.A2(n_3301),
.B1(n_3307),
.B2(n_3262),
.Y(n_3361)
);

BUFx12f_ASAP7_75t_L g3362 ( 
.A(n_3264),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_3280),
.A2(n_3290),
.B1(n_3305),
.B2(n_3310),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_3266),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_3273),
.A2(n_3295),
.B1(n_3271),
.B2(n_3306),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3273),
.A2(n_3295),
.B1(n_3271),
.B2(n_3259),
.Y(n_3366)
);

OAI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_3318),
.A2(n_3323),
.B1(n_3250),
.B2(n_3320),
.Y(n_3367)
);

CKINVDCx5p33_ASAP7_75t_R g3368 ( 
.A(n_3287),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3246),
.Y(n_3369)
);

INVx4_ASAP7_75t_SL g3370 ( 
.A(n_3318),
.Y(n_3370)
);

NOR2xp67_ASAP7_75t_SL g3371 ( 
.A(n_3284),
.B(n_3299),
.Y(n_3371)
);

BUFx4f_ASAP7_75t_SL g3372 ( 
.A(n_3260),
.Y(n_3372)
);

OAI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_3318),
.A2(n_3250),
.B1(n_3243),
.B2(n_3292),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3274),
.A2(n_3243),
.B1(n_3278),
.B2(n_3285),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3294),
.A2(n_3269),
.B1(n_3312),
.B2(n_3326),
.Y(n_3376)
);

OAI222xp33_ASAP7_75t_L g3377 ( 
.A1(n_3294),
.A2(n_3322),
.B1(n_3326),
.B2(n_3269),
.C1(n_3308),
.C2(n_3148),
.Y(n_3377)
);

INVx4_ASAP7_75t_L g3378 ( 
.A(n_3253),
.Y(n_3378)
);

CKINVDCx5p33_ASAP7_75t_R g3379 ( 
.A(n_3249),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_SL g3381 ( 
.A1(n_3297),
.A2(n_3294),
.B1(n_3322),
.B2(n_3326),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3316),
.B(n_3265),
.Y(n_3382)
);

BUFx12f_ASAP7_75t_L g3383 ( 
.A(n_3242),
.Y(n_3383)
);

OR2x2_ASAP7_75t_L g3384 ( 
.A(n_3276),
.B(n_3270),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3385)
);

INVx3_ASAP7_75t_L g3386 ( 
.A(n_3265),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3294),
.A2(n_3269),
.B1(n_3312),
.B2(n_3326),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3294),
.A2(n_3269),
.B1(n_3312),
.B2(n_3326),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3254),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_SL g3392 ( 
.A1(n_3297),
.A2(n_3294),
.B1(n_3322),
.B2(n_3326),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3254),
.Y(n_3393)
);

INVx5_ASAP7_75t_SL g3394 ( 
.A(n_3253),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3297),
.A2(n_3294),
.B(n_3308),
.Y(n_3396)
);

AOI22xp5_ASAP7_75t_SL g3397 ( 
.A1(n_3288),
.A2(n_3325),
.B1(n_3286),
.B2(n_3303),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3399)
);

AND2x4_ASAP7_75t_L g3400 ( 
.A(n_3265),
.B(n_3298),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3401)
);

AOI22xp33_ASAP7_75t_L g3402 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3402)
);

BUFx6f_ASAP7_75t_L g3403 ( 
.A(n_3253),
.Y(n_3403)
);

BUFx4f_ASAP7_75t_L g3404 ( 
.A(n_3253),
.Y(n_3404)
);

AOI22xp33_ASAP7_75t_L g3405 ( 
.A1(n_3297),
.A2(n_3282),
.B1(n_3294),
.B2(n_3283),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3294),
.B(n_3179),
.Y(n_3406)
);

OAI21xp5_ASAP7_75t_SL g3407 ( 
.A1(n_3269),
.A2(n_3153),
.B(n_3251),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_SL g3408 ( 
.A1(n_3297),
.A2(n_3294),
.B1(n_3322),
.B2(n_3326),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3396),
.B(n_3407),
.Y(n_3409)
);

AO21x2_ASAP7_75t_L g3410 ( 
.A1(n_3342),
.A2(n_3347),
.B(n_3338),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_3349),
.Y(n_3411)
);

OR2x2_ASAP7_75t_L g3412 ( 
.A(n_3384),
.B(n_3327),
.Y(n_3412)
);

AO21x2_ASAP7_75t_L g3413 ( 
.A1(n_3347),
.A2(n_3406),
.B(n_3367),
.Y(n_3413)
);

HB1xp67_ASAP7_75t_L g3414 ( 
.A(n_3332),
.Y(n_3414)
);

AO21x2_ASAP7_75t_L g3415 ( 
.A1(n_3367),
.A2(n_3373),
.B(n_3377),
.Y(n_3415)
);

AO221x2_ASAP7_75t_L g3416 ( 
.A1(n_3339),
.A2(n_3377),
.B1(n_3345),
.B2(n_3389),
.C(n_3376),
.Y(n_3416)
);

INVx3_ASAP7_75t_L g3417 ( 
.A(n_3341),
.Y(n_3417)
);

OR2x2_ASAP7_75t_L g3418 ( 
.A(n_3390),
.B(n_3369),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3382),
.B(n_3360),
.Y(n_3419)
);

OR2x6_ASAP7_75t_L g3420 ( 
.A(n_3343),
.B(n_3341),
.Y(n_3420)
);

OR2x6_ASAP7_75t_L g3421 ( 
.A(n_3341),
.B(n_3350),
.Y(n_3421)
);

AO31x2_ASAP7_75t_L g3422 ( 
.A1(n_3358),
.A2(n_3348),
.A3(n_3393),
.B(n_3391),
.Y(n_3422)
);

OA21x2_ASAP7_75t_L g3423 ( 
.A1(n_3375),
.A2(n_3398),
.B(n_3405),
.Y(n_3423)
);

AO21x2_ASAP7_75t_L g3424 ( 
.A1(n_3373),
.A2(n_3344),
.B(n_3340),
.Y(n_3424)
);

BUFx3_ASAP7_75t_L g3425 ( 
.A(n_3346),
.Y(n_3425)
);

BUFx3_ASAP7_75t_L g3426 ( 
.A(n_3346),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3328),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3355),
.Y(n_3428)
);

AO21x2_ASAP7_75t_L g3429 ( 
.A1(n_3361),
.A2(n_3354),
.B(n_3351),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3386),
.B(n_3371),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3352),
.B(n_3397),
.Y(n_3431)
);

INVxp67_ASAP7_75t_R g3432 ( 
.A(n_3394),
.Y(n_3432)
);

OA21x2_ASAP7_75t_L g3433 ( 
.A1(n_3380),
.A2(n_3395),
.B(n_3385),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3329),
.Y(n_3434)
);

BUFx2_ASAP7_75t_L g3435 ( 
.A(n_3372),
.Y(n_3435)
);

AO21x2_ASAP7_75t_L g3436 ( 
.A1(n_3351),
.A2(n_3334),
.B(n_3370),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3352),
.B(n_3366),
.Y(n_3437)
);

OR2x6_ASAP7_75t_L g3438 ( 
.A(n_3356),
.B(n_3403),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_3357),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_SL g3440 ( 
.A1(n_3368),
.A2(n_3370),
.B(n_3331),
.Y(n_3440)
);

OA21x2_ASAP7_75t_L g3441 ( 
.A1(n_3387),
.A2(n_3402),
.B(n_3401),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3381),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3365),
.B(n_3394),
.Y(n_3443)
);

BUFx2_ASAP7_75t_L g3444 ( 
.A(n_3372),
.Y(n_3444)
);

HB1xp67_ASAP7_75t_L g3445 ( 
.A(n_3362),
.Y(n_3445)
);

INVxp67_ASAP7_75t_L g3446 ( 
.A(n_3403),
.Y(n_3446)
);

BUFx12f_ASAP7_75t_L g3447 ( 
.A(n_3403),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3333),
.Y(n_3448)
);

INVx2_ASAP7_75t_SL g3449 ( 
.A(n_3404),
.Y(n_3449)
);

AOI221xp5_ASAP7_75t_L g3450 ( 
.A1(n_3381),
.A2(n_3392),
.B1(n_3408),
.B2(n_3399),
.C(n_3388),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3333),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3357),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3394),
.B(n_3353),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3392),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_3404),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3408),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3336),
.Y(n_3457)
);

OR2x2_ASAP7_75t_L g3458 ( 
.A(n_3359),
.B(n_3374),
.Y(n_3458)
);

OR2x6_ASAP7_75t_L g3459 ( 
.A(n_3331),
.B(n_3378),
.Y(n_3459)
);

INVx4_ASAP7_75t_L g3460 ( 
.A(n_3378),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3330),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3379),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3364),
.Y(n_3463)
);

AO21x2_ASAP7_75t_L g3464 ( 
.A1(n_3336),
.A2(n_3335),
.B(n_3363),
.Y(n_3464)
);

BUFx3_ASAP7_75t_L g3465 ( 
.A(n_3383),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3337),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_3346),
.Y(n_3467)
);

HB1xp67_ASAP7_75t_L g3468 ( 
.A(n_3332),
.Y(n_3468)
);

HB1xp67_ASAP7_75t_L g3469 ( 
.A(n_3332),
.Y(n_3469)
);

OA21x2_ASAP7_75t_L g3470 ( 
.A1(n_3407),
.A2(n_3396),
.B(n_3377),
.Y(n_3470)
);

AOI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3396),
.A2(n_3343),
.B(n_3327),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3396),
.B(n_3407),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3382),
.B(n_3360),
.Y(n_3473)
);

AND2x4_ASAP7_75t_L g3474 ( 
.A(n_3400),
.B(n_3338),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3429),
.B(n_3471),
.Y(n_3475)
);

BUFx2_ASAP7_75t_L g3476 ( 
.A(n_3470),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3429),
.B(n_3471),
.Y(n_3477)
);

HB1xp67_ASAP7_75t_L g3478 ( 
.A(n_3470),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3415),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3429),
.B(n_3470),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3415),
.Y(n_3481)
);

OR2x2_ASAP7_75t_L g3482 ( 
.A(n_3434),
.B(n_3428),
.Y(n_3482)
);

HB1xp67_ASAP7_75t_L g3483 ( 
.A(n_3470),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3434),
.Y(n_3484)
);

INVxp67_ASAP7_75t_L g3485 ( 
.A(n_3425),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3415),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3416),
.B(n_3431),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3464),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3442),
.B(n_3454),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3416),
.B(n_3431),
.Y(n_3490)
);

BUFx2_ASAP7_75t_L g3491 ( 
.A(n_3438),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3416),
.B(n_3443),
.Y(n_3492)
);

NAND2x1_ASAP7_75t_L g3493 ( 
.A(n_3411),
.B(n_3421),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3416),
.B(n_3443),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3419),
.B(n_3473),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3419),
.B(n_3473),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3414),
.B(n_3468),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3469),
.B(n_3422),
.Y(n_3498)
);

BUFx3_ASAP7_75t_L g3499 ( 
.A(n_3425),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3464),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3464),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3442),
.B(n_3454),
.Y(n_3502)
);

BUFx3_ASAP7_75t_L g3503 ( 
.A(n_3426),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3436),
.B(n_3411),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3437),
.B(n_3430),
.Y(n_3505)
);

OAI33xp33_ASAP7_75t_L g3506 ( 
.A1(n_3456),
.A2(n_3457),
.A3(n_3458),
.B1(n_3472),
.B2(n_3409),
.B3(n_3427),
.Y(n_3506)
);

AOI22xp5_ASAP7_75t_L g3507 ( 
.A1(n_3450),
.A2(n_3456),
.B1(n_3457),
.B2(n_3441),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3437),
.B(n_3430),
.Y(n_3508)
);

OR2x2_ASAP7_75t_SL g3509 ( 
.A(n_3423),
.B(n_3433),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3423),
.B(n_3433),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3453),
.B(n_3435),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3435),
.B(n_3444),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_3426),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3423),
.B(n_3433),
.Y(n_3514)
);

BUFx3_ASAP7_75t_L g3515 ( 
.A(n_3467),
.Y(n_3515)
);

AO21x2_ASAP7_75t_L g3516 ( 
.A1(n_3424),
.A2(n_3413),
.B(n_3436),
.Y(n_3516)
);

INVx1_ASAP7_75t_SL g3517 ( 
.A(n_3467),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3444),
.B(n_3420),
.Y(n_3518)
);

BUFx2_ASAP7_75t_L g3519 ( 
.A(n_3438),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3420),
.B(n_3413),
.Y(n_3520)
);

HB1xp67_ASAP7_75t_L g3521 ( 
.A(n_3423),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3458),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3410),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3410),
.Y(n_3524)
);

INVx4_ASAP7_75t_L g3525 ( 
.A(n_3447),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3410),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3413),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3433),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3441),
.B(n_3427),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_3480),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_3480),
.B(n_3475),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3516),
.Y(n_3532)
);

HB1xp67_ASAP7_75t_L g3533 ( 
.A(n_3480),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3476),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3476),
.Y(n_3535)
);

HB1xp67_ASAP7_75t_L g3536 ( 
.A(n_3475),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3475),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3516),
.Y(n_3538)
);

HB1xp67_ASAP7_75t_L g3539 ( 
.A(n_3477),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3478),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3478),
.Y(n_3541)
);

INVx3_ASAP7_75t_L g3542 ( 
.A(n_3477),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3477),
.B(n_3483),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3516),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3483),
.B(n_3420),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_3520),
.Y(n_3546)
);

INVx5_ASAP7_75t_SL g3547 ( 
.A(n_3513),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3516),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3487),
.B(n_3420),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3521),
.Y(n_3550)
);

INVx2_ASAP7_75t_SL g3551 ( 
.A(n_3520),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3487),
.B(n_3421),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3521),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3520),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3487),
.B(n_3421),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3498),
.Y(n_3556)
);

INVx1_ASAP7_75t_SL g3557 ( 
.A(n_3527),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3490),
.B(n_3421),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_3504),
.B(n_3417),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3479),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3479),
.Y(n_3561)
);

INVx3_ASAP7_75t_L g3562 ( 
.A(n_3504),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3509),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3509),
.Y(n_3564)
);

INVx3_ASAP7_75t_L g3565 ( 
.A(n_3504),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3490),
.B(n_3441),
.Y(n_3566)
);

NAND2xp33_ASAP7_75t_SL g3567 ( 
.A(n_3490),
.B(n_3418),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3497),
.B(n_3441),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3479),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3527),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3481),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3492),
.B(n_3412),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3527),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3497),
.B(n_3418),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3481),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3497),
.B(n_3492),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3481),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3486),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3486),
.Y(n_3579)
);

AND2x2_ASAP7_75t_L g3580 ( 
.A(n_3492),
.B(n_3494),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3494),
.B(n_3474),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3486),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3523),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3580),
.B(n_3494),
.Y(n_3584)
);

HB1xp67_ASAP7_75t_L g3585 ( 
.A(n_3530),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3580),
.B(n_3576),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3580),
.A2(n_3507),
.B1(n_3474),
.B2(n_3493),
.Y(n_3587)
);

NAND3xp33_ASAP7_75t_L g3588 ( 
.A(n_3533),
.B(n_3507),
.C(n_3510),
.Y(n_3588)
);

INVx4_ASAP7_75t_L g3589 ( 
.A(n_3542),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3530),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3580),
.B(n_3505),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3566),
.B(n_3488),
.Y(n_3592)
);

OR2x2_ASAP7_75t_L g3593 ( 
.A(n_3533),
.B(n_3482),
.Y(n_3593)
);

AND2x2_ASAP7_75t_L g3594 ( 
.A(n_3576),
.B(n_3505),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3530),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3576),
.B(n_3505),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3530),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3566),
.B(n_3488),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3566),
.B(n_3488),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3576),
.B(n_3508),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3566),
.B(n_3500),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3531),
.B(n_3500),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3543),
.B(n_3508),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3531),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3543),
.B(n_3508),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3563),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3543),
.B(n_3495),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3563),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3563),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3563),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3543),
.B(n_3495),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3564),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3574),
.B(n_3495),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3574),
.B(n_3496),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3531),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3531),
.Y(n_3616)
);

BUFx3_ASAP7_75t_L g3617 ( 
.A(n_3531),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3564),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3574),
.B(n_3552),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3574),
.B(n_3496),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3531),
.B(n_3500),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3552),
.B(n_3496),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3564),
.B(n_3546),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3552),
.B(n_3499),
.Y(n_3624)
);

AND2x2_ASAP7_75t_L g3625 ( 
.A(n_3552),
.B(n_3499),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3564),
.Y(n_3626)
);

NOR3xp33_ASAP7_75t_L g3627 ( 
.A(n_3542),
.B(n_3506),
.C(n_3510),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3536),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3536),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3555),
.B(n_3499),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3537),
.Y(n_3631)
);

AND2x4_ASAP7_75t_SL g3632 ( 
.A(n_3559),
.B(n_3438),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3568),
.B(n_3501),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3555),
.B(n_3503),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3542),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3585),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3585),
.Y(n_3637)
);

BUFx3_ASAP7_75t_L g3638 ( 
.A(n_3623),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3626),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3591),
.B(n_3432),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3627),
.B(n_3568),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3626),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3591),
.B(n_3555),
.Y(n_3643)
);

AND2x2_ASAP7_75t_L g3644 ( 
.A(n_3591),
.B(n_3555),
.Y(n_3644)
);

HB1xp67_ASAP7_75t_L g3645 ( 
.A(n_3593),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3613),
.B(n_3558),
.Y(n_3646)
);

OR2x2_ASAP7_75t_L g3647 ( 
.A(n_3593),
.B(n_3537),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3593),
.B(n_3539),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3613),
.B(n_3432),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3613),
.B(n_3614),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3614),
.B(n_3549),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3623),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3614),
.B(n_3549),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3626),
.Y(n_3654)
);

OR2x2_ASAP7_75t_L g3655 ( 
.A(n_3627),
.B(n_3539),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3620),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3588),
.B(n_3542),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3620),
.B(n_3549),
.Y(n_3658)
);

INVx3_ASAP7_75t_L g3659 ( 
.A(n_3623),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3623),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3620),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3584),
.B(n_3568),
.Y(n_3662)
);

OR2x2_ASAP7_75t_L g3663 ( 
.A(n_3588),
.B(n_3542),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_3619),
.B(n_3549),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3584),
.B(n_3568),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3619),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3619),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3594),
.B(n_3558),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3594),
.B(n_3558),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3594),
.B(n_3596),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3584),
.B(n_3542),
.Y(n_3671)
);

AND2x4_ASAP7_75t_SL g3672 ( 
.A(n_3624),
.B(n_3438),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3633),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3633),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3643),
.Y(n_3675)
);

HB1xp67_ASAP7_75t_L g3676 ( 
.A(n_3657),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3650),
.B(n_3596),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_3641),
.B(n_3506),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3662),
.B(n_3586),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3650),
.B(n_3596),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3643),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3646),
.B(n_3624),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3662),
.B(n_3586),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3643),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3646),
.B(n_3624),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3644),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3670),
.B(n_3600),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3646),
.B(n_3625),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3670),
.B(n_3600),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3641),
.B(n_3525),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3644),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3644),
.B(n_3600),
.Y(n_3692)
);

NAND2x1p5_ASAP7_75t_L g3693 ( 
.A(n_3638),
.B(n_3525),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_3672),
.B(n_3525),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3668),
.B(n_3625),
.Y(n_3695)
);

AND2x4_ASAP7_75t_L g3696 ( 
.A(n_3638),
.B(n_3503),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3652),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3652),
.Y(n_3698)
);

INVx3_ASAP7_75t_L g3699 ( 
.A(n_3657),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3668),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3680),
.B(n_3586),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_3696),
.B(n_3525),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3680),
.B(n_3622),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3676),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3692),
.B(n_3622),
.Y(n_3705)
);

OR2x2_ASAP7_75t_L g3706 ( 
.A(n_3682),
.B(n_3665),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3677),
.B(n_3622),
.Y(n_3707)
);

AOI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3678),
.A2(n_3567),
.B1(n_3522),
.B2(n_3592),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3696),
.B(n_3513),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3687),
.B(n_3669),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_3685),
.B(n_3665),
.Y(n_3711)
);

OR2x2_ASAP7_75t_L g3712 ( 
.A(n_3688),
.B(n_3666),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3696),
.Y(n_3713)
);

OR2x2_ASAP7_75t_L g3714 ( 
.A(n_3695),
.B(n_3666),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3689),
.B(n_3669),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3678),
.B(n_3603),
.Y(n_3716)
);

OR2x2_ASAP7_75t_L g3717 ( 
.A(n_3679),
.B(n_3667),
.Y(n_3717)
);

NAND2x1_ASAP7_75t_L g3718 ( 
.A(n_3697),
.B(n_3440),
.Y(n_3718)
);

AND2x4_ASAP7_75t_SL g3719 ( 
.A(n_3694),
.B(n_3452),
.Y(n_3719)
);

OR2x2_ASAP7_75t_L g3720 ( 
.A(n_3683),
.B(n_3667),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3701),
.B(n_3625),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3703),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3705),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3707),
.B(n_3630),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3710),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3715),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3708),
.B(n_3603),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3708),
.B(n_3603),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3717),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3713),
.B(n_3630),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3719),
.B(n_3630),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_L g3732 ( 
.A(n_3718),
.B(n_3672),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3706),
.B(n_3634),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3711),
.B(n_3672),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3720),
.Y(n_3735)
);

INVx3_ASAP7_75t_L g3736 ( 
.A(n_3712),
.Y(n_3736)
);

INVxp67_ASAP7_75t_L g3737 ( 
.A(n_3709),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3721),
.Y(n_3738)
);

OAI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3730),
.A2(n_3663),
.B1(n_3655),
.B2(n_3572),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3724),
.Y(n_3740)
);

AOI322xp5_ASAP7_75t_L g3741 ( 
.A1(n_3727),
.A2(n_3514),
.A3(n_3567),
.B1(n_3522),
.B2(n_3528),
.C1(n_3501),
.C2(n_3598),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3733),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3736),
.B(n_3634),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3736),
.B(n_3634),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3727),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3731),
.B(n_3503),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_SL g3747 ( 
.A(n_3729),
.B(n_3513),
.Y(n_3747)
);

OR2x2_ASAP7_75t_L g3748 ( 
.A(n_3728),
.B(n_3605),
.Y(n_3748)
);

HB1xp67_ASAP7_75t_L g3749 ( 
.A(n_3725),
.Y(n_3749)
);

NAND2xp33_ASAP7_75t_SL g3750 ( 
.A(n_3743),
.B(n_3513),
.Y(n_3750)
);

OAI22xp33_ASAP7_75t_SL g3751 ( 
.A1(n_3744),
.A2(n_3655),
.B1(n_3663),
.B2(n_3514),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3748),
.B(n_3605),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3749),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3746),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3746),
.Y(n_3755)
);

AOI222xp33_ASAP7_75t_L g3756 ( 
.A1(n_3739),
.A2(n_3501),
.B1(n_3546),
.B2(n_3524),
.C1(n_3523),
.C2(n_3526),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3740),
.B(n_3605),
.Y(n_3757)
);

OAI22xp33_ASAP7_75t_L g3758 ( 
.A1(n_3753),
.A2(n_3676),
.B1(n_3716),
.B2(n_3598),
.Y(n_3758)
);

AND2x2_ASAP7_75t_SL g3759 ( 
.A(n_3757),
.B(n_3735),
.Y(n_3759)
);

XOR2x2_ASAP7_75t_L g3760 ( 
.A(n_3751),
.B(n_3716),
.Y(n_3760)
);

INVxp67_ASAP7_75t_L g3761 ( 
.A(n_3752),
.Y(n_3761)
);

AOI211xp5_ASAP7_75t_SL g3762 ( 
.A1(n_3753),
.A2(n_3745),
.B(n_3738),
.C(n_3704),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3754),
.Y(n_3763)
);

AOI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3756),
.A2(n_3599),
.B1(n_3601),
.B2(n_3592),
.Y(n_3764)
);

AOI211xp5_ASAP7_75t_L g3765 ( 
.A1(n_3750),
.A2(n_3690),
.B(n_3728),
.C(n_3732),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3755),
.A2(n_3601),
.B1(n_3599),
.B2(n_3550),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3757),
.B(n_3558),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3752),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3757),
.B(n_3664),
.Y(n_3769)
);

OAI211xp5_ASAP7_75t_SL g3770 ( 
.A1(n_3753),
.A2(n_3741),
.B(n_3737),
.C(n_3747),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3767),
.A2(n_3699),
.B(n_3704),
.Y(n_3771)
);

A2O1A1Ixp33_ASAP7_75t_L g3772 ( 
.A1(n_3764),
.A2(n_3553),
.B(n_3550),
.C(n_3699),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3769),
.B(n_3664),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3759),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3758),
.B(n_3651),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3766),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3768),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3762),
.B(n_3651),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3760),
.B(n_3653),
.Y(n_3779)
);

OAI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3761),
.A2(n_3690),
.B(n_3660),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3763),
.Y(n_3781)
);

AOI221xp5_ASAP7_75t_SL g3782 ( 
.A1(n_3765),
.A2(n_3698),
.B1(n_3675),
.B2(n_3681),
.C(n_3684),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3770),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3769),
.Y(n_3784)
);

OAI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_3767),
.A2(n_3671),
.B1(n_3616),
.B2(n_3604),
.Y(n_3785)
);

O2A1O1Ixp33_ASAP7_75t_L g3786 ( 
.A1(n_3758),
.A2(n_3699),
.B(n_3645),
.C(n_3553),
.Y(n_3786)
);

OR2x2_ASAP7_75t_L g3787 ( 
.A(n_3767),
.B(n_3671),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3769),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3769),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3769),
.Y(n_3790)
);

AOI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3764),
.A2(n_3553),
.B1(n_3550),
.B2(n_3606),
.Y(n_3791)
);

AOI322xp5_ASAP7_75t_L g3792 ( 
.A1(n_3758),
.A2(n_3522),
.A3(n_3528),
.B1(n_3606),
.B2(n_3609),
.C1(n_3608),
.C2(n_3610),
.Y(n_3792)
);

OAI21xp33_ASAP7_75t_L g3793 ( 
.A1(n_3773),
.A2(n_3700),
.B(n_3691),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3784),
.B(n_3638),
.Y(n_3794)
);

AOI221xp5_ASAP7_75t_L g3795 ( 
.A1(n_3783),
.A2(n_3535),
.B1(n_3534),
.B2(n_3541),
.C(n_3540),
.Y(n_3795)
);

AOI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3774),
.A2(n_3623),
.B1(n_3609),
.B2(n_3610),
.Y(n_3796)
);

INVxp67_ASAP7_75t_L g3797 ( 
.A(n_3778),
.Y(n_3797)
);

HB1xp67_ASAP7_75t_L g3798 ( 
.A(n_3777),
.Y(n_3798)
);

OAI21xp33_ASAP7_75t_L g3799 ( 
.A1(n_3779),
.A2(n_3686),
.B(n_3734),
.Y(n_3799)
);

AOI221xp5_ASAP7_75t_SL g3800 ( 
.A1(n_3771),
.A2(n_3786),
.B1(n_3785),
.B2(n_3780),
.C(n_3636),
.Y(n_3800)
);

NOR4xp25_ASAP7_75t_L g3801 ( 
.A(n_3772),
.B(n_3775),
.C(n_3781),
.D(n_3776),
.Y(n_3801)
);

AOI221xp5_ASAP7_75t_L g3802 ( 
.A1(n_3788),
.A2(n_3535),
.B1(n_3534),
.B2(n_3541),
.C(n_3540),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3790),
.A2(n_3645),
.B(n_3660),
.Y(n_3803)
);

AOI221xp5_ASAP7_75t_L g3804 ( 
.A1(n_3791),
.A2(n_3535),
.B1(n_3534),
.B2(n_3541),
.C(n_3540),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3792),
.B(n_3659),
.Y(n_3805)
);

NAND3xp33_ASAP7_75t_L g3806 ( 
.A(n_3789),
.B(n_3742),
.C(n_3660),
.Y(n_3806)
);

NAND3xp33_ASAP7_75t_SL g3807 ( 
.A(n_3787),
.B(n_3693),
.C(n_3648),
.Y(n_3807)
);

INVxp33_ASAP7_75t_L g3808 ( 
.A(n_3782),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3791),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3784),
.Y(n_3810)
);

OAI21xp5_ASAP7_75t_SL g3811 ( 
.A1(n_3778),
.A2(n_3694),
.B(n_3693),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3784),
.Y(n_3812)
);

OAI21xp33_ASAP7_75t_L g3813 ( 
.A1(n_3773),
.A2(n_3726),
.B(n_3722),
.Y(n_3813)
);

NAND4xp25_ASAP7_75t_L g3814 ( 
.A(n_3782),
.B(n_3702),
.C(n_3723),
.D(n_3714),
.Y(n_3814)
);

AOI221xp5_ASAP7_75t_L g3815 ( 
.A1(n_3783),
.A2(n_3618),
.B1(n_3608),
.B2(n_3612),
.C(n_3674),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3784),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3778),
.A2(n_3659),
.B(n_3637),
.Y(n_3817)
);

INVx1_ASAP7_75t_SL g3818 ( 
.A(n_3773),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3810),
.A2(n_3595),
.B1(n_3590),
.B2(n_3674),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3796),
.B(n_3659),
.Y(n_3820)
);

OAI211xp5_ASAP7_75t_L g3821 ( 
.A1(n_3811),
.A2(n_3659),
.B(n_3636),
.C(n_3637),
.Y(n_3821)
);

OAI21xp33_ASAP7_75t_L g3822 ( 
.A1(n_3812),
.A2(n_3649),
.B(n_3640),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3816),
.A2(n_3528),
.B1(n_3546),
.B2(n_3524),
.Y(n_3823)
);

NAND4xp25_ASAP7_75t_L g3824 ( 
.A(n_3794),
.B(n_3529),
.C(n_3649),
.D(n_3502),
.Y(n_3824)
);

NOR3x1_ASAP7_75t_L g3825 ( 
.A(n_3806),
.B(n_3807),
.C(n_3814),
.Y(n_3825)
);

OAI211xp5_ASAP7_75t_SL g3826 ( 
.A1(n_3797),
.A2(n_3602),
.B(n_3621),
.C(n_3597),
.Y(n_3826)
);

AOI221xp5_ASAP7_75t_L g3827 ( 
.A1(n_3801),
.A2(n_3612),
.B1(n_3618),
.B2(n_3590),
.C(n_3595),
.Y(n_3827)
);

AOI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3818),
.A2(n_3595),
.B1(n_3590),
.B2(n_3673),
.Y(n_3828)
);

AOI31xp33_ASAP7_75t_L g3829 ( 
.A1(n_3808),
.A2(n_3517),
.A3(n_3485),
.B(n_3656),
.Y(n_3829)
);

OAI22xp5_ASAP7_75t_L g3830 ( 
.A1(n_3803),
.A2(n_3616),
.B1(n_3604),
.B2(n_3617),
.Y(n_3830)
);

NOR3xp33_ASAP7_75t_L g3831 ( 
.A(n_3798),
.B(n_3813),
.C(n_3799),
.Y(n_3831)
);

AOI322xp5_ASAP7_75t_L g3832 ( 
.A1(n_3815),
.A2(n_3673),
.A3(n_3621),
.B1(n_3602),
.B2(n_3642),
.C1(n_3551),
.C2(n_3654),
.Y(n_3832)
);

OAI21xp33_ASAP7_75t_L g3833 ( 
.A1(n_3793),
.A2(n_3640),
.B(n_3661),
.Y(n_3833)
);

OAI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_3805),
.A2(n_3604),
.B1(n_3616),
.B2(n_3617),
.Y(n_3834)
);

AOI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_3809),
.A2(n_3597),
.B1(n_3545),
.B2(n_3615),
.Y(n_3835)
);

OAI221xp5_ASAP7_75t_SL g3836 ( 
.A1(n_3817),
.A2(n_3647),
.B1(n_3648),
.B2(n_3656),
.C(n_3661),
.Y(n_3836)
);

OAI321xp33_ASAP7_75t_L g3837 ( 
.A1(n_3795),
.A2(n_3642),
.A3(n_3654),
.B1(n_3639),
.B2(n_3628),
.C(n_3631),
.Y(n_3837)
);

A2O1A1O1Ixp25_ASAP7_75t_L g3838 ( 
.A1(n_3800),
.A2(n_3631),
.B(n_3628),
.C(n_3629),
.D(n_3587),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3802),
.Y(n_3839)
);

OAI21xp5_ASAP7_75t_SL g3840 ( 
.A1(n_3804),
.A2(n_3632),
.B(n_3658),
.Y(n_3840)
);

OAI21xp5_ASAP7_75t_SL g3841 ( 
.A1(n_3811),
.A2(n_3632),
.B(n_3658),
.Y(n_3841)
);

OAI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3810),
.A2(n_3654),
.B(n_3639),
.Y(n_3842)
);

OAI221xp5_ASAP7_75t_L g3843 ( 
.A1(n_3841),
.A2(n_3647),
.B1(n_3617),
.B2(n_3629),
.C(n_3615),
.Y(n_3843)
);

OAI221xp5_ASAP7_75t_L g3844 ( 
.A1(n_3827),
.A2(n_3615),
.B1(n_3589),
.B2(n_3519),
.C(n_3491),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3824),
.A2(n_3615),
.B1(n_3635),
.B2(n_3545),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3823),
.B(n_3639),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3835),
.B(n_3653),
.Y(n_3847)
);

NAND2xp33_ASAP7_75t_L g3848 ( 
.A(n_3831),
.B(n_3513),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3832),
.B(n_3557),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_SL g3850 ( 
.A(n_3828),
.B(n_3513),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3837),
.A2(n_3635),
.B(n_3545),
.Y(n_3851)
);

AOI211xp5_ASAP7_75t_L g3852 ( 
.A1(n_3836),
.A2(n_3587),
.B(n_3545),
.C(n_3581),
.Y(n_3852)
);

AOI211xp5_ASAP7_75t_L g3853 ( 
.A1(n_3821),
.A2(n_3581),
.B(n_3635),
.C(n_3572),
.Y(n_3853)
);

OAI321xp33_ASAP7_75t_L g3854 ( 
.A1(n_3826),
.A2(n_3551),
.A3(n_3526),
.B1(n_3524),
.B2(n_3523),
.C(n_3554),
.Y(n_3854)
);

AOI221xp5_ASAP7_75t_L g3855 ( 
.A1(n_3830),
.A2(n_3551),
.B1(n_3546),
.B2(n_3557),
.C(n_3589),
.Y(n_3855)
);

OAI221xp5_ASAP7_75t_L g3856 ( 
.A1(n_3840),
.A2(n_3589),
.B1(n_3491),
.B2(n_3519),
.C(n_3551),
.Y(n_3856)
);

AOI22xp33_ASAP7_75t_L g3857 ( 
.A1(n_3834),
.A2(n_3554),
.B1(n_3526),
.B2(n_3565),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3820),
.A2(n_3589),
.B(n_3556),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3829),
.B(n_3517),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_SL g3860 ( 
.A(n_3859),
.B(n_3822),
.Y(n_3860)
);

INVxp33_ASAP7_75t_SL g3861 ( 
.A(n_3847),
.Y(n_3861)
);

NOR2x1_ASAP7_75t_L g3862 ( 
.A(n_3848),
.B(n_3842),
.Y(n_3862)
);

INVxp67_ASAP7_75t_L g3863 ( 
.A(n_3850),
.Y(n_3863)
);

AOI211xp5_ASAP7_75t_L g3864 ( 
.A1(n_3843),
.A2(n_3839),
.B(n_3833),
.C(n_3819),
.Y(n_3864)
);

NOR3xp33_ASAP7_75t_L g3865 ( 
.A(n_3849),
.B(n_3846),
.C(n_3854),
.Y(n_3865)
);

OAI211xp5_ASAP7_75t_L g3866 ( 
.A1(n_3858),
.A2(n_3838),
.B(n_3825),
.C(n_3589),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3855),
.A2(n_3562),
.B1(n_3565),
.B2(n_3554),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3845),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3844),
.Y(n_3869)
);

NOR2x1_ASAP7_75t_L g3870 ( 
.A(n_3851),
.B(n_3515),
.Y(n_3870)
);

NAND3xp33_ASAP7_75t_L g3871 ( 
.A(n_3853),
.B(n_3502),
.C(n_3489),
.Y(n_3871)
);

INVxp67_ASAP7_75t_SL g3872 ( 
.A(n_3857),
.Y(n_3872)
);

NAND3xp33_ASAP7_75t_SL g3873 ( 
.A(n_3852),
.B(n_3557),
.C(n_3489),
.Y(n_3873)
);

NOR2x1p5_ASAP7_75t_L g3874 ( 
.A(n_3856),
.B(n_3515),
.Y(n_3874)
);

NAND4xp25_ASAP7_75t_L g3875 ( 
.A(n_3864),
.B(n_3529),
.C(n_3515),
.D(n_3512),
.Y(n_3875)
);

O2A1O1Ixp33_ASAP7_75t_L g3876 ( 
.A1(n_3861),
.A2(n_3556),
.B(n_3581),
.C(n_3482),
.Y(n_3876)
);

AOI211x1_ASAP7_75t_L g3877 ( 
.A1(n_3866),
.A2(n_3611),
.B(n_3607),
.C(n_3581),
.Y(n_3877)
);

OAI211xp5_ASAP7_75t_SL g3878 ( 
.A1(n_3862),
.A2(n_3582),
.B(n_3560),
.C(n_3561),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3870),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_L g3880 ( 
.A(n_3873),
.B(n_3465),
.Y(n_3880)
);

NAND3xp33_ASAP7_75t_L g3881 ( 
.A(n_3865),
.B(n_3560),
.C(n_3561),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3874),
.B(n_3513),
.Y(n_3882)
);

OAI221xp5_ASAP7_75t_L g3883 ( 
.A1(n_3867),
.A2(n_3562),
.B1(n_3565),
.B2(n_3607),
.C(n_3611),
.Y(n_3883)
);

NOR2x1_ASAP7_75t_L g3884 ( 
.A(n_3868),
.B(n_3465),
.Y(n_3884)
);

NAND3xp33_ASAP7_75t_L g3885 ( 
.A(n_3860),
.B(n_3561),
.C(n_3560),
.Y(n_3885)
);

AOI22x1_ASAP7_75t_L g3886 ( 
.A1(n_3872),
.A2(n_3611),
.B1(n_3607),
.B2(n_3512),
.Y(n_3886)
);

NAND3xp33_ASAP7_75t_SL g3887 ( 
.A(n_3863),
.B(n_3578),
.C(n_3575),
.Y(n_3887)
);

OAI211xp5_ASAP7_75t_SL g3888 ( 
.A1(n_3869),
.A2(n_3575),
.B(n_3577),
.C(n_3582),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_SL g3889 ( 
.A(n_3871),
.B(n_3447),
.Y(n_3889)
);

NAND4xp25_ASAP7_75t_L g3890 ( 
.A(n_3864),
.B(n_3512),
.C(n_3485),
.D(n_3582),
.Y(n_3890)
);

AOI221xp5_ASAP7_75t_L g3891 ( 
.A1(n_3873),
.A2(n_3562),
.B1(n_3565),
.B2(n_3559),
.C(n_3554),
.Y(n_3891)
);

OR3x1_ASAP7_75t_L g3892 ( 
.A(n_3873),
.B(n_3632),
.C(n_3547),
.Y(n_3892)
);

NOR2x1_ASAP7_75t_L g3893 ( 
.A(n_3884),
.B(n_3562),
.Y(n_3893)
);

O2A1O1Ixp33_ASAP7_75t_L g3894 ( 
.A1(n_3879),
.A2(n_3449),
.B(n_3455),
.C(n_3548),
.Y(n_3894)
);

NOR2x1_ASAP7_75t_L g3895 ( 
.A(n_3892),
.B(n_3562),
.Y(n_3895)
);

AND2x4_ASAP7_75t_L g3896 ( 
.A(n_3882),
.B(n_3439),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3886),
.Y(n_3897)
);

O2A1O1Ixp33_ASAP7_75t_L g3898 ( 
.A1(n_3880),
.A2(n_3449),
.B(n_3455),
.C(n_3548),
.Y(n_3898)
);

INVxp67_ASAP7_75t_SL g3899 ( 
.A(n_3882),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3877),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3885),
.Y(n_3901)
);

NOR2xp67_ASAP7_75t_L g3902 ( 
.A(n_3887),
.B(n_3417),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3883),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3876),
.B(n_3570),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3878),
.Y(n_3905)
);

AND2x4_ASAP7_75t_L g3906 ( 
.A(n_3881),
.B(n_3439),
.Y(n_3906)
);

AND3x4_ASAP7_75t_L g3907 ( 
.A(n_3889),
.B(n_3559),
.C(n_3452),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3890),
.Y(n_3908)
);

NOR2x1_ASAP7_75t_L g3909 ( 
.A(n_3875),
.B(n_3562),
.Y(n_3909)
);

AND5x1_ASAP7_75t_L g3910 ( 
.A(n_3894),
.B(n_3891),
.C(n_3888),
.D(n_3544),
.E(n_3532),
.Y(n_3910)
);

INVxp33_ASAP7_75t_L g3911 ( 
.A(n_3895),
.Y(n_3911)
);

NAND3xp33_ASAP7_75t_SL g3912 ( 
.A(n_3900),
.B(n_3571),
.C(n_3579),
.Y(n_3912)
);

NOR3xp33_ASAP7_75t_L g3913 ( 
.A(n_3899),
.B(n_3897),
.C(n_3908),
.Y(n_3913)
);

NOR2x1_ASAP7_75t_L g3914 ( 
.A(n_3905),
.B(n_3893),
.Y(n_3914)
);

NAND3xp33_ASAP7_75t_SL g3915 ( 
.A(n_3901),
.B(n_3571),
.C(n_3579),
.Y(n_3915)
);

NAND3xp33_ASAP7_75t_SL g3916 ( 
.A(n_3903),
.B(n_3571),
.C(n_3579),
.Y(n_3916)
);

NAND4xp25_ASAP7_75t_L g3917 ( 
.A(n_3896),
.B(n_3569),
.C(n_3578),
.D(n_3577),
.Y(n_3917)
);

NAND3xp33_ASAP7_75t_SL g3918 ( 
.A(n_3904),
.B(n_3578),
.C(n_3577),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3909),
.B(n_3570),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3902),
.B(n_3570),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_R g3921 ( 
.A1(n_3910),
.A2(n_3907),
.B1(n_3906),
.B2(n_3898),
.Y(n_3921)
);

AND3x4_ASAP7_75t_L g3922 ( 
.A(n_3913),
.B(n_3559),
.C(n_3532),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3919),
.Y(n_3923)
);

NAND5xp2_ASAP7_75t_L g3924 ( 
.A(n_3911),
.B(n_3575),
.C(n_3569),
.D(n_3583),
.E(n_3518),
.Y(n_3924)
);

NOR2x1_ASAP7_75t_L g3925 ( 
.A(n_3914),
.B(n_3565),
.Y(n_3925)
);

NOR3xp33_ASAP7_75t_L g3926 ( 
.A(n_3916),
.B(n_3460),
.C(n_3569),
.Y(n_3926)
);

AOI22xp33_ASAP7_75t_L g3927 ( 
.A1(n_3925),
.A2(n_3915),
.B1(n_3912),
.B2(n_3918),
.Y(n_3927)
);

AND3x2_ASAP7_75t_L g3928 ( 
.A(n_3923),
.B(n_3920),
.C(n_3445),
.Y(n_3928)
);

AO211x2_ASAP7_75t_L g3929 ( 
.A1(n_3921),
.A2(n_3917),
.B(n_3583),
.C(n_3484),
.Y(n_3929)
);

OR3x2_ASAP7_75t_L g3930 ( 
.A(n_3928),
.B(n_3924),
.C(n_3922),
.Y(n_3930)
);

HB1xp67_ASAP7_75t_L g3931 ( 
.A(n_3929),
.Y(n_3931)
);

OAI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3930),
.A2(n_3927),
.B1(n_3926),
.B2(n_3547),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3932),
.A2(n_3931),
.B1(n_3547),
.B2(n_3573),
.Y(n_3933)
);

OAI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3933),
.A2(n_3573),
.B(n_3570),
.Y(n_3934)
);

OAI22x1_ASAP7_75t_L g3935 ( 
.A1(n_3934),
.A2(n_3460),
.B1(n_3466),
.B2(n_3463),
.Y(n_3935)
);

INVxp67_ASAP7_75t_L g3936 ( 
.A(n_3935),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3936),
.Y(n_3937)
);

NAND4xp25_ASAP7_75t_L g3938 ( 
.A(n_3937),
.B(n_3460),
.C(n_3466),
.D(n_3511),
.Y(n_3938)
);

OAI22xp5_ASAP7_75t_SL g3939 ( 
.A1(n_3938),
.A2(n_3459),
.B1(n_3451),
.B2(n_3448),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3939),
.A2(n_3511),
.B(n_3573),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3940),
.Y(n_3941)
);

OAI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3941),
.A2(n_3462),
.B1(n_3461),
.B2(n_3463),
.Y(n_3942)
);

OAI221xp5_ASAP7_75t_R g3943 ( 
.A1(n_3942),
.A2(n_3532),
.B1(n_3538),
.B2(n_3548),
.C(n_3544),
.Y(n_3943)
);

AOI21xp33_ASAP7_75t_SL g3944 ( 
.A1(n_3943),
.A2(n_3462),
.B(n_3461),
.Y(n_3944)
);

AOI211xp5_ASAP7_75t_L g3945 ( 
.A1(n_3944),
.A2(n_3448),
.B(n_3451),
.C(n_3446),
.Y(n_3945)
);


endmodule