module fake_netlist_6_1932_n_2068 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2068);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2068;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2017;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_3),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_146),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_29),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_61),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_5),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_89),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_52),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_53),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_77),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_88),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_78),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_6),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_16),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_14),
.Y(n_233)
);

BUFx2_ASAP7_75t_R g234 ( 
.A(n_19),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_49),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_64),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_170),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_72),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_123),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_44),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_59),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_98),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_18),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_113),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_103),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_134),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_109),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_81),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_96),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_60),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_176),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_64),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_186),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_26),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_106),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_50),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_22),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_76),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_108),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_172),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_9),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_49),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_153),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_117),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_41),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_188),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_51),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_133),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_151),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_25),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_156),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_120),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_25),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_142),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_194),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_37),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_167),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_179),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_58),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_28),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_112),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_6),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_130),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_66),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_148),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_48),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

INVxp67_ASAP7_75t_R g306 ( 
.A(n_40),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_185),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_136),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_44),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_21),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_93),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_182),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_181),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_114),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_161),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_126),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_55),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_94),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_122),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_33),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_33),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_9),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_19),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_152),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_4),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_83),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_87),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_72),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_99),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_199),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_41),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_35),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_11),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_155),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_75),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_1),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_100),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_169),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_202),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_21),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_197),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_34),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_129),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_165),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_67),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_57),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_5),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_163),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_60),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_0),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_195),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_47),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_18),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_45),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_30),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_42),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_63),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_3),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_174),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_24),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_29),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_2),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_196),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_84),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_85),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_192),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_138),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_54),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_69),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_191),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_140),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_4),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_69),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_22),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_54),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_24),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_141),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_50),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_1),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_154),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_55),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_39),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_70),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_171),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_183),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_46),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_32),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_90),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_101),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_111),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_119),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_39),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_68),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_128),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_61),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_145),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_66),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_46),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_160),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_104),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_11),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_127),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_178),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_37),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_31),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_162),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_268),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_268),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_225),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_318),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_212),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_318),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_208),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_253),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_322),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_206),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_212),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_210),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_214),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_214),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_215),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_292),
.B(n_0),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_249),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_218),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_343),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_219),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_292),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_269),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_269),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_205),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_227),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_211),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_224),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_213),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_225),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_227),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_221),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_233),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_228),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_223),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_226),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_241),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_281),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_235),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_236),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_228),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_230),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_231),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_341),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_242),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_231),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_295),
.B(n_2),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_237),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_240),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_241),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_240),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_R g466 ( 
.A(n_312),
.B(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_248),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_255),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_248),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_250),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_250),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_265),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_243),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_251),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_251),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_281),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_275),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_254),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_254),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_295),
.B(n_327),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_360),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_281),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_232),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_246),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_262),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_277),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_327),
.B(n_7),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_256),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_360),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_280),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_262),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_241),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_341),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_258),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_263),
.B(n_7),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_259),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_354),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_263),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_207),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_270),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_261),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_282),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_301),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_264),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_287),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_270),
.B(n_8),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_272),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_273),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_288),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_272),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_274),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_300),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_274),
.B(n_8),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_279),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_283),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_285),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_241),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_464),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_241),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_427),
.B(n_301),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

CKINVDCx8_ASAP7_75t_R g530 ( 
.A(n_481),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_434),
.A2(n_222),
.B1(n_266),
.B2(n_229),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_416),
.B(n_216),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_461),
.B(n_217),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_435),
.A2(n_344),
.B1(n_352),
.B2(n_358),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_413),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_487),
.B(n_217),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_301),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_286),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_422),
.A2(n_425),
.B(n_424),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_503),
.B(n_289),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_482),
.B(n_290),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_493),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_493),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_482),
.B(n_330),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_493),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_495),
.B(n_312),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_437),
.B(n_330),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_442),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_506),
.B(n_217),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_459),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_465),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_421),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_469),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_470),
.B(n_293),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_474),
.B(n_475),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_478),
.A2(n_312),
.B(n_372),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_491),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_498),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_500),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_436),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_444),
.A2(n_306),
.B1(n_363),
.B2(n_362),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_507),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_513),
.B(n_312),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_499),
.B(n_330),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_419),
.B(n_296),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_483),
.B(n_405),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_421),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_489),
.B(n_405),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_423),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_423),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_565),
.A2(n_306),
.B1(n_387),
.B2(n_466),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_524),
.B(n_405),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_438),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_546),
.B(n_552),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_538),
.A2(n_417),
.B1(n_441),
.B2(n_414),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_567),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_524),
.B(n_598),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_426),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_520),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_564),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_562),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_426),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_562),
.B(n_341),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_538),
.A2(n_417),
.B1(n_308),
.B2(n_313),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_595),
.C(n_592),
.Y(n_622)
);

INVx4_ASAP7_75t_SL g623 ( 
.A(n_562),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_524),
.B(n_598),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_573),
.B(n_598),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_595),
.B(n_429),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_541),
.B(n_440),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_562),
.A2(n_216),
.B1(n_347),
.B2(n_257),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_562),
.A2(n_216),
.B1(n_347),
.B2(n_257),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_555),
.B(n_517),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_567),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_520),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_527),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_567),
.Y(n_636)
);

INVxp33_ASAP7_75t_L g637 ( 
.A(n_593),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_562),
.A2(n_347),
.B1(n_357),
.B2(n_257),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_518),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_545),
.B(n_560),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_545),
.B(n_560),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_562),
.A2(n_374),
.B1(n_357),
.B2(n_284),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_522),
.A2(n_448),
.B1(n_449),
.B2(n_445),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_555),
.B(n_429),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_584),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_573),
.B(n_432),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_528),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_594),
.B(n_432),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_573),
.B(n_439),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_560),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_524),
.B(n_276),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_533),
.Y(n_655)
);

BUFx4f_ASAP7_75t_L g656 ( 
.A(n_562),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_571),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_520),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_533),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_544),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_533),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_545),
.B(n_439),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_526),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_SL g665 ( 
.A1(n_524),
.A2(n_308),
.B1(n_313),
.B2(n_299),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_562),
.A2(n_374),
.B1(n_357),
.B2(n_284),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_529),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_571),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_544),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_571),
.Y(n_672)
);

INVx6_ASAP7_75t_L g673 ( 
.A(n_563),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_599),
.B(n_446),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_517),
.B(n_446),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_523),
.B(n_452),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_599),
.B(n_452),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_562),
.B(n_341),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_568),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_522),
.A2(n_455),
.B1(n_473),
.B2(n_462),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_599),
.B(n_484),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_523),
.B(n_453),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_566),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_529),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_591),
.B(n_488),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_534),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_594),
.B(n_453),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_571),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_596),
.B(n_458),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_534),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_582),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_524),
.B(n_276),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_521),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_575),
.B(n_458),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_521),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_582),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_589),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_593),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_596),
.B(n_468),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_566),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_525),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_530),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_524),
.B(n_276),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_582),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_591),
.B(n_494),
.Y(n_707)
);

INVxp33_ASAP7_75t_L g708 ( 
.A(n_593),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_597),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_525),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_589),
.B(n_468),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_519),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_582),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_589),
.A2(n_374),
.B1(n_380),
.B2(n_207),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_582),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_592),
.A2(n_321),
.B1(n_238),
.B2(n_245),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_530),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_596),
.B(n_472),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_590),
.B(n_472),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_590),
.B(n_477),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_587),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_551),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_544),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_544),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_596),
.B(n_477),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_544),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_530),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_587),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_597),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_587),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_587),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_587),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_551),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_543),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_547),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_589),
.A2(n_380),
.B1(n_377),
.B2(n_324),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_551),
.Y(n_742)
);

BUFx10_ASAP7_75t_L g743 ( 
.A(n_519),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_596),
.B(n_486),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_547),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_566),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_588),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_569),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_574),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_575),
.B(n_496),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_588),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_646),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_610),
.B(n_589),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_652),
.B(n_590),
.Y(n_755)
);

NOR3xp33_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_559),
.C(n_527),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_737),
.A2(n_738),
.B(n_742),
.C(n_699),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_656),
.B(n_341),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_656),
.B(n_393),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_699),
.A2(n_589),
.B1(n_504),
.B2(n_508),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_653),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_719),
.B(n_486),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_601),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_637),
.B(n_597),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_673),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_601),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_618),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_702),
.A2(n_589),
.B1(n_239),
.B2(n_247),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_702),
.B(n_238),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_708),
.B(n_501),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_628),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_628),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_737),
.A2(n_589),
.B(n_578),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_607),
.B(n_559),
.C(n_527),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_686),
.A2(n_589),
.B1(n_515),
.B2(n_516),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_679),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_656),
.B(n_393),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_589),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_707),
.A2(n_750),
.B1(n_641),
.B2(n_640),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_675),
.B(n_514),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_618),
.B(n_698),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_618),
.B(n_393),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_722),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_680),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_726),
.Y(n_785)
);

AOI221xp5_ASAP7_75t_L g786 ( 
.A1(n_611),
.A2(n_585),
.B1(n_336),
.B2(n_244),
.C(n_247),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_640),
.B(n_588),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_650),
.B(n_559),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_748),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_618),
.B(n_578),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_749),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_490),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_618),
.B(n_393),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_747),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_738),
.A2(n_239),
.B(n_260),
.C(n_244),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_641),
.B(n_588),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_663),
.B(n_537),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_652),
.B(n_566),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_715),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_490),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_566),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_751),
.Y(n_802)
);

AOI22x1_ASAP7_75t_L g803 ( 
.A1(n_742),
.A2(n_590),
.B1(n_505),
.B2(n_509),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_698),
.B(n_393),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_751),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_715),
.A2(n_536),
.B(n_577),
.C(n_574),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_673),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_673),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_673),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_698),
.B(n_393),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_710),
.B(n_733),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_710),
.B(n_566),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_733),
.B(n_572),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_627),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_SL g815 ( 
.A1(n_704),
.A2(n_428),
.B1(n_430),
.B2(n_418),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_502),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_627),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_698),
.A2(n_678),
.B(n_620),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_698),
.B(n_572),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_639),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_645),
.B(n_572),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_695),
.B(n_502),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_606),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_623),
.B(n_572),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_725),
.B(n_572),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_682),
.Y(n_826)
);

INVx8_ASAP7_75t_L g827 ( 
.A(n_654),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_725),
.B(n_572),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_612),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_623),
.B(n_630),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_722),
.B(n_590),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_635),
.B(n_537),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_623),
.B(n_572),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_623),
.B(n_572),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_563),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_676),
.B(n_540),
.Y(n_836)
);

INVx8_ASAP7_75t_L g837 ( 
.A(n_654),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_612),
.Y(n_838)
);

AND2x6_ASAP7_75t_SL g839 ( 
.A(n_683),
.B(n_260),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_625),
.B(n_505),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_609),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_642),
.B(n_563),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_723),
.B(n_540),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_631),
.B(n_550),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_614),
.A2(n_585),
.B1(n_532),
.B2(n_539),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_723),
.A2(n_550),
.B1(n_563),
.B2(n_509),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_668),
.B(n_563),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_716),
.B(n_570),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_638),
.B(n_303),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_613),
.B(n_570),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_633),
.B(n_570),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_633),
.B(n_576),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_739),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_636),
.B(n_576),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_622),
.A2(n_267),
.B(n_271),
.C(n_291),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_604),
.B(n_650),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_646),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_639),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_688),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_657),
.B(n_576),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_712),
.B(n_372),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_657),
.B(n_581),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_688),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_670),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_621),
.A2(n_536),
.B(n_577),
.C(n_580),
.Y(n_865)
);

BUFx12f_ASAP7_75t_SL g866 ( 
.A(n_654),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_670),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_672),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_674),
.B(n_586),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_614),
.A2(n_238),
.B1(n_396),
.B2(n_245),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_665),
.B(n_376),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_713),
.B(n_532),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_677),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_648),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_672),
.Y(n_875)
);

BUFx12f_ASAP7_75t_L g876 ( 
.A(n_713),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_689),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_644),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_651),
.B(n_539),
.C(n_579),
.Y(n_879)
);

NAND3xp33_ASAP7_75t_L g880 ( 
.A(n_690),
.B(n_580),
.C(n_579),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_620),
.A2(n_586),
.B(n_583),
.C(n_581),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_644),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_689),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_692),
.B(n_581),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_700),
.B(n_302),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_647),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_704),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_692),
.B(n_583),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_614),
.A2(n_321),
.B1(n_245),
.B2(n_252),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_647),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_697),
.A2(n_396),
.B(n_317),
.C(n_369),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_706),
.B(n_376),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_717),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_721),
.B(n_209),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_L g895 ( 
.A(n_719),
.B(n_305),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_654),
.B(n_583),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_649),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_649),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_717),
.B(n_736),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_729),
.B(n_220),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_744),
.A2(n_353),
.B1(n_370),
.B2(n_340),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_713),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_736),
.B(n_714),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_694),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_714),
.B(n_309),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_655),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_694),
.B(n_535),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_696),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_743),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_696),
.B(n_535),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_703),
.B(n_542),
.Y(n_911)
);

AO22x2_ASAP7_75t_L g912 ( 
.A1(n_718),
.A2(n_321),
.B1(n_317),
.B2(n_252),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_703),
.B(n_542),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_711),
.B(n_548),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_711),
.B(n_548),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_693),
.B(n_310),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_724),
.B(n_553),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_753),
.A2(n_678),
.B(n_624),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_752),
.B(n_731),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_797),
.B(n_743),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_857),
.B(n_731),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_779),
.B(n_614),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_778),
.A2(n_624),
.B(n_603),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_823),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_857),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_799),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_755),
.B(n_624),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_832),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_799),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_870),
.A2(n_338),
.B(n_299),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_768),
.A2(n_760),
.B1(n_775),
.B2(n_894),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_755),
.B(n_624),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_831),
.B(n_693),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_792),
.B(n_724),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_773),
.A2(n_734),
.B(n_732),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_841),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_827),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_767),
.A2(n_603),
.B(n_602),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_819),
.A2(n_739),
.B(n_734),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_767),
.A2(n_818),
.B(n_768),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_799),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_781),
.A2(n_603),
.B(n_602),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_799),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_792),
.B(n_800),
.Y(n_944)
);

NAND2x1_ASAP7_75t_L g945 ( 
.A(n_829),
.B(n_600),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_794),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_781),
.A2(n_684),
.B(n_602),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_825),
.A2(n_701),
.B(n_684),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_800),
.B(n_732),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_757),
.A2(n_735),
.B(n_578),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_826),
.B(n_831),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_787),
.B(n_735),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_802),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_828),
.A2(n_701),
.B(n_684),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_816),
.B(n_743),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_827),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_600),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_765),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_764),
.B(n_600),
.Y(n_959)
);

AOI222xp33_ASAP7_75t_L g960 ( 
.A1(n_786),
.A2(n_367),
.B1(n_336),
.B2(n_331),
.C1(n_324),
.C2(n_307),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_830),
.A2(n_746),
.B(n_701),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_780),
.B(n_608),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_780),
.B(n_811),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_821),
.A2(n_746),
.B(n_616),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_894),
.A2(n_605),
.B1(n_681),
.B2(n_643),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_900),
.B(n_608),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_900),
.B(n_608),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_754),
.B(n_658),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_761),
.B(n_658),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_819),
.A2(n_660),
.B(n_655),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_776),
.B(n_658),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_816),
.B(n_693),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_783),
.B(n_856),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_856),
.B(n_612),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_771),
.A2(n_605),
.B1(n_693),
.B2(n_705),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_843),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_805),
.Y(n_977)
);

AO21x1_ASAP7_75t_L g978 ( 
.A1(n_889),
.A2(n_342),
.B(n_338),
.Y(n_978)
);

AO21x1_ASAP7_75t_L g979 ( 
.A1(n_861),
.A2(n_368),
.B(n_342),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_842),
.A2(n_616),
.B(n_612),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_864),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_SL g982 ( 
.A(n_876),
.B(n_234),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_806),
.A2(n_671),
.B(n_667),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_765),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_847),
.A2(n_835),
.B(n_798),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_784),
.B(n_667),
.Y(n_986)
);

CKINVDCx10_ASAP7_75t_R g987 ( 
.A(n_815),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_867),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_812),
.A2(n_616),
.B(n_612),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_772),
.B(n_705),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_887),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_785),
.B(n_667),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_874),
.B(n_664),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_813),
.A2(n_626),
.B(n_616),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_861),
.A2(n_720),
.B(n_671),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_758),
.A2(n_634),
.B(n_626),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_789),
.B(n_671),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_758),
.A2(n_634),
.B(n_626),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_868),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_791),
.B(n_720),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_822),
.A2(n_605),
.B1(n_705),
.B2(n_718),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_869),
.B(n_720),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_869),
.B(n_822),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_859),
.B(n_705),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_759),
.A2(n_634),
.B(n_626),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_844),
.A2(n_605),
.B(n_685),
.C(n_669),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_865),
.B(n_727),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_844),
.B(n_727),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_759),
.A2(n_634),
.B(n_626),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_866),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_904),
.B(n_727),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_875),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_756),
.B(n_774),
.Y(n_1013)
);

AO21x1_ASAP7_75t_L g1014 ( 
.A1(n_777),
.A2(n_401),
.B(n_368),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_908),
.B(n_730),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_840),
.B(n_730),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_840),
.B(n_730),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_788),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_863),
.B(n_740),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_896),
.B(n_873),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_829),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_777),
.A2(n_659),
.B(n_634),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_896),
.B(n_659),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_877),
.B(n_740),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_770),
.B(n_740),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_883),
.B(n_745),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_899),
.A2(n_745),
.B(n_662),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_899),
.A2(n_745),
.B(n_662),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_769),
.B(n_664),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_829),
.A2(n_661),
.B(n_659),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_770),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_902),
.B(n_360),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_879),
.B(n_323),
.C(n_311),
.Y(n_1034)
);

OAI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_901),
.A2(n_326),
.B(n_325),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_845),
.A2(n_401),
.B(n_334),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_829),
.A2(n_838),
.B(n_848),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_807),
.B(n_659),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_763),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_769),
.B(n_666),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_850),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_769),
.B(n_669),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_795),
.A2(n_377),
.B(n_331),
.C(n_398),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_838),
.A2(n_661),
.B(n_659),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_769),
.B(n_685),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_851),
.B(n_687),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_838),
.A2(n_709),
.B(n_661),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_808),
.B(n_661),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_809),
.A2(n_718),
.B1(n_687),
.B2(n_691),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_766),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_795),
.A2(n_367),
.B(n_400),
.C(n_398),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_855),
.A2(n_916),
.B(n_881),
.C(n_846),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_762),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_824),
.A2(n_728),
.B(n_709),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_852),
.B(n_691),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_824),
.A2(n_728),
.B(n_709),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_845),
.B(n_328),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_855),
.A2(n_378),
.B(n_307),
.C(n_381),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_854),
.B(n_718),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_833),
.A2(n_728),
.B(n_709),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_827),
.B(n_267),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_833),
.A2(n_728),
.B(n_549),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_834),
.A2(n_728),
.B(n_549),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_837),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_860),
.B(n_660),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_872),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_834),
.A2(n_801),
.B(n_903),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_862),
.A2(n_549),
.B(n_547),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_884),
.A2(n_549),
.B(n_547),
.Y(n_1069)
);

NOR2xp67_ASAP7_75t_L g1070 ( 
.A(n_909),
.B(n_314),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_888),
.A2(n_891),
.B(n_790),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_803),
.B(n_252),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_814),
.B(n_278),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_817),
.B(n_278),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_907),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_820),
.B(n_278),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_858),
.B(n_317),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_885),
.B(n_335),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_878),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_882),
.B(n_369),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_886),
.B(n_369),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_849),
.A2(n_558),
.B(n_547),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_890),
.B(n_396),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_917),
.A2(n_558),
.B(n_547),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_897),
.B(n_315),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_853),
.Y(n_1086)
);

AO21x1_ASAP7_75t_L g1087 ( 
.A1(n_871),
.A2(n_892),
.B(n_836),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_916),
.B(n_339),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_839),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_837),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_898),
.B(n_316),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_906),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_880),
.A2(n_294),
.B(n_271),
.C(n_291),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_910),
.A2(n_558),
.B(n_547),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_871),
.B(n_345),
.C(n_350),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_837),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_895),
.B(n_294),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_911),
.A2(n_558),
.B(n_547),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_892),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_905),
.A2(n_375),
.B1(n_320),
.B2(n_329),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_790),
.B(n_384),
.C(n_355),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_913),
.A2(n_558),
.B(n_549),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_914),
.B(n_319),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_920),
.B(n_912),
.Y(n_1104)
);

BUFx4f_ASAP7_75t_L g1105 ( 
.A(n_1096),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_944),
.B(n_853),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_SL g1107 ( 
.A(n_1096),
.B(n_782),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_981),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1003),
.A2(n_912),
.B1(n_915),
.B2(n_810),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1088),
.A2(n_782),
.B(n_810),
.C(n_804),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_976),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_946),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_931),
.A2(n_297),
.B1(n_298),
.B2(n_304),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_946),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_912),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_963),
.B(n_793),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1066),
.B(n_793),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1041),
.B(n_804),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_925),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_953),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_925),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1075),
.B(n_1025),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1025),
.B(n_332),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_929),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1036),
.A2(n_973),
.B(n_965),
.C(n_1088),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_940),
.A2(n_985),
.B(n_918),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_922),
.A2(n_389),
.B1(n_364),
.B2(n_371),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1001),
.A2(n_390),
.B1(n_346),
.B2(n_348),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_972),
.A2(n_385),
.B1(n_394),
.B2(n_395),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_929),
.B(n_934),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_923),
.A2(n_558),
.B(n_549),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_973),
.B(n_333),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_991),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1078),
.A2(n_391),
.B(n_297),
.C(n_298),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_929),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_1072),
.A2(n_1087),
.B(n_979),
.C(n_962),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_949),
.B(n_337),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_988),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_964),
.A2(n_558),
.B(n_549),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_953),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_977),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_948),
.A2(n_558),
.B(n_549),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1057),
.A2(n_392),
.B1(n_304),
.B2(n_378),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1078),
.B(n_349),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_988),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_977),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_974),
.A2(n_399),
.B1(n_356),
.B2(n_382),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1018),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_999),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_954),
.A2(n_531),
.B(n_553),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1092),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_990),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1057),
.A2(n_381),
.B1(n_391),
.B2(n_392),
.Y(n_1153)
);

BUFx8_ASAP7_75t_SL g1154 ( 
.A(n_1010),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_980),
.A2(n_531),
.B(n_557),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1032),
.B(n_359),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1032),
.B(n_361),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_955),
.B(n_360),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_957),
.A2(n_531),
.B(n_557),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_974),
.A2(n_561),
.B(n_557),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_929),
.B(n_404),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1096),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1096),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_952),
.A2(n_531),
.B(n_556),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1006),
.A2(n_531),
.B(n_556),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_999),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1037),
.A2(n_561),
.B(n_556),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_951),
.B(n_365),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_993),
.B(n_407),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_366),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1028),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_927),
.A2(n_408),
.B1(n_403),
.B2(n_373),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1013),
.B(n_379),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_951),
.B(n_383),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1039),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_933),
.B(n_217),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_932),
.A2(n_406),
.B1(n_388),
.B2(n_397),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1020),
.B(n_386),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1020),
.B(n_402),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1013),
.B(n_990),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_924),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1016),
.A2(n_410),
.B1(n_409),
.B2(n_400),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1052),
.A2(n_561),
.B(n_554),
.C(n_543),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1052),
.A2(n_554),
.B(n_543),
.C(n_13),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_936),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_SL g1186 ( 
.A(n_1089),
.B(n_554),
.C(n_12),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_943),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1004),
.A2(n_10),
.B(n_13),
.C(n_15),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1017),
.A2(n_204),
.B1(n_200),
.B2(n_198),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_960),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1004),
.B(n_17),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1012),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_921),
.B(n_193),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1092),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1039),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_933),
.A2(n_189),
.B1(n_187),
.B2(n_177),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_961),
.A2(n_1002),
.B(n_1030),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_926),
.B(n_175),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_926),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1050),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_975),
.A2(n_173),
.B1(n_164),
.B2(n_157),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_R g1202 ( 
.A(n_1053),
.B(n_147),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1040),
.A2(n_143),
.B(n_139),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1034),
.B(n_23),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_919),
.B(n_132),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_941),
.A2(n_116),
.B1(n_115),
.B2(n_110),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1019),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_959),
.B(n_27),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1019),
.B(n_27),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1064),
.B(n_91),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_SL g1211 ( 
.A(n_982),
.B(n_1064),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1050),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1079),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_943),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1086),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1099),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1093),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1046),
.B(n_38),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1042),
.A2(n_97),
.B(n_92),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1097),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_941),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1095),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1045),
.A2(n_80),
.B(n_79),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1035),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1055),
.B(n_53),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1061),
.B(n_56),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_968),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_969),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_971),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1023),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1067),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_986),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_970),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1071),
.A2(n_74),
.B(n_63),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_966),
.B(n_62),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_967),
.B(n_62),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1061),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_958),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1065),
.B(n_65),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1021),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1007),
.B(n_1008),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1090),
.B(n_65),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_939),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1023),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_1246)
);

AOI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1085),
.A2(n_71),
.B(n_73),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_992),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_958),
.B(n_984),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1021),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_984),
.B(n_997),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1090),
.B(n_937),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1103),
.B(n_1070),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_987),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_950),
.A2(n_983),
.B(n_935),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_937),
.B(n_956),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1059),
.B(n_945),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1061),
.B(n_956),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1093),
.B(n_1058),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_942),
.A2(n_947),
.B(n_994),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1126),
.A2(n_930),
.A3(n_978),
.B(n_1014),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1119),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1125),
.A2(n_995),
.B(n_1081),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1134),
.A2(n_1058),
.B(n_1043),
.C(n_1051),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1111),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1250),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1158),
.B(n_1043),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_1083),
.B(n_1080),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1181),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1133),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_R g1271 ( 
.A(n_1194),
.B(n_1091),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1197),
.A2(n_989),
.B(n_938),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_SL g1273 ( 
.A1(n_1225),
.A2(n_1051),
.B(n_1038),
.C(n_1048),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1152),
.A2(n_1074),
.B(n_1077),
.C(n_1076),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1148),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1170),
.B(n_1000),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1184),
.A2(n_1048),
.B(n_1038),
.C(n_1026),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1131),
.A2(n_1022),
.B(n_996),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1173),
.A2(n_1180),
.B1(n_1190),
.B2(n_1191),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_998),
.B(n_1005),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1110),
.A2(n_1073),
.A3(n_1082),
.B(n_1009),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1156),
.B(n_1049),
.Y(n_1282)
);

AO32x2_ASAP7_75t_L g1283 ( 
.A1(n_1109),
.A2(n_1027),
.A3(n_1029),
.B1(n_1069),
.B2(n_1068),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_SL g1284 ( 
.A(n_1241),
.B(n_1024),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1122),
.B(n_1242),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1242),
.A2(n_1031),
.B(n_1044),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1207),
.B(n_1011),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1156),
.B(n_1100),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1252),
.B(n_1015),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1142),
.A2(n_1047),
.B(n_1054),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1243),
.B(n_1056),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1207),
.B(n_1060),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1255),
.A2(n_1094),
.B(n_1098),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1108),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1179),
.B(n_1062),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1241),
.B(n_1063),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1167),
.A2(n_1084),
.B(n_1102),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1165),
.A2(n_1232),
.A3(n_1234),
.B(n_1245),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_1139),
.B(n_1150),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1255),
.A2(n_1249),
.B(n_1251),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1136),
.A2(n_1183),
.B(n_1106),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1255),
.A2(n_1249),
.B(n_1251),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1241),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1236),
.A2(n_1237),
.B(n_1130),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1305)
);

NOR4xp25_ASAP7_75t_L g1306 ( 
.A(n_1190),
.B(n_1113),
.C(n_1223),
.D(n_1188),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1185),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1121),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1130),
.A2(n_1164),
.B(n_1152),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1159),
.A2(n_1203),
.B(n_1220),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1180),
.A2(n_1191),
.B1(n_1113),
.B2(n_1104),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1144),
.A2(n_1168),
.B(n_1178),
.C(n_1219),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1211),
.B(n_1221),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1157),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1224),
.A2(n_1239),
.B(n_1198),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1230),
.B(n_1233),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1239),
.A2(n_1198),
.B(n_1140),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1241),
.A2(n_1123),
.B(n_1118),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1154),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1137),
.A2(n_1248),
.B(n_1135),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_SL g1321 ( 
.A1(n_1218),
.A2(n_1208),
.B(n_1201),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1138),
.B(n_1145),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1157),
.B(n_1168),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1178),
.B(n_1115),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1171),
.B(n_1112),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1221),
.B(n_1253),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1176),
.A2(n_1193),
.B1(n_1174),
.B2(n_1161),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1135),
.A2(n_1257),
.B(n_1161),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1192),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1240),
.A2(n_1226),
.B(n_1209),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1199),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1189),
.A2(n_1246),
.A3(n_1128),
.B(n_1182),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1132),
.A2(n_1149),
.A3(n_1146),
.B(n_1114),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1169),
.A2(n_1120),
.B(n_1166),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1176),
.A2(n_1129),
.B1(n_1127),
.B2(n_1172),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1141),
.B(n_1259),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1105),
.A2(n_1231),
.B(n_1199),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1231),
.A2(n_1247),
.B(n_1196),
.C(n_1217),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1175),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1210),
.A2(n_1250),
.B(n_1252),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1195),
.A2(n_1212),
.B(n_1200),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1244),
.A2(n_1143),
.B(n_1153),
.C(n_1204),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1258),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1186),
.A2(n_1217),
.B(n_1223),
.C(n_1177),
.Y(n_1344)
);

INVxp67_ASAP7_75t_SL g1345 ( 
.A(n_1124),
.Y(n_1345)
);

AO21x1_ASAP7_75t_L g1346 ( 
.A1(n_1206),
.A2(n_1147),
.B(n_1214),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1143),
.A2(n_1153),
.B1(n_1210),
.B2(n_1238),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1213),
.B(n_1222),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1256),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1107),
.A2(n_1216),
.B(n_1117),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1105),
.B(n_1205),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1250),
.A2(n_1124),
.B(n_1215),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1250),
.A2(n_1124),
.B(n_1215),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1124),
.B(n_1162),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1256),
.B(n_1254),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1162),
.Y(n_1356)
);

BUFx10_ASAP7_75t_L g1357 ( 
.A(n_1162),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1162),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1227),
.A2(n_1187),
.B(n_1205),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1187),
.A2(n_1163),
.B(n_1151),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1163),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1163),
.A2(n_1126),
.A3(n_1184),
.B(n_1110),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1163),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1202),
.B(n_1122),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1202),
.A2(n_1126),
.B(n_1260),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_607),
.B2(n_780),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1126),
.A2(n_1184),
.A3(n_1110),
.B(n_1242),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1125),
.A2(n_1136),
.B(n_1242),
.Y(n_1372)
);

CKINVDCx16_ASAP7_75t_R g1373 ( 
.A(n_1133),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1105),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1122),
.B(n_944),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1130),
.A2(n_1160),
.B(n_1197),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_1088),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_607),
.B2(n_780),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1126),
.A2(n_1184),
.A3(n_1110),
.B(n_1242),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1181),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1108),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_629),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1133),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1125),
.A2(n_931),
.B(n_1110),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1126),
.A2(n_656),
.B(n_944),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_629),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_1088),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1126),
.A2(n_1184),
.A3(n_1110),
.B(n_1242),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1397)
);

AO32x2_ASAP7_75t_L g1398 ( 
.A1(n_1109),
.A2(n_931),
.A3(n_1246),
.B1(n_1182),
.B2(n_889),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1111),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1400)
);

AOI221x1_ASAP7_75t_L g1401 ( 
.A1(n_1235),
.A2(n_944),
.B1(n_931),
.B2(n_1184),
.C(n_1232),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1126),
.A2(n_1184),
.A3(n_1110),
.B(n_1242),
.Y(n_1402)
);

INVx3_ASAP7_75t_SL g1403 ( 
.A(n_1133),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_629),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1126),
.A2(n_656),
.B(n_618),
.Y(n_1405)
);

CKINVDCx8_ASAP7_75t_R g1406 ( 
.A(n_1256),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1158),
.B(n_826),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1119),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1190),
.A2(n_944),
.B1(n_1003),
.B2(n_768),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1119),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1133),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1190),
.A2(n_944),
.B1(n_1003),
.B2(n_768),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_SL g1413 ( 
.A(n_1194),
.B(n_857),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1122),
.B(n_944),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_SL g1415 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_1225),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1119),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_629),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1252),
.B(n_937),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_607),
.B2(n_780),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1125),
.B(n_944),
.C(n_1003),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1194),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_SL g1423 ( 
.A1(n_1125),
.A2(n_944),
.B(n_1003),
.C(n_1225),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1131),
.A2(n_1160),
.B(n_1260),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1158),
.B(n_826),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1133),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1126),
.A2(n_1260),
.B(n_1197),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1133),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_1378),
.B2(n_1419),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1428),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1409),
.A2(n_1412),
.B1(n_1367),
.B2(n_1311),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1288),
.A2(n_1412),
.B1(n_1409),
.B2(n_1314),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1294),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1374),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1374),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1307),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1374),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1420),
.A2(n_1282),
.B1(n_1425),
.B2(n_1407),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1262),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1410),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1285),
.A2(n_1414),
.B1(n_1375),
.B2(n_1342),
.Y(n_1441)
);

INVx8_ASAP7_75t_L g1442 ( 
.A(n_1361),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1420),
.A2(n_1324),
.B1(n_1267),
.B2(n_1335),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1321),
.A2(n_1276),
.B1(n_1364),
.B2(n_1313),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1422),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1270),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1364),
.A2(n_1347),
.B1(n_1359),
.B2(n_1330),
.Y(n_1447)
);

BUFx8_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1329),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1373),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1285),
.A2(n_1375),
.B1(n_1414),
.B2(n_1382),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1359),
.A2(n_1330),
.B1(n_1327),
.B2(n_1372),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1306),
.A2(n_1403),
.B1(n_1406),
.B2(n_1411),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1372),
.A2(n_1295),
.B1(n_1275),
.B2(n_1343),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1357),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1357),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1351),
.A2(n_1326),
.B1(n_1399),
.B2(n_1346),
.Y(n_1457)
);

INVx11_ASAP7_75t_L g1458 ( 
.A(n_1340),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1380),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1356),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1331),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1356),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1291),
.A2(n_1289),
.B1(n_1320),
.B2(n_1304),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1365),
.B1(n_1336),
.B2(n_1349),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1306),
.A2(n_1386),
.B1(n_1344),
.B2(n_1305),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1381),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1305),
.B(n_1316),
.Y(n_1467)
);

BUFx4_ASAP7_75t_R g1468 ( 
.A(n_1416),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1385),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1339),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1365),
.A2(n_1336),
.B1(n_1316),
.B2(n_1292),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1292),
.A2(n_1287),
.B1(n_1318),
.B2(n_1413),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1401),
.A2(n_1355),
.B1(n_1287),
.B2(n_1337),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1354),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1377),
.A2(n_1393),
.B1(n_1417),
.B2(n_1392),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1325),
.Y(n_1476)
);

AND2x4_ASAP7_75t_SL g1477 ( 
.A(n_1418),
.B(n_1408),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1426),
.A2(n_1308),
.B1(n_1360),
.B2(n_1350),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1328),
.A2(n_1322),
.B1(n_1341),
.B2(n_1303),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1418),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1309),
.A2(n_1334),
.B1(n_1389),
.B2(n_1341),
.Y(n_1481)
);

OAI21xp33_ASAP7_75t_L g1482 ( 
.A1(n_1404),
.A2(n_1312),
.B(n_1309),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1389),
.A2(n_1301),
.B1(n_1302),
.B2(n_1300),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1356),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1348),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1354),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1363),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1338),
.A2(n_1398),
.B1(n_1301),
.B2(n_1415),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1333),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1333),
.Y(n_1491)
);

CKINVDCx11_ASAP7_75t_R g1492 ( 
.A(n_1271),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1266),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1358),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1358),
.B(n_1317),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1345),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1352),
.A2(n_1353),
.B1(n_1296),
.B2(n_1286),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1296),
.A2(n_1286),
.B1(n_1398),
.B2(n_1423),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1263),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1284),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1264),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1315),
.B(n_1310),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1298),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1273),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1398),
.A2(n_1332),
.B1(n_1427),
.B2(n_1402),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1362),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1277),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1332),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_R g1509 ( 
.A1(n_1332),
.A2(n_1379),
.B1(n_1402),
.B2(n_1395),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1272),
.A2(n_1397),
.B1(n_1391),
.B2(n_1371),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1370),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1427),
.A2(n_1395),
.B1(n_1379),
.B2(n_1370),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1268),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1268),
.A2(n_1293),
.B1(n_1384),
.B2(n_1390),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1274),
.A2(n_1405),
.B1(n_1394),
.B2(n_1387),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1379),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1402),
.B(n_1261),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1299),
.A2(n_1368),
.B1(n_1421),
.B2(n_1400),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1283),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1376),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1261),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1366),
.A2(n_1424),
.B1(n_1396),
.B2(n_1388),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1278),
.Y(n_1523)
);

CKINVDCx11_ASAP7_75t_R g1524 ( 
.A(n_1283),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1283),
.A2(n_1281),
.B1(n_1369),
.B2(n_1383),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1280),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1290),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1297),
.A2(n_1323),
.B1(n_1412),
.B2(n_1409),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1374),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1367),
.A2(n_1419),
.B1(n_1378),
.B2(n_944),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1279),
.A2(n_1190),
.B1(n_944),
.B2(n_1409),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1374),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1269),
.Y(n_1535)
);

INVx6_ASAP7_75t_L g1536 ( 
.A(n_1374),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1537)
);

BUFx10_ASAP7_75t_L g1538 ( 
.A(n_1270),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1428),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1374),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1279),
.A2(n_1190),
.B1(n_944),
.B2(n_1409),
.Y(n_1541)
);

CKINVDCx9p33_ASAP7_75t_R g1542 ( 
.A(n_1319),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1265),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1262),
.Y(n_1544)
);

INVx8_ASAP7_75t_L g1545 ( 
.A(n_1361),
.Y(n_1545)
);

INVx5_ASAP7_75t_L g1546 ( 
.A(n_1374),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1262),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1367),
.A2(n_944),
.B1(n_1419),
.B2(n_1378),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1279),
.A2(n_1190),
.B1(n_944),
.B2(n_1367),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1262),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1323),
.A2(n_1409),
.B1(n_1412),
.B2(n_944),
.Y(n_1551)
);

BUFx5_ASAP7_75t_L g1552 ( 
.A(n_1357),
.Y(n_1552)
);

BUFx10_ASAP7_75t_L g1553 ( 
.A(n_1270),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1428),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1275),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1285),
.B(n_1375),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1323),
.A2(n_1409),
.B1(n_1412),
.B2(n_944),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1269),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1294),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1418),
.B(n_1252),
.Y(n_1562)
);

BUFx10_ASAP7_75t_L g1563 ( 
.A(n_1270),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1428),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1566)
);

OAI22x1_ASAP7_75t_L g1567 ( 
.A1(n_1367),
.A2(n_1419),
.B1(n_1378),
.B2(n_1180),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1262),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1279),
.A2(n_1190),
.B1(n_944),
.B2(n_1409),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1294),
.Y(n_1571)
);

INVx6_ASAP7_75t_L g1572 ( 
.A(n_1374),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1294),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1279),
.A2(n_1323),
.B1(n_944),
.B2(n_1367),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1374),
.Y(n_1575)
);

INVx5_ASAP7_75t_L g1576 ( 
.A(n_1374),
.Y(n_1576)
);

BUFx10_ASAP7_75t_L g1577 ( 
.A(n_1270),
.Y(n_1577)
);

CKINVDCx6p67_ASAP7_75t_R g1578 ( 
.A(n_1403),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1351),
.B(n_1241),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1523),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1508),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1549),
.A2(n_1541),
.B1(n_1532),
.B2(n_1569),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1490),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1458),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1491),
.Y(n_1585)
);

INVxp33_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1503),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1511),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1506),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1495),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1520),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1516),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1524),
.B(n_1528),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1521),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1486),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1517),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1502),
.A2(n_1518),
.B(n_1515),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1517),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1509),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1461),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1455),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1467),
.B(n_1558),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1461),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1495),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1532),
.A2(n_1569),
.B1(n_1541),
.B2(n_1431),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1528),
.B(n_1465),
.Y(n_1606)
);

CKINVDCx14_ASAP7_75t_R g1607 ( 
.A(n_1539),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1465),
.B(n_1551),
.Y(n_1608)
);

BUFx2_ASAP7_75t_SL g1609 ( 
.A(n_1437),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1500),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1513),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1431),
.A2(n_1531),
.B1(n_1429),
.B2(n_1548),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1551),
.B(n_1559),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1436),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1504),
.Y(n_1615)
);

BUFx4f_ASAP7_75t_SL g1616 ( 
.A(n_1430),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1452),
.B(n_1483),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1513),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1543),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1559),
.B(n_1432),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1510),
.A2(n_1498),
.B(n_1515),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1558),
.A2(n_1533),
.B(n_1529),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1522),
.A2(n_1514),
.B(n_1525),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1525),
.A2(n_1527),
.B(n_1526),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1519),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1474),
.B(n_1443),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1441),
.B(n_1537),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1479),
.A2(n_1497),
.B(n_1482),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1519),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1507),
.B(n_1453),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1519),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1507),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1519),
.Y(n_1633)
);

OAI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1475),
.A2(n_1570),
.B(n_1557),
.C(n_1565),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1441),
.B(n_1505),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1449),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1459),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1535),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1560),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1566),
.A2(n_1574),
.B1(n_1444),
.B2(n_1447),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1507),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1455),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1501),
.A2(n_1567),
.B1(n_1499),
.B2(n_1578),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1474),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1438),
.A2(n_1475),
.B1(n_1454),
.B2(n_1473),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1485),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1505),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1556),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1512),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1487),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1476),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1512),
.Y(n_1652)
);

AOI222xp33_ASAP7_75t_L g1653 ( 
.A1(n_1451),
.A2(n_1554),
.B1(n_1445),
.B2(n_1492),
.C1(n_1457),
.C2(n_1472),
.Y(n_1653)
);

CKINVDCx6p67_ASAP7_75t_R g1654 ( 
.A(n_1542),
.Y(n_1654)
);

BUFx12f_ASAP7_75t_L g1655 ( 
.A(n_1564),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1481),
.A2(n_1463),
.B(n_1471),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1489),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1466),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1489),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1470),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1433),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1451),
.A2(n_1478),
.B(n_1464),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1561),
.Y(n_1663)
);

BUFx5_ASAP7_75t_L g1664 ( 
.A(n_1562),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1579),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1496),
.A2(n_1493),
.B1(n_1480),
.B2(n_1579),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1571),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1484),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1484),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1573),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1494),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1488),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1440),
.A2(n_1547),
.B1(n_1568),
.B2(n_1550),
.C(n_1439),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1562),
.B(n_1460),
.Y(n_1674)
);

AO21x1_ASAP7_75t_SL g1675 ( 
.A1(n_1552),
.A2(n_1468),
.B(n_1437),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1450),
.A2(n_1480),
.B1(n_1448),
.B2(n_1544),
.Y(n_1676)
);

INVx6_ASAP7_75t_L g1677 ( 
.A(n_1437),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1552),
.A2(n_1456),
.B(n_1455),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1552),
.A2(n_1456),
.B(n_1545),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1462),
.A2(n_1456),
.B(n_1469),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1437),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1546),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1546),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1546),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1576),
.B(n_1534),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1534),
.B(n_1540),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1448),
.A2(n_1577),
.B1(n_1538),
.B2(n_1563),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1435),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1442),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1435),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1446),
.A2(n_1575),
.B(n_1530),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1530),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1477),
.B(n_1575),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1434),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1434),
.Y(n_1695)
);

BUFx4f_ASAP7_75t_SL g1696 ( 
.A(n_1538),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1536),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1442),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1577),
.A2(n_1553),
.B1(n_1563),
.B2(n_1545),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1644),
.B(n_1536),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1582),
.A2(n_1605),
.B1(n_1612),
.B2(n_1645),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1639),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1607),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1623),
.A2(n_1442),
.B(n_1545),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1612),
.A2(n_1582),
.B(n_1634),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1595),
.B(n_1643),
.Y(n_1709)
);

OR2x6_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1691),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1640),
.A2(n_1627),
.B(n_1622),
.C(n_1653),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1626),
.B(n_1672),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1595),
.B(n_1648),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1622),
.A2(n_1608),
.B(n_1606),
.C(n_1613),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1595),
.B(n_1674),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1599),
.B(n_1600),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1672),
.B(n_1593),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1617),
.A2(n_1656),
.B(n_1608),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1593),
.B(n_1619),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_SL g1722 ( 
.A1(n_1666),
.A2(n_1673),
.B(n_1642),
.C(n_1601),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1617),
.A2(n_1656),
.B(n_1606),
.Y(n_1723)
);

AO32x2_ASAP7_75t_L g1724 ( 
.A1(n_1601),
.A2(n_1642),
.A3(n_1647),
.B1(n_1649),
.B2(n_1652),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1613),
.A2(n_1630),
.B(n_1635),
.C(n_1620),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1616),
.Y(n_1726)
);

BUFx12f_ASAP7_75t_L g1727 ( 
.A(n_1655),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1620),
.A2(n_1635),
.B1(n_1657),
.B2(n_1659),
.C(n_1652),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1597),
.A2(n_1623),
.B(n_1621),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1654),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1628),
.A2(n_1621),
.B(n_1617),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1630),
.A2(n_1628),
.B(n_1657),
.C(n_1659),
.Y(n_1732)
);

O2A1O1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1630),
.A2(n_1628),
.B(n_1632),
.C(n_1641),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1632),
.A2(n_1641),
.B(n_1581),
.C(n_1610),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1678),
.B(n_1636),
.Y(n_1735)
);

AOI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1649),
.A2(n_1647),
.B(n_1610),
.C(n_1615),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1691),
.B(n_1680),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1650),
.B(n_1651),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1695),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1654),
.B(n_1696),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1630),
.A2(n_1610),
.B1(n_1668),
.B2(n_1669),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1668),
.A2(n_1669),
.B1(n_1687),
.B2(n_1699),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1584),
.A2(n_1665),
.B(n_1624),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1638),
.B(n_1614),
.Y(n_1745)
);

AO32x2_ASAP7_75t_L g1746 ( 
.A1(n_1596),
.A2(n_1598),
.A3(n_1594),
.B1(n_1618),
.B2(n_1611),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1691),
.B(n_1680),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1668),
.A2(n_1669),
.B1(n_1676),
.B2(n_1615),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_SL g1749 ( 
.A1(n_1665),
.A2(n_1683),
.B(n_1580),
.C(n_1604),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_L g1750 ( 
.A(n_1667),
.B(n_1658),
.C(n_1660),
.D(n_1584),
.Y(n_1750)
);

AO32x2_ASAP7_75t_L g1751 ( 
.A1(n_1596),
.A2(n_1598),
.A3(n_1594),
.B1(n_1618),
.B2(n_1611),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1680),
.A2(n_1615),
.B1(n_1632),
.B2(n_1641),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1584),
.A2(n_1621),
.B1(n_1641),
.B2(n_1632),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1665),
.A2(n_1698),
.B(n_1689),
.C(n_1615),
.Y(n_1754)
);

BUFx4f_ASAP7_75t_SL g1755 ( 
.A(n_1689),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1583),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1615),
.A2(n_1664),
.B1(n_1689),
.B2(n_1698),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1609),
.B(n_1698),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1729),
.B(n_1625),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1711),
.A2(n_1625),
.B1(n_1629),
.B2(n_1631),
.C(n_1633),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1707),
.A2(n_1702),
.B1(n_1718),
.B2(n_1723),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1756),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1703),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1707),
.A2(n_1675),
.B1(n_1664),
.B2(n_1667),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1735),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1710),
.B(n_1633),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1747),
.B(n_1604),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1702),
.A2(n_1675),
.B1(n_1664),
.B2(n_1670),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1718),
.A2(n_1664),
.B1(n_1670),
.B2(n_1661),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1745),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1723),
.A2(n_1664),
.B1(n_1663),
.B2(n_1661),
.Y(n_1776)
);

AOI222xp33_ASAP7_75t_L g1777 ( 
.A1(n_1728),
.A2(n_1646),
.B1(n_1663),
.B2(n_1697),
.C1(n_1694),
.C2(n_1688),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1737),
.Y(n_1778)
);

INVx4_ASAP7_75t_L g1779 ( 
.A(n_1747),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1746),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1709),
.A2(n_1646),
.B1(n_1697),
.B2(n_1694),
.Y(n_1781)
);

NAND4xp25_ASAP7_75t_L g1782 ( 
.A(n_1731),
.B(n_1695),
.C(n_1692),
.D(n_1690),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1746),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.B(n_1588),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1751),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_1587),
.Y(n_1786)
);

NOR2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1750),
.B(n_1683),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1757),
.B(n_1760),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1751),
.B(n_1589),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1732),
.A2(n_1677),
.B1(n_1690),
.B2(n_1692),
.C(n_1684),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1753),
.B(n_1590),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1738),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1705),
.B(n_1585),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1771),
.B(n_1744),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1716),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1763),
.B(n_1752),
.Y(n_1796)
);

AOI33xp33_ASAP7_75t_L g1797 ( 
.A1(n_1763),
.A2(n_1725),
.A3(n_1722),
.B1(n_1736),
.B2(n_1733),
.B3(n_1721),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1785),
.B(n_1720),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1784),
.Y(n_1799)
);

INVx5_ASAP7_75t_SL g1800 ( 
.A(n_1771),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1784),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1764),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1784),
.Y(n_1803)
);

AO21x2_ASAP7_75t_L g1804 ( 
.A1(n_1791),
.A2(n_1753),
.B(n_1761),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1785),
.B(n_1712),
.Y(n_1805)
);

INVx5_ASAP7_75t_SL g1806 ( 
.A(n_1771),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1790),
.A2(n_1752),
.B1(n_1748),
.B2(n_1759),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1779),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1779),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1786),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1786),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1772),
.A2(n_1748),
.B1(n_1713),
.B2(n_1743),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1789),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1789),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1764),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1780),
.Y(n_1817)
);

OAI31xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1790),
.A2(n_1741),
.A3(n_1743),
.B(n_1750),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1791),
.B(n_1736),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1793),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1772),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1766),
.B(n_1724),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1764),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1708),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1779),
.B(n_1769),
.Y(n_1825)
);

AOI21xp33_ASAP7_75t_L g1826 ( 
.A1(n_1777),
.A2(n_1749),
.B(n_1741),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1765),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1775),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1792),
.B(n_1708),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1780),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1769),
.B(n_1724),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1820),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1795),
.B(n_1788),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1813),
.B(n_1778),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1822),
.B(n_1783),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1820),
.Y(n_1836)
);

AND2x2_ASAP7_75t_SL g1837 ( 
.A(n_1797),
.B(n_1774),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1813),
.B(n_1778),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1795),
.B(n_1788),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1813),
.B(n_1778),
.Y(n_1840)
);

BUFx10_ASAP7_75t_L g1841 ( 
.A(n_1802),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1813),
.B(n_1778),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1817),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1816),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1816),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1825),
.B(n_1779),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1801),
.B(n_1779),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1828),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1816),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1801),
.B(n_1779),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1821),
.B(n_1704),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1811),
.B(n_1769),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1821),
.B(n_1740),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1811),
.B(n_1768),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1820),
.Y(n_1856)
);

AO21x1_ASAP7_75t_SL g1857 ( 
.A1(n_1826),
.A2(n_1767),
.B(n_1773),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1823),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1812),
.B(n_1727),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1823),
.Y(n_1860)
);

NAND4xp25_ASAP7_75t_L g1861 ( 
.A(n_1797),
.B(n_1777),
.C(n_1762),
.D(n_1781),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1809),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1822),
.B(n_1783),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1828),
.Y(n_1864)
);

NOR2x1_ASAP7_75t_L g1865 ( 
.A(n_1819),
.B(n_1796),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1799),
.B(n_1770),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1825),
.B(n_1771),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1794),
.B(n_1771),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1799),
.B(n_1770),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1815),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1830),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1827),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1795),
.B(n_1788),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1803),
.B(n_1810),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1800),
.Y(n_1876)
);

OR2x6_ASAP7_75t_L g1877 ( 
.A(n_1865),
.B(n_1819),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1848),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1867),
.B(n_1800),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1835),
.B(n_1863),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1835),
.B(n_1798),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1837),
.B(n_1812),
.Y(n_1882)
);

NAND2x1_ASAP7_75t_L g1883 ( 
.A(n_1865),
.B(n_1831),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1841),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1867),
.B(n_1800),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1844),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1848),
.Y(n_1887)
);

INVx3_ASAP7_75t_R g1888 ( 
.A(n_1846),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1851),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1862),
.Y(n_1890)
);

AND3x2_ASAP7_75t_L g1891 ( 
.A(n_1859),
.B(n_1818),
.C(n_1809),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1841),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1845),
.Y(n_1894)
);

NAND2x1_ASAP7_75t_L g1895 ( 
.A(n_1867),
.B(n_1831),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1867),
.B(n_1800),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1837),
.B(n_1829),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1863),
.B(n_1798),
.Y(n_1899)
);

NAND2x1_ASAP7_75t_L g1900 ( 
.A(n_1846),
.B(n_1831),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1849),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1849),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1833),
.B(n_1798),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1841),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1858),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1838),
.B(n_1806),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1861),
.B(n_1829),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1833),
.B(n_1824),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1838),
.B(n_1806),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1838),
.B(n_1806),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1861),
.B(n_1818),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_R g1915 ( 
.A(n_1854),
.B(n_1726),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1841),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1847),
.A2(n_1807),
.B(n_1826),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

INVxp67_ASAP7_75t_SL g1919 ( 
.A(n_1862),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1839),
.B(n_1824),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1839),
.B(n_1824),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1877),
.B(n_1862),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1877),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1875),
.A2(n_1807),
.B1(n_1804),
.B2(n_1791),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1877),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1878),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1877),
.B(n_1868),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1890),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1883),
.B(n_1873),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_L g1930 ( 
.A(n_1914),
.B(n_1781),
.C(n_1762),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1898),
.B(n_1910),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1915),
.Y(n_1932)
);

AND2x4_ASAP7_75t_SL g1933 ( 
.A(n_1887),
.B(n_1846),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1886),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1882),
.B(n_1719),
.Y(n_1935)
);

INVx4_ASAP7_75t_L g1936 ( 
.A(n_1890),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1883),
.B(n_1880),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1889),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1903),
.B(n_1868),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1892),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1911),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1894),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1903),
.B(n_1868),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1917),
.B(n_1864),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1906),
.B(n_1868),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1896),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1891),
.B(n_1864),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1906),
.B(n_1868),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1880),
.B(n_1873),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1919),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1901),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1908),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1918),
.A2(n_1804),
.B1(n_1794),
.B2(n_1787),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1908),
.B(n_1840),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1876),
.B(n_1846),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1911),
.B(n_1815),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1909),
.B(n_1840),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1920),
.B(n_1815),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1926),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1950),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1924),
.A2(n_1895),
.B1(n_1900),
.B2(n_1734),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1936),
.B(n_1884),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1940),
.Y(n_1963)
);

OAI32xp33_ASAP7_75t_L g1964 ( 
.A1(n_1947),
.A2(n_1871),
.A3(n_1853),
.B1(n_1843),
.B2(n_1884),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_SL g1965 ( 
.A(n_1938),
.B(n_1900),
.C(n_1895),
.Y(n_1965)
);

AOI33xp33_ASAP7_75t_L g1966 ( 
.A1(n_1952),
.A2(n_1905),
.A3(n_1902),
.B1(n_1907),
.B2(n_1916),
.B3(n_1893),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1930),
.A2(n_1921),
.B1(n_1920),
.B2(n_1806),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1954),
.B(n_1909),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1936),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1954),
.B(n_1912),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1944),
.A2(n_1782),
.B1(n_1759),
.B2(n_1758),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1931),
.A2(n_1905),
.B(n_1893),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1938),
.A2(n_1857),
.B1(n_1804),
.B2(n_1913),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1932),
.Y(n_1974)
);

AOI21xp33_ASAP7_75t_L g1975 ( 
.A1(n_1923),
.A2(n_1916),
.B(n_1913),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1925),
.A2(n_1912),
.B(n_1879),
.Y(n_1976)
);

AOI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1928),
.A2(n_1885),
.B1(n_1876),
.B2(n_1897),
.C(n_1879),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_L g1978 ( 
.A(n_1936),
.B(n_1782),
.C(n_1904),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1941),
.B(n_1921),
.Y(n_1979)
);

INVx1_ASAP7_75t_SL g1980 ( 
.A(n_1933),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1940),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1934),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1953),
.A2(n_1804),
.B1(n_1885),
.B2(n_1897),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1935),
.A2(n_1853),
.B(n_1843),
.Y(n_1984)
);

AND2x4_ASAP7_75t_SL g1985 ( 
.A(n_1922),
.B(n_1846),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1960),
.Y(n_1986)
);

AOI321xp33_ASAP7_75t_L g1987 ( 
.A1(n_1964),
.A2(n_1928),
.A3(n_1927),
.B1(n_1941),
.B2(n_1922),
.C(n_1937),
.Y(n_1987)
);

NAND2x2_ASAP7_75t_L g1988 ( 
.A(n_1979),
.B(n_1937),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1959),
.Y(n_1989)
);

NAND3xp33_ASAP7_75t_L g1990 ( 
.A(n_1973),
.B(n_1922),
.C(n_1942),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1963),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1981),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1974),
.B(n_1957),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1969),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1983),
.A2(n_1929),
.B1(n_1949),
.B2(n_1927),
.Y(n_1995)
);

OAI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1973),
.A2(n_1957),
.B(n_1933),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1965),
.A2(n_1955),
.B1(n_1943),
.B2(n_1939),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1969),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1961),
.A2(n_1955),
.B1(n_1943),
.B2(n_1939),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1970),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1982),
.Y(n_2001)
);

NAND2x1_ASAP7_75t_L g2002 ( 
.A(n_1962),
.B(n_1955),
.Y(n_2002)
);

OAI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1980),
.A2(n_1929),
.B1(n_1949),
.B2(n_1948),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1971),
.A2(n_1804),
.B1(n_1946),
.B2(n_1951),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1978),
.B(n_1984),
.Y(n_2005)
);

OAI322xp33_ASAP7_75t_L g2006 ( 
.A1(n_1971),
.A2(n_1958),
.A3(n_1956),
.B1(n_1881),
.B2(n_1899),
.C1(n_1904),
.C2(n_1871),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1994),
.B(n_1966),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1993),
.B(n_1975),
.Y(n_2008)
);

NOR2xp67_ASAP7_75t_L g2009 ( 
.A(n_1997),
.B(n_1970),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1989),
.B(n_1976),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2000),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1998),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1986),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_2005),
.B(n_1972),
.Y(n_2014)
);

XNOR2xp5_ASAP7_75t_L g2015 ( 
.A(n_2003),
.B(n_1999),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_2002),
.B(n_1968),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1996),
.B(n_1966),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_L g2018 ( 
.A(n_1987),
.B(n_1977),
.C(n_1967),
.D(n_1948),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1990),
.B(n_1881),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2014),
.B(n_1995),
.C(n_2001),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2008),
.B(n_2010),
.Y(n_2021)
);

NOR3xp33_ASAP7_75t_L g2022 ( 
.A(n_2017),
.B(n_1992),
.C(n_1991),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_L g2023 ( 
.A(n_2018),
.B(n_2006),
.C(n_2004),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_2009),
.B(n_1985),
.Y(n_2024)
);

NAND4xp25_ASAP7_75t_L g2025 ( 
.A(n_2007),
.B(n_2004),
.C(n_1988),
.D(n_1945),
.Y(n_2025)
);

OAI211xp5_ASAP7_75t_SL g2026 ( 
.A1(n_2007),
.A2(n_1700),
.B(n_1958),
.C(n_1956),
.Y(n_2026)
);

AOI221x1_ASAP7_75t_L g2027 ( 
.A1(n_2012),
.A2(n_1945),
.B1(n_1888),
.B2(n_1730),
.C(n_1985),
.Y(n_2027)
);

NOR2x1_ASAP7_75t_L g2028 ( 
.A(n_2013),
.B(n_1847),
.Y(n_2028)
);

NOR3x1_ASAP7_75t_L g2029 ( 
.A(n_2011),
.B(n_2019),
.C(n_2015),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_SL g2030 ( 
.A1(n_2016),
.A2(n_1888),
.B1(n_1755),
.B2(n_1808),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_2019),
.B(n_1899),
.Y(n_2031)
);

NAND3xp33_ASAP7_75t_L g2032 ( 
.A(n_2014),
.B(n_1808),
.C(n_1847),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2023),
.B(n_1850),
.Y(n_2033)
);

NAND4xp25_ASAP7_75t_L g2034 ( 
.A(n_2029),
.B(n_1754),
.C(n_1808),
.D(n_1758),
.Y(n_2034)
);

NOR2xp67_ASAP7_75t_L g2035 ( 
.A(n_2024),
.B(n_2031),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_2020),
.A2(n_1808),
.B1(n_1809),
.B2(n_1794),
.Y(n_2036)
);

NAND4xp25_ASAP7_75t_L g2037 ( 
.A(n_2021),
.B(n_2025),
.C(n_2022),
.D(n_2027),
.Y(n_2037)
);

AOI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2026),
.A2(n_1850),
.B1(n_1870),
.B2(n_1840),
.C(n_1842),
.Y(n_2038)
);

AOI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_2037),
.A2(n_2032),
.B1(n_2030),
.B2(n_2028),
.C(n_1850),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2033),
.A2(n_1870),
.B(n_1715),
.Y(n_2040)
);

OAI31xp33_ASAP7_75t_L g2041 ( 
.A1(n_2034),
.A2(n_1787),
.A3(n_1842),
.B(n_1830),
.Y(n_2041)
);

AOI222xp33_ASAP7_75t_L g2042 ( 
.A1(n_2035),
.A2(n_1842),
.B1(n_1815),
.B2(n_1855),
.C1(n_1852),
.C2(n_1814),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_SL g2043 ( 
.A1(n_2036),
.A2(n_2038),
.B(n_1767),
.Y(n_2043)
);

OAI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2037),
.A2(n_1808),
.B1(n_1773),
.B2(n_1856),
.C(n_1836),
.Y(n_2044)
);

OAI211xp5_ASAP7_75t_SL g2045 ( 
.A1(n_2033),
.A2(n_1706),
.B(n_1739),
.C(n_1774),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2039),
.Y(n_2046)
);

XOR2xp5_ASAP7_75t_L g2047 ( 
.A(n_2040),
.B(n_1717),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2044),
.Y(n_2048)
);

BUFx3_ASAP7_75t_L g2049 ( 
.A(n_2041),
.Y(n_2049)
);

NOR2x1p5_ASAP7_75t_L g2050 ( 
.A(n_2043),
.B(n_1808),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2045),
.B(n_1858),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2046),
.A2(n_2042),
.B(n_1776),
.C(n_1805),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_1701),
.C(n_1686),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2049),
.B(n_1855),
.Y(n_2054)
);

AO22x2_ASAP7_75t_L g2055 ( 
.A1(n_2054),
.A2(n_2048),
.B1(n_2047),
.B2(n_2050),
.Y(n_2055)
);

AO22x2_ASAP7_75t_L g2056 ( 
.A1(n_2055),
.A2(n_2053),
.B1(n_2052),
.B2(n_2051),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2056),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2056),
.A2(n_1856),
.B1(n_1832),
.B2(n_1836),
.Y(n_2058)
);

AO22x2_ASAP7_75t_L g2059 ( 
.A1(n_2057),
.A2(n_1836),
.B1(n_1856),
.B2(n_1832),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2058),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2060),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2059),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2061),
.A2(n_1855),
.B1(n_1852),
.B2(n_1869),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2062),
.A2(n_1832),
.B(n_1872),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_2064),
.A2(n_1874),
.B(n_1852),
.Y(n_2065)
);

OAI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_2065),
.A2(n_2063),
.B1(n_1860),
.B2(n_1872),
.Y(n_2066)
);

OAI221xp5_ASAP7_75t_R g2067 ( 
.A1(n_2066),
.A2(n_1776),
.B1(n_1874),
.B2(n_1869),
.C(n_1866),
.Y(n_2067)
);

AOI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2067),
.A2(n_1685),
.B(n_1681),
.C(n_1682),
.Y(n_2068)
);


endmodule