module fake_netlist_1_9488_n_626 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_626);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_626;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g85 ( .A(n_46), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_32), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_68), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_50), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_70), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_53), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_44), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_48), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_49), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_77), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_2), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_14), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_27), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_9), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_55), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_61), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_82), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_23), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_20), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_51), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_12), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_65), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_5), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_74), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_7), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_58), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_24), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_75), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_28), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_108), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_89), .B(n_38), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_108), .B(n_1), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_128), .B(n_1), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_88), .B(n_2), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_90), .B(n_39), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_88), .B(n_3), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_92), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_122), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_94), .A2(n_3), .B(n_4), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_128), .B(n_5), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_101), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_131), .Y(n_157) );
AO22x2_ASAP7_75t_L g158 ( .A1(n_137), .A2(n_127), .B1(n_126), .B2(n_101), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_129), .B(n_100), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_129), .Y(n_160) );
NAND2xp33_ASAP7_75t_SL g161 ( .A(n_129), .B(n_95), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_140), .B(n_109), .Y(n_162) );
AND2x6_ASAP7_75t_L g163 ( .A(n_137), .B(n_114), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_137), .B(n_114), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_140), .B(n_96), .Y(n_165) );
INVxp67_ASAP7_75t_SL g166 ( .A(n_143), .Y(n_166) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_150), .B(n_115), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_143), .B(n_147), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_150), .B(n_115), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_137), .B(n_100), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_147), .B(n_127), .C(n_126), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_153), .B(n_123), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_137), .B(n_123), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_153), .B(n_97), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_150), .B(n_110), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_155), .B(n_98), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_155), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_159), .B(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_151), .B1(n_135), .B2(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_166), .B(n_145), .Y(n_195) );
NOR2x1p5_ASAP7_75t_L g196 ( .A(n_160), .B(n_103), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_159), .B(n_85), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_107), .B1(n_138), .B2(n_142), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_159), .B(n_151), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_169), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g202 ( .A1(n_181), .A2(n_102), .B1(n_120), .B2(n_124), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_166), .A2(n_151), .B(n_154), .C(n_152), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_187), .B(n_151), .Y(n_204) );
BUFx12f_ASAP7_75t_L g205 ( .A(n_181), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_158), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_162), .B(n_138), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_159), .B(n_142), .Y(n_209) );
BUFx4f_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_171), .B(n_136), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_187), .B(n_130), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_183), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_161), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_176), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_165), .B(n_130), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_130), .B(n_144), .C(n_133), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_177), .B(n_105), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_171), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_183), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
NOR2xp33_ASAP7_75t_R g231 ( .A(n_183), .B(n_119), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_190), .A2(n_134), .B(n_139), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_172), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_206), .B(n_178), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_230), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_232), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_209), .B(n_208), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_208), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_235), .B(n_165), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_232), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_180), .B1(n_163), .B2(n_164), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_205), .B(n_185), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_230), .B(n_177), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_206), .A2(n_112), .B1(n_179), .B2(n_186), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_230), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_235), .A2(n_177), .B(n_178), .C(n_179), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_205), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_236), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_199), .A2(n_164), .B1(n_163), .B2(n_180), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_194), .A2(n_163), .B1(n_180), .B2(n_164), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_207), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_197), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_209), .A2(n_164), .B1(n_163), .B2(n_180), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_209), .B(n_182), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_230), .B(n_177), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_197), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_209), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_210), .B(n_182), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
AO22x1_ASAP7_75t_L g265 ( .A1(n_233), .A2(n_163), .B1(n_180), .B2(n_164), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g266 ( .A1(n_202), .A2(n_116), .B1(n_113), .B2(n_186), .C(n_184), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_200), .B(n_164), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_195), .A2(n_191), .B(n_171), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_200), .B(n_164), .Y(n_269) );
AOI21xp33_ASAP7_75t_L g270 ( .A1(n_198), .A2(n_191), .B(n_171), .Y(n_270) );
INVxp67_ASAP7_75t_SL g271 ( .A(n_210), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_210), .Y(n_273) );
BUFx8_ASAP7_75t_L g274 ( .A(n_200), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_200), .B(n_164), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_194), .A2(n_184), .B1(n_167), .B2(n_175), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_192), .A2(n_180), .B1(n_134), .B2(n_139), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_225), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_SL g281 ( .A1(n_203), .A2(n_117), .B(n_136), .C(n_152), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_243), .A2(n_196), .B1(n_218), .B2(n_225), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g285 ( .A1(n_274), .A2(n_231), .B1(n_210), .B2(n_225), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_257), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_241), .B(n_237), .Y(n_287) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_244), .A2(n_196), .B1(n_225), .B2(n_221), .C1(n_204), .C2(n_121), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_257), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_180), .B1(n_234), .B2(n_222), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_251), .A2(n_278), .B(n_268), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_261), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_274), .Y(n_294) );
INVx8_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_255), .A2(n_213), .B1(n_220), .B2(n_228), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_255), .A2(n_228), .B1(n_214), .B2(n_211), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_253), .A2(n_180), .B1(n_234), .B2(n_217), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_252), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_244), .B(n_228), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_249), .B(n_237), .Y(n_301) );
AOI22xp33_ASAP7_75t_SL g302 ( .A1(n_274), .A2(n_139), .B1(n_134), .B2(n_167), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_262), .B(n_193), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_276), .B(n_193), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_256), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_248), .B(n_237), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_274), .A2(n_217), .B1(n_222), .B2(n_229), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_248), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_272), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_247), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_279), .B(n_201), .Y(n_313) );
CKINVDCx8_ASAP7_75t_R g314 ( .A(n_248), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_254), .A2(n_214), .B1(n_226), .B2(n_201), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_266), .A2(n_223), .B1(n_211), .B2(n_226), .C(n_215), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_259), .Y(n_318) );
BUFx8_ASAP7_75t_SL g319 ( .A(n_240), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_280), .A2(n_215), .B1(n_229), .B2(n_222), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_267), .B(n_217), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_288), .A2(n_260), .B1(n_269), .B2(n_275), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_300), .B(n_282), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_311), .A2(n_314), .B1(n_285), .B2(n_296), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_307), .A2(n_283), .B1(n_282), .B2(n_260), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_284), .A2(n_260), .B1(n_283), .B2(n_264), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_311), .B(n_264), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_310), .A2(n_260), .B1(n_264), .B2(n_134), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_310), .A2(n_139), .B1(n_134), .B2(n_258), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_300), .A2(n_277), .B1(n_278), .B2(n_238), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_307), .A2(n_238), .B1(n_273), .B2(n_250), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_318), .B(n_294), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_292), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_312), .A2(n_139), .B1(n_134), .B2(n_270), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_314), .A2(n_273), .B1(n_250), .B2(n_239), .Y(n_336) );
INVx5_ASAP7_75t_SL g337 ( .A(n_308), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_292), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_299), .A2(n_246), .B1(n_265), .B2(n_263), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_139), .B1(n_134), .B2(n_217), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_306), .B(n_222), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_293), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_321), .A2(n_139), .B1(n_134), .B2(n_239), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_295), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_301), .A2(n_265), .B(n_281), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
AOI222xp33_ASAP7_75t_L g348 ( .A1(n_306), .A2(n_121), .B1(n_110), .B2(n_111), .C1(n_118), .C2(n_122), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_313), .B(n_167), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_313), .A2(n_139), .B1(n_150), .B2(n_144), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_286), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_305), .B(n_136), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_333), .B(n_295), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_325), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_326), .A2(n_305), .B1(n_317), .B2(n_118), .C(n_111), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_325), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g357 ( .A1(n_324), .A2(n_297), .A3(n_315), .B(n_317), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_295), .B1(n_287), .B2(n_308), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_331), .A2(n_320), .B1(n_308), .B2(n_289), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_327), .A2(n_295), .B1(n_287), .B2(n_308), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_339), .B(n_289), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_345), .A2(n_295), .B1(n_287), .B2(n_308), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g363 ( .A(n_348), .B(n_340), .C(n_339), .D(n_343), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_345), .B(n_291), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_351), .Y(n_366) );
NAND3xp33_ASAP7_75t_L g367 ( .A(n_346), .B(n_302), .C(n_320), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_331), .A2(n_309), .B1(n_304), .B2(n_290), .C(n_298), .Y(n_368) );
OAI31xp33_ASAP7_75t_L g369 ( .A1(n_323), .A2(n_287), .A3(n_175), .B(n_149), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_328), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_334), .B(n_303), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_323), .B(n_349), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_349), .B(n_150), .Y(n_373) );
AOI33xp33_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_132), .A3(n_133), .B1(n_144), .B2(n_141), .B3(n_152), .Y(n_374) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_347), .A2(n_132), .B(n_133), .C(n_149), .Y(n_375) );
OAI221xp5_ASAP7_75t_SL g376 ( .A1(n_350), .A2(n_141), .B1(n_154), .B2(n_152), .C(n_149), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_345), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_328), .A2(n_303), .B1(n_150), .B2(n_175), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_334), .A2(n_106), .B(n_154), .C(n_141), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_337), .A2(n_139), .B1(n_132), .B2(n_154), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g382 ( .A1(n_338), .A2(n_332), .B1(n_350), .B2(n_352), .C1(n_336), .C2(n_342), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_355), .B(n_338), .C(n_122), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_337), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_366), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_370), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_370), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_377), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_337), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_365), .B(n_352), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_377), .B(n_303), .Y(n_392) );
AO21x2_ASAP7_75t_L g393 ( .A1(n_378), .A2(n_141), .B(n_149), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_366), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_356), .B(n_337), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_355), .A2(n_364), .B1(n_359), .B2(n_376), .C1(n_358), .C2(n_372), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_303), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_365), .B(n_329), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_366), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_372), .B(n_341), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_357), .A2(n_330), .B1(n_303), .B2(n_335), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_379), .B(n_6), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_357), .A2(n_344), .B1(n_104), .B2(n_146), .C(n_148), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_382), .A2(n_125), .B(n_156), .C(n_148), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_361), .B(n_148), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_379), .B(n_7), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_8), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_361), .B(n_148), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
OAI211xp5_ASAP7_75t_SL g414 ( .A1(n_353), .A2(n_148), .B(n_156), .C(n_188), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_363), .A2(n_156), .B(n_271), .C(n_239), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_377), .B(n_156), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_416), .B(n_364), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_410), .B(n_375), .C(n_380), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_401), .B(n_364), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_416), .B(n_364), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_418), .B(n_364), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_405), .B(n_373), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_418), .B(n_371), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_410), .A2(n_375), .A3(n_359), .B1(n_367), .B2(n_12), .B3(n_13), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_410), .B(n_397), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_388), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_367), .A3(n_10), .B1(n_11), .B2(n_13), .B3(n_15), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_389), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_389), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_407), .B(n_377), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_383), .A2(n_368), .B1(n_380), .B2(n_360), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g439 ( .A(n_407), .B(n_362), .C(n_369), .D(n_374), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_386), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_386), .B(n_373), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_388), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_387), .B(n_369), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_387), .B(n_8), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_10), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_385), .B(n_30), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_409), .B(n_368), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_398), .B(n_15), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_409), .B(n_376), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_409), .B(n_16), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_16), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
OAI31xp33_ASAP7_75t_SL g458 ( .A1(n_383), .A2(n_382), .A3(n_18), .B(n_19), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_417), .B(n_156), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_415), .A2(n_381), .B(n_212), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_396), .Y(n_462) );
OAI31xp33_ASAP7_75t_L g463 ( .A1(n_397), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_463) );
BUFx2_ASAP7_75t_SL g464 ( .A(n_385), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_396), .B(n_20), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_443), .B(n_392), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_423), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_429), .B(n_415), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_445), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_421), .Y(n_472) );
NAND2x1_ASAP7_75t_SL g473 ( .A(n_465), .B(n_417), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_419), .B(n_413), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_419), .B(n_413), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_455), .B(n_391), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_439), .A2(n_403), .B1(n_406), .B2(n_384), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_442), .B(n_391), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_457), .B(n_384), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_453), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_442), .B(n_384), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_457), .B(n_390), .Y(n_482) );
INVx4_ASAP7_75t_SL g483 ( .A(n_448), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_458), .A2(n_406), .B(n_392), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_461), .B(n_395), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_426), .B(n_395), .Y(n_488) );
BUFx2_ASAP7_75t_SL g489 ( .A(n_443), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_434), .A2(n_404), .B1(n_392), .B2(n_403), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_424), .B(n_413), .Y(n_491) );
NOR2x1p5_ASAP7_75t_L g492 ( .A(n_422), .B(n_393), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_427), .B(n_385), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_463), .A2(n_414), .B(n_392), .C(n_404), .Y(n_495) );
AOI32xp33_ASAP7_75t_L g496 ( .A1(n_420), .A2(n_414), .A3(n_400), .B1(n_394), .B2(n_24), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_424), .B(n_400), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_452), .B(n_393), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_435), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_430), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_437), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_449), .B(n_393), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_463), .A2(n_394), .B(n_393), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_440), .B(n_394), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_447), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_433), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_425), .B(n_21), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_456), .B(n_22), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_452), .A2(n_23), .B(n_25), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_25), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_478), .B(n_446), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_500), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_474), .B(n_425), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_471), .B(n_450), .Y(n_516) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_483), .B(n_462), .Y(n_517) );
AND4x1_ASAP7_75t_L g518 ( .A(n_511), .B(n_428), .C(n_431), .D(n_436), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_507), .B(n_444), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_469), .B(n_456), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_489), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_480), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_505), .A2(n_436), .B(n_422), .C(n_460), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g524 ( .A1(n_485), .A2(n_459), .B(n_462), .C(n_451), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_484), .Y(n_525) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_496), .A2(n_451), .B1(n_466), .B2(n_459), .C(n_464), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g527 ( .A(n_510), .B(n_466), .C(n_448), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_469), .A2(n_464), .B1(n_448), .B2(n_438), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_475), .B(n_448), .Y(n_529) );
XNOR2x2_ASAP7_75t_L g530 ( .A(n_498), .B(n_26), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_475), .B(n_31), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_491), .B(n_33), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_486), .B(n_34), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_494), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_499), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_35), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_481), .B(n_37), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_493), .B(n_41), .Y(n_539) );
AOI21xp33_ASAP7_75t_L g540 ( .A1(n_512), .A2(n_42), .B(n_43), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_470), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_SL g542 ( .A1(n_495), .A2(n_188), .B(n_174), .C(n_173), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_499), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
NAND2xp33_ASAP7_75t_R g547 ( .A(n_483), .B(n_47), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_483), .B(n_171), .Y(n_548) );
OAI32xp33_ASAP7_75t_L g549 ( .A1(n_486), .A2(n_490), .A3(n_467), .B1(n_503), .B2(n_501), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_477), .B(n_52), .Y(n_550) );
XOR2xp5_ASAP7_75t_L g551 ( .A(n_488), .B(n_54), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
AOI211xp5_ASAP7_75t_L g553 ( .A1(n_509), .A2(n_250), .B(n_245), .C(n_240), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_476), .A2(n_168), .B1(n_173), .B2(n_174), .C(n_188), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_472), .Y(n_556) );
O2A1O1Ixp5_ASAP7_75t_SL g557 ( .A1(n_467), .A2(n_56), .B(n_57), .C(n_59), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_497), .A2(n_245), .B1(n_240), .B2(n_242), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_495), .A2(n_242), .B(n_168), .C(n_64), .Y(n_559) );
OAI311xp33_ASAP7_75t_L g560 ( .A1(n_492), .A2(n_60), .A3(n_62), .B1(n_66), .C1(n_67), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_472), .A2(n_191), .B1(n_245), .B2(n_240), .C(n_250), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_508), .A2(n_191), .B1(n_245), .B2(n_240), .C(n_72), .Y(n_562) );
XOR2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_69), .Y(n_563) );
AOI211x1_ASAP7_75t_L g564 ( .A1(n_504), .A2(n_73), .B(n_76), .C(n_79), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_471), .B(n_80), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_505), .B(n_81), .C(n_83), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g567 ( .A1(n_505), .A2(n_84), .B(n_212), .C(n_216), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_505), .A2(n_212), .B1(n_216), .B2(n_227), .C(n_429), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_500), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_500), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_480), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_505), .A2(n_212), .B1(n_216), .B2(n_227), .C(n_458), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_505), .A2(n_227), .B(n_216), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_480), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_505), .A2(n_216), .B1(n_227), .B2(n_212), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_500), .B(n_212), .Y(n_576) );
OAI211xp5_ASAP7_75t_SL g577 ( .A1(n_496), .A2(n_227), .B(n_458), .C(n_463), .Y(n_577) );
NOR4xp75_ASAP7_75t_L g578 ( .A(n_572), .B(n_526), .C(n_548), .D(n_575), .Y(n_578) );
OAI22xp5_ASAP7_75t_SL g579 ( .A1(n_521), .A2(n_551), .B1(n_572), .B2(n_517), .Y(n_579) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_514), .B(n_524), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_520), .A2(n_569), .B1(n_568), .B2(n_549), .C1(n_570), .C2(n_523), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_520), .A2(n_566), .B1(n_577), .B2(n_519), .Y(n_582) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_573), .A2(n_568), .B(n_550), .C(n_527), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g584 ( .A1(n_550), .A2(n_547), .B(n_542), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_546), .B(n_545), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_541), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_556), .Y(n_587) );
AOI21xp33_ASAP7_75t_L g588 ( .A1(n_547), .A2(n_542), .B(n_567), .Y(n_588) );
INVxp33_ASAP7_75t_SL g589 ( .A(n_544), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_543), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_517), .A2(n_573), .B1(n_536), .B2(n_528), .Y(n_591) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_548), .B(n_536), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_536), .A2(n_553), .B1(n_538), .B2(n_516), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_563), .B(n_518), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_530), .A2(n_539), .B1(n_537), .B2(n_532), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_513), .B(n_552), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_539), .A2(n_532), .B1(n_531), .B2(n_537), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_533), .Y(n_598) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_579), .A2(n_559), .B(n_560), .C(n_533), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_590), .Y(n_600) );
AO22x2_ASAP7_75t_L g601 ( .A1(n_591), .A2(n_564), .B1(n_555), .B2(n_574), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_580), .B(n_515), .Y(n_602) );
NAND4xp75_ASAP7_75t_L g603 ( .A(n_582), .B(n_592), .C(n_584), .D(n_588), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_540), .B(n_531), .C(n_562), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g605 ( .A1(n_581), .A2(n_529), .B1(n_562), .B2(n_558), .C(n_565), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_595), .B(n_534), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_589), .A2(n_593), .B(n_583), .Y(n_607) );
NOR3x2_ASAP7_75t_L g608 ( .A(n_578), .B(n_557), .C(n_554), .Y(n_608) );
OAI22x1_ASAP7_75t_L g609 ( .A1(n_598), .A2(n_535), .B1(n_522), .B2(n_571), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_607), .B(n_593), .C(n_597), .D(n_576), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_603), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_601), .A2(n_585), .B1(n_586), .B2(n_587), .C(n_525), .Y(n_612) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_599), .B(n_561), .C(n_596), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_606), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_602), .B(n_529), .Y(n_615) );
OR4x2_ASAP7_75t_L g616 ( .A(n_613), .B(n_601), .C(n_605), .D(n_604), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_611), .B(n_608), .C(n_600), .Y(n_617) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_614), .Y(n_618) );
OR3x1_ASAP7_75t_L g619 ( .A(n_616), .B(n_610), .C(n_612), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_618), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_620), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_619), .A2(n_617), .B1(n_615), .B2(n_609), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_621), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_622), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_624), .B(n_619), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_625), .A2(n_620), .B(n_623), .Y(n_626) );
endmodule