module fake_jpeg_21283_n_75 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_55;
wire n_64;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_73;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_74;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_55)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_29),
.B1(n_38),
.B2(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_22),
.A2(n_24),
.B1(n_26),
.B2(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_44),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_23),
.C(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_59),
.C(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_59),
.B1(n_52),
.B2(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_35),
.B(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_32),
.C(n_28),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_34),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B(n_27),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_24),
.B(n_26),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_54),
.B(n_47),
.C(n_40),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_54),
.Y(n_75)
);


endmodule