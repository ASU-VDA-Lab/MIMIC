module fake_jpeg_3461_n_633 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_633);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_633;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_61),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_8),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_117),
.B(n_125),
.Y(n_147)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_66),
.Y(n_190)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_71),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_25),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_102),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_76),
.B(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_82),
.Y(n_179)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_84),
.Y(n_203)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_90),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_23),
.A2(n_7),
.B(n_16),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_111),
.B(n_0),
.Y(n_213)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_46),
.B(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_36),
.B(n_17),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_55),
.B(n_57),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_7),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_45),
.B1(n_50),
.B2(n_44),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_134),
.A2(n_175),
.B1(n_196),
.B2(n_0),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_54),
.B1(n_125),
.B2(n_65),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_148),
.A2(n_153),
.B(n_165),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_31),
.B1(n_56),
.B2(n_24),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_150),
.B(n_185),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_152),
.A2(n_166),
.B(n_168),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_62),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_50),
.B1(n_34),
.B2(n_53),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_34),
.B1(n_48),
.B2(n_36),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_61),
.B(n_57),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_171),
.B(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_59),
.B(n_24),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_206),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_69),
.A2(n_48),
.B1(n_56),
.B2(n_26),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_70),
.B(n_38),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_73),
.B(n_38),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_47),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_40),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_186),
.B(n_187),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_77),
.B(n_28),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_86),
.Y(n_192)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_123),
.A2(n_40),
.B1(n_31),
.B2(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_95),
.A2(n_34),
.B1(n_44),
.B2(n_26),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_99),
.B(n_28),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_15),
.Y(n_263)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_108),
.B(n_10),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_218),
.B(n_219),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_121),
.B(n_10),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_76),
.A2(n_55),
.B1(n_49),
.B2(n_42),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_16),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_223),
.A2(n_254),
.B1(n_176),
.B2(n_208),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_224),
.A2(n_232),
.B1(n_166),
.B2(n_220),
.Y(n_314)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_228),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_148),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_229),
.A2(n_248),
.B1(n_261),
.B2(n_283),
.Y(n_316)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_234),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_235),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_238),
.B(n_288),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_132),
.Y(n_239)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_240),
.Y(n_343)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVx3_ASAP7_75t_SL g340 ( 
.A(n_241),
.Y(n_340)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_187),
.B(n_3),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_243),
.Y(n_353)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_138),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_247),
.B(n_232),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_138),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_129),
.Y(n_249)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_168),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_254)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_260),
.A2(n_262),
.B1(n_264),
.B2(n_291),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_157),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_188),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g344 ( 
.A1(n_263),
.A2(n_270),
.B(n_299),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_194),
.A2(n_131),
.B1(n_162),
.B2(n_146),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_147),
.B(n_133),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_184),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_267),
.B(n_268),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_145),
.Y(n_269)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_147),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_164),
.Y(n_272)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_275),
.Y(n_324)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_181),
.Y(n_277)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_185),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_279),
.B(n_289),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_165),
.A2(n_153),
.B1(n_219),
.B2(n_209),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_200),
.Y(n_284)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_206),
.A2(n_205),
.B1(n_202),
.B2(n_169),
.Y(n_285)
);

AO22x1_ASAP7_75t_SL g339 ( 
.A1(n_285),
.A2(n_217),
.B1(n_203),
.B2(n_130),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_164),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_287),
.Y(n_309)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_178),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_141),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_136),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_197),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_294),
.B(n_295),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_199),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_137),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_298),
.Y(n_347)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_210),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_297),
.B(n_302),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_159),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_143),
.B(n_142),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_149),
.B(n_179),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_301),
.Y(n_356)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_195),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_210),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_160),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_327),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

OAI22x1_ASAP7_75t_SL g322 ( 
.A1(n_233),
.A2(n_158),
.B1(n_174),
.B2(n_161),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_242),
.B1(n_245),
.B2(n_298),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_248),
.B(n_182),
.CI(n_215),
.CON(n_325),
.SN(n_325)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_325),
.B(n_275),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_243),
.B(n_135),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_330),
.A2(n_338),
.B1(n_271),
.B2(n_280),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_243),
.B(n_176),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_339),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_229),
.A2(n_217),
.B1(n_204),
.B2(n_158),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_235),
.A2(n_203),
.B1(n_130),
.B2(n_139),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_270),
.B(n_139),
.C(n_286),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_352),
.C(n_249),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_231),
.B(n_139),
.C(n_278),
.Y(n_352)
);

AO22x1_ASAP7_75t_SL g354 ( 
.A1(n_285),
.A2(n_283),
.B1(n_227),
.B2(n_223),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_355),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_263),
.B(n_252),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_333),
.A2(n_227),
.B1(n_239),
.B2(n_237),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_373),
.B1(n_378),
.B2(n_323),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_316),
.A2(n_354),
.B1(n_345),
.B2(n_353),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_363),
.A2(n_365),
.B1(n_380),
.B2(n_407),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_316),
.A2(n_224),
.B1(n_237),
.B2(n_247),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_333),
.B(n_344),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_367),
.A2(n_374),
.B(n_404),
.Y(n_435)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_313),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_375),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_371),
.B(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_357),
.Y(n_372)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_372),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_309),
.A2(n_246),
.B1(n_236),
.B2(n_241),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_358),
.A2(n_264),
.B(n_262),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_359),
.Y(n_375)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_345),
.A2(n_226),
.B1(n_265),
.B2(n_281),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_306),
.Y(n_383)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_384),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_255),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_406),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_350),
.Y(n_410)
);

AO22x2_ASAP7_75t_SL g387 ( 
.A1(n_345),
.A2(n_253),
.B1(n_251),
.B2(n_291),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_388),
.Y(n_424)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_389),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_276),
.C(n_244),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_392),
.C(n_402),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_311),
.C(n_320),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_393),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_354),
.A2(n_322),
.B1(n_339),
.B2(n_327),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_394),
.A2(n_397),
.B1(n_400),
.B2(n_405),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_339),
.A2(n_228),
.B1(n_287),
.B2(n_272),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_399),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_314),
.B1(n_325),
.B2(n_335),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_305),
.B(n_256),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_401),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_258),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_324),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_323),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_329),
.A2(n_257),
.B(n_274),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_314),
.A2(n_284),
.B1(n_297),
.B2(n_302),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_260),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_319),
.A2(n_314),
.B1(n_307),
.B2(n_310),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_412),
.C(n_421),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_312),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_395),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_422),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_363),
.A2(n_307),
.B1(n_326),
.B2(n_340),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_426),
.B1(n_431),
.B2(n_389),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_392),
.B(n_390),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_404),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_368),
.A2(n_326),
.B1(n_340),
.B2(n_334),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_391),
.A2(n_303),
.B(n_360),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_427),
.A2(n_436),
.B(n_443),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_376),
.B(n_361),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_438),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_368),
.A2(n_303),
.B1(n_360),
.B2(n_321),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_377),
.A2(n_331),
.B1(n_321),
.B2(n_304),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_318),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_399),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_437),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_364),
.A2(n_310),
.B1(n_337),
.B2(n_318),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_442),
.A2(n_372),
.B1(n_381),
.B2(n_369),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_391),
.A2(n_341),
.B(n_304),
.Y(n_443)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_430),
.Y(n_448)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_446),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_451),
.B(n_454),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_422),
.A2(n_364),
.B(n_374),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_452),
.A2(n_457),
.B(n_463),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_408),
.Y(n_453)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_453),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_408),
.Y(n_454)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_435),
.A2(n_411),
.B(n_424),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_418),
.B(n_370),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_458),
.B(n_470),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_409),
.A2(n_394),
.B1(n_400),
.B2(n_397),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_459),
.A2(n_444),
.B1(n_439),
.B2(n_437),
.Y(n_516)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_461),
.Y(n_506)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_462),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_435),
.A2(n_377),
.B(n_405),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_385),
.Y(n_464)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_424),
.A2(n_406),
.B(n_365),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_465),
.A2(n_479),
.B(n_427),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_477),
.B1(n_478),
.B2(n_480),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_367),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_418),
.B(n_361),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_402),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_472),
.Y(n_500)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_414),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_473),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_414),
.B(n_382),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_474),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_383),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_410),
.C(n_443),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_425),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_476),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_428),
.A2(n_387),
.B1(n_403),
.B2(n_396),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_416),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_425),
.A2(n_393),
.B(n_387),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_428),
.A2(n_387),
.B1(n_398),
.B2(n_384),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_366),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_440),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_413),
.B(n_388),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_482),
.A2(n_460),
.B1(n_473),
.B2(n_462),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_468),
.A2(n_424),
.B1(n_413),
.B2(n_433),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_483),
.A2(n_491),
.B(n_504),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_459),
.A2(n_409),
.B1(n_433),
.B2(n_420),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_484),
.A2(n_485),
.B1(n_510),
.B2(n_516),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_465),
.A2(n_426),
.B1(n_412),
.B2(n_442),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_429),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_487),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_455),
.B(n_429),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_457),
.A2(n_465),
.B1(n_480),
.B2(n_477),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_493),
.A2(n_452),
.B1(n_469),
.B2(n_463),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_499),
.C(n_509),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_455),
.B(n_445),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_496),
.B(n_469),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_498),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_416),
.C(n_423),
.Y(n_499)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_434),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_448),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_452),
.A2(n_434),
.B(n_432),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_423),
.C(n_432),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_449),
.A2(n_444),
.B1(n_439),
.B2(n_417),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_454),
.C(n_453),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_520),
.C(n_543),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_449),
.C(n_460),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_521),
.B(n_530),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_510),
.Y(n_523)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_523),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_491),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_525),
.B(n_529),
.Y(n_560)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_526),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_527),
.B(n_534),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_505),
.A2(n_484),
.B1(n_503),
.B2(n_492),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_528),
.A2(n_493),
.B1(n_513),
.B2(n_500),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_532),
.Y(n_552)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_535),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_496),
.B(n_469),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_507),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_536),
.A2(n_539),
.B1(n_542),
.B2(n_485),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_495),
.B(n_447),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_519),
.Y(n_558)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_507),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_538),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_505),
.A2(n_476),
.B1(n_456),
.B2(n_447),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_490),
.A2(n_482),
.B1(n_470),
.B2(n_464),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_451),
.C(n_467),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_481),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_494),
.Y(n_553)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_545),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_542),
.A2(n_483),
.B1(n_492),
.B2(n_516),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_547),
.A2(n_524),
.B1(n_528),
.B2(n_536),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_517),
.B(n_502),
.C(n_514),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_549),
.B(n_550),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_517),
.B(n_489),
.C(n_511),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_529),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_561),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_553),
.B(n_558),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_525),
.A2(n_488),
.B(n_504),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_555),
.A2(n_540),
.B(n_467),
.Y(n_577)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_556),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_518),
.B(n_489),
.C(n_494),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_543),
.C(n_544),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_518),
.B(n_488),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_537),
.B(n_513),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_562),
.B(n_527),
.C(n_474),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_531),
.B1(n_458),
.B2(n_539),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_567),
.A2(n_568),
.B1(n_578),
.B2(n_564),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_556),
.A2(n_524),
.B1(n_515),
.B2(n_541),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_520),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_571),
.B(n_572),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_573),
.A2(n_561),
.B1(n_553),
.B2(n_550),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_522),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_566),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_577),
.A2(n_436),
.B(n_466),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_565),
.B(n_472),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_SL g579 ( 
.A(n_560),
.B(n_534),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_566),
.B(n_461),
.Y(n_595)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_552),
.Y(n_580)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_580),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_532),
.Y(n_582)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_582),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_548),
.A2(n_540),
.B1(n_466),
.B2(n_479),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_547),
.B1(n_560),
.B2(n_555),
.Y(n_585)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_584),
.B(n_549),
.C(n_574),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_585),
.B(n_595),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_546),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_588),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_570),
.A2(n_564),
.B1(n_554),
.B2(n_562),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_591),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_592),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_546),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_581),
.B(n_558),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_596),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_569),
.B(n_415),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_597),
.B(n_578),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_599),
.A2(n_577),
.B(n_582),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_603),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_594),
.B(n_591),
.Y(n_603)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_606),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_586),
.B(n_570),
.C(n_575),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_609),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_590),
.B(n_593),
.C(n_575),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_589),
.B(n_580),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_610),
.A2(n_587),
.B(n_585),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_598),
.A2(n_579),
.B(n_584),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_611),
.A2(n_608),
.B1(n_602),
.B2(n_508),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_612),
.B(n_614),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_573),
.C(n_599),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_601),
.C(n_609),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_615),
.A2(n_508),
.B(n_450),
.Y(n_621)
);

AO21x1_ASAP7_75t_SL g616 ( 
.A1(n_604),
.A2(n_583),
.B(n_478),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_616),
.A2(n_617),
.B(n_602),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_620),
.B(n_621),
.C(n_622),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_613),
.B(n_618),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_SL g627 ( 
.A(n_623),
.B(n_624),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_613),
.B(n_379),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_625),
.A2(n_626),
.B(n_349),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_622),
.B(n_619),
.C(n_616),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_629),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_627),
.A2(n_349),
.B(n_351),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_630),
.A2(n_351),
.B(n_343),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_332),
.C(n_328),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_332),
.B(n_328),
.Y(n_633)
);


endmodule