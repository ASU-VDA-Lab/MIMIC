module fake_jpeg_3295_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_51),
.B(n_46),
.C(n_49),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx12f_ASAP7_75t_SL g69 ( 
.A(n_59),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_54),
.B1(n_47),
.B2(n_50),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_0),
.Y(n_78)
);

OR2x4_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_60),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_54),
.B1(n_48),
.B2(n_50),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_87),
.B1(n_68),
.B2(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_55),
.B1(n_45),
.B2(n_41),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_41),
.B1(n_45),
.B2(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_93),
.Y(n_120)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_86),
.B1(n_79),
.B2(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_28),
.B1(n_37),
.B2(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_6),
.Y(n_117)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_25),
.C(n_38),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_26),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_119),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_27),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_126),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_109),
.C(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_17),
.B(n_34),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_14),
.B(n_32),
.C(n_31),
.D(n_30),
.Y(n_128)
);

OA21x2_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_129),
.B(n_120),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_11),
.B(n_39),
.C(n_9),
.D(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_115),
.B1(n_105),
.B2(n_112),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_134),
.B(n_138),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_132),
.B1(n_131),
.B2(n_124),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_137),
.C(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_141),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_124),
.B(n_123),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_148),
.A2(n_133),
.B(n_8),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_7),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_9),
.Y(n_151)
);


endmodule