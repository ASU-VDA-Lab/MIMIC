module fake_jpeg_26505_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_6),
.A2(n_15),
.B(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_21),
.A2(n_33),
.B1(n_18),
.B2(n_29),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_14),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_46),
.Y(n_66)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_18),
.B1(n_33),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_61),
.B1(n_71),
.B2(n_24),
.Y(n_91)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_18),
.B1(n_33),
.B2(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_65),
.Y(n_88)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_70),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_20),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_32),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_89),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_94),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_23),
.B(n_34),
.C(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_48),
.B(n_36),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_92),
.B1(n_70),
.B2(n_60),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_47),
.B1(n_27),
.B2(n_26),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_26),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_11),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_25),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_64),
.B1(n_55),
.B2(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_93),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_4),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_111),
.B1(n_123),
.B2(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_55),
.B1(n_52),
.B2(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_100),
.B1(n_80),
.B2(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_51),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2x1_ASAP7_75t_R g117 ( 
.A(n_88),
.B(n_1),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_85),
.B(n_86),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_2),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_76),
.B1(n_4),
.B2(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_120),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_137),
.B1(n_138),
.B2(n_104),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_117),
.C(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_86),
.C(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_142),
.B1(n_106),
.B2(n_122),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_96),
.B1(n_90),
.B2(n_80),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_79),
.B(n_101),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_138),
.B(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_113),
.B1(n_108),
.B2(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_97),
.B1(n_95),
.B2(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_97),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_150),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_112),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_7),
.B(n_8),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_134),
.C(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_149),
.C(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_143),
.B(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_174),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_137),
.C(n_144),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_143),
.B(n_150),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_166),
.C(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_180),
.Y(n_185)
);

OAI21x1_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_158),
.B(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_163),
.C(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_170),
.C(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_172),
.C(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_183),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_185),
.A3(n_155),
.B1(n_165),
.B2(n_9),
.C(n_106),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_165),
.C(n_9),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_191),
.Y(n_194)
);


endmodule