module fake_netlist_6_424_n_818 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_818);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_818;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_33),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_37),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_57),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_49),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_29),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_11),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_4),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_101),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_7),
.B(n_83),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_63),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_56),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_74),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_11),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_2),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_38),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_21),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_35),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_75),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_111),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_51),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_70),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_77),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_157),
.B(n_44),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_106),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_95),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_31),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_0),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_0),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_184),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_188),
.B(n_4),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_5),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_8),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_9),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_9),
.Y(n_262)
);

OAI22x1_ASAP7_75t_R g263 ( 
.A1(n_181),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_263)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_177),
.A2(n_10),
.B(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g272 ( 
.A(n_197),
.B(n_13),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_203),
.B(n_23),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_218),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_193),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_15),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_191),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

AO21x2_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_228),
.B(n_221),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_217),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_226),
.C(n_176),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_190),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_224),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_226),
.Y(n_296)
);

BUFx6f_ASAP7_75t_SL g297 ( 
.A(n_237),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_229),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_190),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_232),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_247),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

AND3x2_ASAP7_75t_L g306 ( 
.A(n_237),
.B(n_236),
.C(n_233),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_257),
.A2(n_212),
.B1(n_227),
.B2(n_225),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_250),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_253),
.B(n_175),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_241),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_251),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_243),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_256),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

AND3x2_ASAP7_75t_L g327 ( 
.A(n_253),
.B(n_16),
.C(n_17),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_272),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_248),
.B(n_183),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_262),
.B1(n_260),
.B2(n_254),
.C(n_274),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_269),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_269),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_331),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_280),
.Y(n_342)
);

NOR2x1p5_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_240),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_280),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_280),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_288),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_262),
.C(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_280),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_286),
.B(n_254),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_242),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_286),
.B(n_288),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_242),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_242),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

NOR2x1p5_ASAP7_75t_L g366 ( 
.A(n_297),
.B(n_249),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_303),
.Y(n_367)
);

O2A1O1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_304),
.A2(n_275),
.B(n_271),
.C(n_277),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_289),
.B(n_273),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_258),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_295),
.B(n_260),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_307),
.B(n_185),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_259),
.C(n_267),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_286),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_305),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_317),
.B(n_189),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_284),
.B(n_258),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_334),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_324),
.B(n_196),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_297),
.B(n_276),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_312),
.B(n_258),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_285),
.B(n_200),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_298),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_297),
.B(n_276),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_330),
.B(n_202),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_258),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_330),
.B(n_204),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_322),
.B(n_207),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_332),
.B(n_209),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_315),
.B(n_247),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_247),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_332),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_335),
.A2(n_351),
.B1(n_348),
.B2(n_343),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_299),
.B(n_319),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_397),
.A2(n_264),
.B1(n_248),
.B2(n_270),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_334),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_319),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_357),
.A2(n_299),
.B(n_328),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_264),
.B(n_279),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_374),
.A2(n_264),
.B1(n_279),
.B2(n_283),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_354),
.B(n_216),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_299),
.B(n_328),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_339),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_375),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_373),
.A2(n_316),
.B1(n_309),
.B2(n_311),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_372),
.A2(n_299),
.B(n_329),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_306),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_345),
.A2(n_299),
.B(n_329),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_337),
.A2(n_326),
.B(n_291),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_386),
.B(n_219),
.Y(n_427)
);

O2A1O1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_368),
.A2(n_311),
.B(n_309),
.C(n_321),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_327),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_386),
.B(n_222),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_380),
.A2(n_326),
.B(n_287),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_392),
.B(n_234),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_342),
.A2(n_291),
.B(n_287),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_399),
.A2(n_401),
.B(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

NOR2x1p5_ASAP7_75t_SL g444 ( 
.A(n_382),
.B(n_316),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_378),
.B(n_321),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_344),
.A2(n_276),
.B(n_263),
.C(n_247),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_369),
.A2(n_276),
.B(n_247),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_344),
.A2(n_338),
.B(n_392),
.C(n_352),
.Y(n_449)
);

O2A1O1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_393),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_398),
.A2(n_395),
.B(n_393),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_400),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_373),
.A2(n_97),
.B(n_172),
.Y(n_453)
);

AOI33xp33_ASAP7_75t_L g454 ( 
.A1(n_353),
.A2(n_19),
.A3(n_21),
.B1(n_24),
.B2(n_25),
.B3(n_26),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_395),
.A2(n_27),
.B(n_28),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_363),
.B(n_30),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_379),
.A2(n_32),
.B(n_36),
.C(n_40),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_379),
.B(n_41),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_336),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_350),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_364),
.A2(n_42),
.B(n_43),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_358),
.B(n_45),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_341),
.B(n_46),
.Y(n_463)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_355),
.A2(n_47),
.B(n_48),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_347),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_388),
.A2(n_50),
.B(n_52),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_394),
.A2(n_53),
.B(n_54),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_383),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_366),
.B(n_60),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_383),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_381),
.B(n_61),
.Y(n_472)
);

OAI21x1_ASAP7_75t_SL g473 ( 
.A1(n_453),
.A2(n_62),
.B(n_64),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_442),
.A2(n_391),
.B(n_360),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_411),
.A2(n_391),
.B(n_360),
.Y(n_475)
);

AOI21xp33_ASAP7_75t_L g476 ( 
.A1(n_403),
.A2(n_396),
.B(n_385),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_396),
.B1(n_385),
.B2(n_381),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_413),
.A2(n_391),
.B(n_69),
.C(n_71),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g479 ( 
.A1(n_403),
.A2(n_391),
.B(n_72),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_405),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_420),
.B(n_68),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

AOI21xp33_ASAP7_75t_L g484 ( 
.A1(n_431),
.A2(n_73),
.B(n_78),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_402),
.B(n_79),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_435),
.A2(n_80),
.B(n_81),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_410),
.B(n_82),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_406),
.Y(n_491)
);

AO21x1_ASAP7_75t_L g492 ( 
.A1(n_416),
.A2(n_453),
.B(n_409),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_84),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_408),
.A2(n_85),
.B(n_86),
.Y(n_496)
);

AO31x2_ASAP7_75t_L g497 ( 
.A1(n_416),
.A2(n_87),
.A3(n_88),
.B(n_89),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_438),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

NAND2x1_ASAP7_75t_L g501 ( 
.A(n_423),
.B(n_93),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_451),
.A2(n_94),
.B(n_98),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_100),
.B(n_102),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_450),
.A2(n_103),
.B(n_105),
.C(n_107),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_108),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_418),
.A2(n_173),
.B(n_113),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_422),
.A2(n_168),
.B(n_114),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_417),
.B(n_112),
.Y(n_510)
);

O2A1O1Ixp33_ASAP7_75t_SL g511 ( 
.A1(n_457),
.A2(n_115),
.B(n_116),
.C(n_118),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_121),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_439),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_425),
.A2(n_167),
.B(n_130),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_SL g518 ( 
.A(n_446),
.B(n_128),
.C(n_132),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_133),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_452),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_434),
.A2(n_134),
.B(n_135),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_413),
.A2(n_136),
.B(n_137),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_459),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_421),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_138),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_469),
.B(n_139),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_412),
.A2(n_141),
.B(n_142),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_520),
.A2(n_472),
.B(n_421),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_454),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_482),
.B(n_415),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_469),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_495),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_458),
.C(n_427),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_474),
.A2(n_472),
.B(n_463),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_517),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_475),
.A2(n_463),
.B(n_426),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_489),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_432),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_508),
.A2(n_456),
.B(n_466),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_500),
.Y(n_550)
);

INVx6_ASAP7_75t_L g551 ( 
.A(n_481),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_491),
.B(n_437),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_525),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_494),
.Y(n_554)
);

OAI21x1_ASAP7_75t_SL g555 ( 
.A1(n_473),
.A2(n_464),
.B(n_455),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_495),
.B(n_448),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g557 ( 
.A1(n_492),
.A2(n_440),
.B(n_447),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_519),
.B(n_461),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_476),
.A2(n_468),
.B(n_436),
.Y(n_559)
);

AOI22x1_ASAP7_75t_L g560 ( 
.A1(n_524),
.A2(n_428),
.B1(n_144),
.B2(n_145),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_485),
.A2(n_143),
.B(n_146),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_493),
.B(n_147),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_509),
.A2(n_148),
.B(n_149),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_496),
.A2(n_151),
.B(n_154),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_507),
.B(n_155),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_479),
.A2(n_158),
.B(n_160),
.Y(n_567)
);

OA21x2_ASAP7_75t_L g568 ( 
.A1(n_516),
.A2(n_162),
.B(n_163),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_495),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_519),
.A2(n_165),
.B(n_166),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_527),
.B(n_487),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_506),
.B(n_513),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_518),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_510),
.B(n_513),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_530),
.A2(n_477),
.B(n_488),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_503),
.A2(n_521),
.B(n_501),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_528),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_521),
.A2(n_504),
.B(n_523),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_538),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_577),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_525),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_541),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_561),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_573),
.A2(n_529),
.B1(n_527),
.B2(n_510),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_544),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_550),
.Y(n_588)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

CKINVDCx6p67_ASAP7_75t_R g591 ( 
.A(n_554),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_528),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_535),
.A2(n_514),
.B1(n_498),
.B2(n_484),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_553),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_573),
.A2(n_574),
.B1(n_572),
.B2(n_567),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_542),
.A2(n_478),
.B(n_497),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_551),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_497),
.B(n_487),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_548),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_497),
.B(n_487),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_552),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_567),
.A2(n_505),
.B(n_511),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_540),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_569),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_540),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_487),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_576),
.A2(n_487),
.B(n_519),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_543),
.A2(n_535),
.B1(n_546),
.B2(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_556),
.B(n_536),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_565),
.A2(n_578),
.B(n_539),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_577),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

AO21x1_ASAP7_75t_L g620 ( 
.A1(n_531),
.A2(n_562),
.B(n_563),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_535),
.B(n_536),
.Y(n_621)
);

AO21x2_ASAP7_75t_L g622 ( 
.A1(n_531),
.A2(n_555),
.B(n_547),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_580),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_610),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_580),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_560),
.B1(n_563),
.B2(n_566),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_587),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_590),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_602),
.B(n_534),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_590),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_621),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_617),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_617),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_604),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_611),
.B(n_534),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_551),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_613),
.B(n_551),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_621),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_579),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_595),
.A2(n_562),
.B1(n_559),
.B2(n_536),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_583),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_559),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_607),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_582),
.B(n_592),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_593),
.A2(n_558),
.B1(n_570),
.B2(n_568),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_599),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_609),
.B(n_568),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_570),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_588),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_599),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_621),
.B(n_568),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_596),
.B(n_558),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_600),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_621),
.B(n_592),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_607),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_584),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_589),
.B(n_615),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_618),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_594),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_610),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_622),
.Y(n_664)
);

AO31x2_ASAP7_75t_L g665 ( 
.A1(n_620),
.A2(n_597),
.A3(n_622),
.B(n_601),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_622),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_597),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_615),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_656),
.B(n_615),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_637),
.A2(n_591),
.B1(n_603),
.B2(n_619),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_628),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_635),
.B(n_605),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_608),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_630),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_643),
.B(n_598),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_643),
.B(n_646),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_635),
.B(n_591),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_646),
.B(n_598),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_671),
.B(n_631),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_629),
.B(n_614),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_623),
.B(n_581),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_638),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_630),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_623),
.B(n_581),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_632),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_671),
.B(n_581),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_626),
.B(n_618),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_633),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_633),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_658),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_648),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_625),
.B(n_618),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_625),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_659),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_644),
.B(n_618),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_606),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_629),
.B(n_606),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_634),
.B(n_645),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_644),
.B(n_651),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_686),
.B(n_667),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_689),
.B(n_653),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_699),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_681),
.B(n_680),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_690),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_702),
.B(n_634),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_709),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_690),
.Y(n_717)
);

AND2x6_ASAP7_75t_SL g718 ( 
.A(n_706),
.B(n_655),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_685),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_686),
.B(n_667),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_681),
.B(n_653),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_702),
.B(n_654),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_674),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_699),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_682),
.B(n_650),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_680),
.B(n_664),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_692),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_704),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_698),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_682),
.B(n_665),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_683),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_704),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_672),
.B(n_666),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_684),
.B(n_641),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_684),
.B(n_641),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_711),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_722),
.B(n_709),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_712),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_725),
.B(n_673),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_712),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_721),
.B(n_708),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_716),
.B(n_711),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_724),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_724),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_716),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_728),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_728),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_725),
.B(n_705),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_723),
.B(n_678),
.Y(n_749)
);

AOI21xp33_ASAP7_75t_L g750 ( 
.A1(n_739),
.A2(n_731),
.B(n_719),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_739),
.A2(n_725),
.B1(n_695),
.B2(n_705),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_689),
.B1(n_715),
.B2(n_735),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_749),
.B(n_721),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_748),
.A2(n_705),
.B1(n_711),
.B2(n_733),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_737),
.B(n_713),
.Y(n_756)
);

OAI21xp33_ASAP7_75t_L g757 ( 
.A1(n_741),
.A2(n_734),
.B(n_729),
.Y(n_757)
);

OAI33xp33_ASAP7_75t_L g758 ( 
.A1(n_738),
.A2(n_707),
.A3(n_730),
.B1(n_710),
.B2(n_720),
.B3(n_732),
.Y(n_758)
);

OAI21xp33_ASAP7_75t_L g759 ( 
.A1(n_741),
.A2(n_687),
.B(n_713),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_743),
.A2(n_730),
.B(n_705),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_751),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_752),
.A2(n_650),
.B1(n_736),
.B2(n_689),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_750),
.A2(n_718),
.B(n_742),
.C(n_745),
.Y(n_763)
);

OR4x1_ASAP7_75t_L g764 ( 
.A(n_758),
.B(n_747),
.C(n_744),
.D(n_732),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_753),
.A2(n_746),
.B1(n_740),
.B2(n_678),
.C(n_745),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_757),
.B1(n_759),
.B2(n_760),
.C(n_756),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_763),
.A2(n_755),
.B1(n_742),
.B2(n_672),
.Y(n_767)
);

AOI311xp33_ASAP7_75t_L g768 ( 
.A1(n_764),
.A2(n_718),
.A3(n_639),
.B(n_636),
.C(n_708),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_762),
.A2(n_754),
.B1(n_745),
.B2(n_746),
.C(n_640),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_761),
.B(n_703),
.Y(n_770)
);

OAI221xp5_ASAP7_75t_SL g771 ( 
.A1(n_763),
.A2(n_676),
.B1(n_710),
.B2(n_720),
.C(n_716),
.Y(n_771)
);

AOI322xp5_ASAP7_75t_L g772 ( 
.A1(n_766),
.A2(n_742),
.A3(n_726),
.B1(n_639),
.B2(n_703),
.C1(n_700),
.C2(n_714),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_771),
.B(n_660),
.C(n_663),
.Y(n_773)
);

AOI21xp33_ASAP7_75t_SL g774 ( 
.A1(n_767),
.A2(n_769),
.B(n_768),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_770),
.Y(n_775)
);

NAND4xp25_ASAP7_75t_L g776 ( 
.A(n_771),
.B(n_700),
.C(n_693),
.D(n_688),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_SL g777 ( 
.A(n_775),
.B(n_727),
.Y(n_777)
);

AO22x2_ASAP7_75t_L g778 ( 
.A1(n_773),
.A2(n_647),
.B1(n_693),
.B2(n_717),
.Y(n_778)
);

NOR3x1_ASAP7_75t_L g779 ( 
.A(n_776),
.B(n_694),
.C(n_675),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_779),
.B(n_774),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_SL g781 ( 
.A(n_778),
.B(n_772),
.C(n_660),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_777),
.B(n_660),
.C(n_663),
.Y(n_782)
);

XOR2xp5_ASAP7_75t_L g783 ( 
.A(n_780),
.B(n_669),
.Y(n_783)
);

NOR4xp25_ASAP7_75t_L g784 ( 
.A(n_781),
.B(n_661),
.C(n_663),
.D(n_651),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_782),
.Y(n_785)
);

AOI221xp5_ASAP7_75t_SL g786 ( 
.A1(n_780),
.A2(n_691),
.B1(n_688),
.B2(n_694),
.C(n_675),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_780),
.B(n_660),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_780),
.B(n_726),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_788),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_785),
.B(n_727),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_783),
.Y(n_792)
);

NAND4xp75_ASAP7_75t_L g793 ( 
.A(n_786),
.B(n_784),
.C(n_691),
.D(n_661),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_788),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_787),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_792),
.A2(n_794),
.B1(n_789),
.B2(n_790),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_795),
.A2(n_650),
.B(n_627),
.Y(n_797)
);

XNOR2x1_ASAP7_75t_L g798 ( 
.A(n_795),
.B(n_650),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_791),
.A2(n_714),
.B1(n_717),
.B2(n_649),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_791),
.B(n_627),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_798),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_796),
.B(n_793),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_800),
.B(n_677),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_797),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_799),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_SL g806 ( 
.A1(n_796),
.A2(n_642),
.B(n_677),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_802),
.A2(n_697),
.B1(n_679),
.B2(n_696),
.Y(n_807)
);

OAI21xp33_ASAP7_75t_L g808 ( 
.A1(n_801),
.A2(n_697),
.B(n_679),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_805),
.A2(n_696),
.B1(n_692),
.B2(n_701),
.Y(n_809)
);

AOI21xp33_ASAP7_75t_SL g810 ( 
.A1(n_804),
.A2(n_642),
.B(n_668),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_806),
.A2(n_668),
.B(n_652),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_807),
.A2(n_803),
.B1(n_701),
.B2(n_649),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_811),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_SL g814 ( 
.A1(n_813),
.A2(n_809),
.B1(n_808),
.B2(n_810),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_812),
.A2(n_664),
.B1(n_662),
.B2(n_624),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_815),
.A2(n_670),
.B(n_665),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_816),
.B(n_814),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_817),
.A2(n_624),
.B1(n_662),
.B2(n_670),
.Y(n_818)
);


endmodule