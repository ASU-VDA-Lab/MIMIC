module fake_jpeg_5807_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_45),
.B1(n_32),
.B2(n_34),
.Y(n_54)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_48),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_47),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_26),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_15),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_19),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_72),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_19),
.B1(n_16),
.B2(n_20),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_68),
.B1(n_28),
.B2(n_5),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_73),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_22),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_77),
.B(n_65),
.C(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_74),
.Y(n_92)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_33),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_31),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_31),
.B1(n_28),
.B2(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_0),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_41),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_103),
.Y(n_116)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_43),
.C(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_1),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_3),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_4),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_81),
.B1(n_80),
.B2(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_107),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_84),
.C(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_72),
.B1(n_57),
.B2(n_58),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_105),
.B1(n_86),
.B2(n_107),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_79),
.B(n_35),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_94),
.B(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_35),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_106),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_57),
.B1(n_4),
.B2(n_58),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_138),
.B(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_137),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_135),
.B1(n_144),
.B2(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_117),
.B1(n_114),
.B2(n_116),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_102),
.B(n_84),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_4),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_127),
.C(n_108),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_125),
.B1(n_121),
.B2(n_109),
.Y(n_145)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_153),
.C(n_157),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_110),
.B(n_124),
.C(n_120),
.D(n_112),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_156),
.A3(n_137),
.B1(n_142),
.B2(n_138),
.C1(n_130),
.C2(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_119),
.C(n_124),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_158),
.B1(n_135),
.B2(n_144),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_R g156 ( 
.A(n_144),
.B(n_70),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_89),
.C(n_115),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_136),
.B(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_141),
.Y(n_163)
);

XOR2x1_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_168),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_130),
.C(n_131),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_147),
.C(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_171),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_154),
.B1(n_158),
.B2(n_160),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_179),
.B(n_170),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_162),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.C(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_172),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_179),
.C(n_143),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule