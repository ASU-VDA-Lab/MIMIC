module fake_jpeg_14914_n_57 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_13),
.B1(n_1),
.B2(n_4),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_31),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_5),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI21x1_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_51),
.CON(n_52),
.SN(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_6),
.C(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_47),
.B1(n_11),
.B2(n_16),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_10),
.B1(n_17),
.B2(n_18),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_19),
.C(n_21),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_22),
.B(n_23),
.Y(n_57)
);


endmodule