module fake_jpeg_273_n_399 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_399);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_45),
.B(n_61),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_50),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_28),
.B(n_33),
.Y(n_104)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_3),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_76),
.Y(n_118)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_80),
.Y(n_96)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_35),
.B1(n_41),
.B2(n_39),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_99),
.B1(n_100),
.B2(n_116),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_25),
.B1(n_38),
.B2(n_27),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_78),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_38),
.B1(n_27),
.B2(n_21),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_38),
.B1(n_27),
.B2(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_59),
.B1(n_64),
.B2(n_62),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_77),
.B1(n_75),
.B2(n_68),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_104),
.A2(n_8),
.B(n_9),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_26),
.B1(n_36),
.B2(n_32),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_118),
.B(n_90),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_111),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_63),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_36),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_32),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_123),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_43),
.B(n_33),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_43),
.B(n_20),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_20),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_28),
.B1(n_20),
.B2(n_7),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_60),
.B1(n_54),
.B2(n_79),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_135),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_136),
.Y(n_226)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_168),
.B1(n_171),
.B2(n_111),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_161),
.Y(n_189)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_147),
.B(n_169),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_149),
.B(n_150),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_63),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_58),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_178),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_176),
.B1(n_133),
.B2(n_125),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_55),
.B1(n_44),
.B2(n_7),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_162),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_97),
.B(n_3),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_170),
.Y(n_209)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_167),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_118),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_173),
.Y(n_222)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_11),
.C(n_101),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_99),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_180),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_119),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_10),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_10),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_202),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_185),
.A2(n_194),
.B1(n_208),
.B2(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_98),
.B1(n_121),
.B2(n_89),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_191),
.B1(n_217),
.B2(n_156),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_98),
.B1(n_121),
.B2(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_192),
.B(n_189),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_138),
.A2(n_107),
.B1(n_130),
.B2(n_120),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_119),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_203),
.B(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_130),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_120),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_140),
.A2(n_124),
.B1(n_110),
.B2(n_126),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_142),
.B(n_110),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_171),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_144),
.A2(n_125),
.B1(n_126),
.B2(n_101),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_141),
.B(n_11),
.Y(n_219)
);

AOI22x1_ASAP7_75t_SL g224 ( 
.A1(n_157),
.A2(n_122),
.B1(n_127),
.B2(n_168),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_136),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_166),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_227),
.B(n_235),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_197),
.C(n_214),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_190),
.B1(n_185),
.B2(n_184),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_229),
.A2(n_240),
.B1(n_217),
.B2(n_191),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

AO21x2_ASAP7_75t_SL g233 ( 
.A1(n_190),
.A2(n_162),
.B(n_157),
.Y(n_233)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_233),
.A2(n_188),
.B1(n_162),
.B2(n_197),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_157),
.B(n_153),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_259),
.B(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_173),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_238),
.B(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_190),
.A2(n_162),
.B1(n_171),
.B2(n_152),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_170),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_248),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_253),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_197),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_137),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_228),
.Y(n_281)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_160),
.B(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_207),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_151),
.B(n_159),
.C(n_165),
.D(n_174),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_221),
.A3(n_211),
.B1(n_218),
.B2(n_219),
.C1(n_209),
.C2(n_214),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_249),
.B(n_261),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_234),
.B(n_229),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_266),
.A2(n_233),
.B(n_257),
.Y(n_299)
);

AOI22x1_ASAP7_75t_SL g269 ( 
.A1(n_233),
.A2(n_240),
.B1(n_232),
.B2(n_253),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_269),
.A2(n_271),
.B(n_275),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_270),
.A2(n_282),
.B1(n_293),
.B2(n_200),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_203),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_226),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_292),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_255),
.A2(n_198),
.B1(n_207),
.B2(n_205),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_223),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_285),
.B(n_288),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_201),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.C(n_294),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_193),
.C(n_201),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_244),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_198),
.B1(n_215),
.B2(n_158),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_195),
.C(n_216),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_266),
.A2(n_233),
.B1(n_243),
.B2(n_237),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_296),
.A2(n_304),
.B1(n_313),
.B2(n_289),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_307),
.B(n_265),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_248),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_273),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_249),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_310),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_242),
.C(n_246),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_303),
.C(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_231),
.C(n_236),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_245),
.B1(n_254),
.B2(n_239),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_312),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_260),
.C(n_251),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_282),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_250),
.C(n_256),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.C(n_292),
.Y(n_325)
);

OAI322xp33_ASAP7_75t_L g339 ( 
.A1(n_309),
.A2(n_284),
.A3(n_268),
.B1(n_274),
.B2(n_277),
.C1(n_275),
.C2(n_134),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_225),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_195),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_215),
.B1(n_200),
.B2(n_226),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_269),
.B1(n_289),
.B2(n_287),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_216),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_181),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_317),
.Y(n_327)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_278),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_134),
.B(n_213),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_275),
.B(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_272),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_324),
.B(n_337),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_333),
.C(n_336),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_331),
.B1(n_334),
.B2(n_338),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_329),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_300),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_311),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_267),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_289),
.B1(n_271),
.B2(n_293),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_272),
.C(n_278),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_291),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_296),
.A2(n_313),
.B1(n_305),
.B2(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_339),
.B(n_320),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_340),
.A2(n_316),
.B1(n_311),
.B2(n_318),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_307),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_356),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_307),
.B1(n_314),
.B2(n_297),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_275),
.B1(n_274),
.B2(n_213),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_295),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_277),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_330),
.Y(n_362)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_308),
.C(n_303),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_323),
.C(n_328),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_338),
.A2(n_297),
.B1(n_311),
.B2(n_310),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_354),
.A2(n_355),
.B1(n_335),
.B2(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_295),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_358),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_344),
.B1(n_352),
.B2(n_343),
.Y(n_373)
);

OAI221xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_356),
.B1(n_213),
.B2(n_134),
.C(n_127),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_357),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_363),
.B(n_364),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_333),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_365),
.B(n_122),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_329),
.C(n_332),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_368),
.C(n_372),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_353),
.C(n_349),
.Y(n_368)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_275),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_342),
.C(n_358),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_373),
.A2(n_371),
.B1(n_360),
.B2(n_361),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_346),
.Y(n_374)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_376),
.B(n_378),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_354),
.C(n_351),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_367),
.C(n_366),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_370),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_384),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_372),
.C(n_366),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_386),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_359),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_375),
.C(n_379),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_377),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_393),
.B(n_394),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_391),
.B(n_385),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_385),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_390),
.C(n_376),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_396),
.B(n_397),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_398),
.Y(n_399)
);


endmodule