module fake_jpeg_7584_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_21),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_15),
.CON(n_40),
.SN(n_40)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_59)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_24),
.B(n_20),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_22),
.C(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_60),
.B1(n_35),
.B2(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_30),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_17),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_20),
.B1(n_27),
.B2(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_27),
.B1(n_16),
.B2(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_74),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_18),
.B1(n_32),
.B2(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_77),
.B(n_78),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_19),
.B1(n_17),
.B2(n_44),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_82),
.B(n_87),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_47),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_95),
.C(n_31),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_91),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_90),
.B1(n_111),
.B2(n_67),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_35),
.B1(n_33),
.B2(n_25),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_47),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_46),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_105),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_25),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_115),
.Y(n_142)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_67),
.B1(n_66),
.B2(n_52),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_54),
.A2(n_33),
.B1(n_25),
.B2(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_26),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_15),
.B(n_11),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_86),
.B(n_97),
.C(n_78),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_91),
.B1(n_93),
.B2(n_109),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_144),
.B1(n_108),
.B2(n_107),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_83),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_56),
.C(n_48),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_137),
.C(n_138),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_82),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_10),
.B(n_15),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_139),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_80),
.B(n_14),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_56),
.C(n_61),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_52),
.B1(n_29),
.B2(n_33),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_94),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_151),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_143),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_155),
.B1(n_157),
.B2(n_160),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_163),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_88),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_98),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_177),
.B(n_145),
.Y(n_192)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_164),
.B1(n_121),
.B2(n_117),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_162),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_99),
.B1(n_113),
.B2(n_94),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_89),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_179),
.B1(n_160),
.B2(n_155),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_120),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_173),
.C(n_129),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_95),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_120),
.A2(n_95),
.B(n_101),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_109),
.B1(n_101),
.B2(n_102),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_122),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_177),
.B1(n_167),
.B2(n_171),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_142),
.B1(n_123),
.B2(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_182),
.A2(n_190),
.B1(n_201),
.B2(n_213),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_184),
.C(n_189),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_137),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_130),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_123),
.B1(n_132),
.B2(n_121),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_195),
.B(n_174),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_116),
.B(n_132),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_81),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_117),
.B1(n_116),
.B2(n_129),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.C(n_211),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_29),
.C(n_14),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_141),
.B(n_14),
.C(n_11),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_159),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_148),
.B(n_150),
.C(n_153),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_29),
.A3(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_141),
.B1(n_92),
.B2(n_81),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_153),
.B(n_165),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_230),
.B(n_185),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_220),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_180),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_188),
.B(n_152),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_147),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_225),
.C(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_237),
.B1(n_238),
.B2(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_163),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_235),
.B(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_154),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_158),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_171),
.C(n_170),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_151),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_195),
.A2(n_157),
.B(n_92),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_239),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_197),
.B(n_0),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_208),
.B1(n_210),
.B2(n_209),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_242),
.A2(n_244),
.B1(n_251),
.B2(n_256),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_235),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_209),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_247),
.B(n_222),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_191),
.B1(n_181),
.B2(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_228),
.B1(n_236),
.B2(n_214),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_214),
.A2(n_206),
.B1(n_212),
.B2(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_184),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_247),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_203),
.C(n_211),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_223),
.C(n_225),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_232),
.CI(n_226),
.CON(n_263),
.SN(n_263)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_261),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_252),
.B1(n_253),
.B2(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_226),
.C(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_189),
.C(n_234),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_275),
.B(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_230),
.B(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_248),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_237),
.C(n_238),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_279),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_2),
.C(n_3),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_3),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_298),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_245),
.B1(n_270),
.B2(n_242),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_257),
.B1(n_244),
.B2(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_295),
.B1(n_279),
.B2(n_254),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_243),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_257),
.B1(n_245),
.B2(n_248),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_251),
.B1(n_258),
.B2(n_263),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_281),
.B1(n_278),
.B2(n_280),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_300),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_294),
.B(n_249),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_254),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_268),
.C(n_269),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_286),
.B(n_266),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_312),
.B(n_288),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_295),
.B(n_293),
.C(n_292),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_319)
);

OAI221xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_296),
.B1(n_298),
.B2(n_291),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_300),
.B1(n_302),
.B2(n_311),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_297),
.B(n_299),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_319),
.B(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_323),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_285),
.B1(n_306),
.B2(n_7),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_327),
.C(n_328),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_285),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_313),
.B(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_8),
.C(n_318),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_8),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_330),
.A2(n_324),
.B(n_322),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_332),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_329),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_317),
.B(n_328),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_319),
.Y(n_339)
);


endmodule