module fake_jpeg_28872_n_448 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_17),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_57),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_82),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_16),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_16),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_34),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_95),
.B(n_100),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_132),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_109),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_34),
.B1(n_28),
.B2(n_20),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_41),
.B1(n_42),
.B2(n_40),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_113),
.B1(n_42),
.B2(n_70),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_42),
.B1(n_30),
.B2(n_40),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_30),
.B1(n_22),
.B2(n_40),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_127),
.B1(n_80),
.B2(n_78),
.Y(n_148)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_30),
.B1(n_44),
.B2(n_24),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_24),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_103),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_151),
.Y(n_179)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_27),
.B(n_38),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_33),
.C(n_111),
.Y(n_195)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_139),
.B1(n_110),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_65),
.B1(n_115),
.B2(n_93),
.Y(n_186)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_164),
.B1(n_178),
.B2(n_104),
.Y(n_197)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_159),
.Y(n_187)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_52),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_27),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_27),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_168),
.Y(n_194)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_27),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_170),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_173),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_96),
.B(n_77),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_175),
.Y(n_196)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_177),
.Y(n_198)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_20),
.C(n_38),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_92),
.B1(n_55),
.B2(n_59),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_92),
.B1(n_47),
.B2(n_53),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_173),
.B1(n_116),
.B2(n_93),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_205),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_154),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_116),
.B1(n_137),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_172),
.B1(n_167),
.B2(n_163),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_120),
.Y(n_202)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_133),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_213),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_180),
.B1(n_181),
.B2(n_189),
.Y(n_234)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g236 ( 
.A(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_154),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_216),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_215),
.A2(n_222),
.B(n_204),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_175),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_158),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_217),
.B(n_219),
.C(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_149),
.C(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_224),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_163),
.B1(n_144),
.B2(n_157),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_225),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_185),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_227),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_186),
.B(n_15),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_173),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_239),
.B1(n_254),
.B2(n_222),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_189),
.C(n_203),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_241),
.C(n_251),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_202),
.B1(n_192),
.B2(n_191),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_206),
.C(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_202),
.B1(n_107),
.B2(n_105),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_242),
.A2(n_211),
.B1(n_229),
.B2(n_231),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_207),
.B1(n_191),
.B2(n_188),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_212),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_212),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_206),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_191),
.B1(n_137),
.B2(n_136),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_213),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_204),
.B1(n_184),
.B2(n_182),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_236),
.B1(n_244),
.B2(n_226),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_254),
.B(n_256),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_260),
.B(n_261),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_262),
.B(n_282),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_209),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_264),
.A2(n_288),
.B1(n_263),
.B2(n_287),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_210),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_266),
.B(n_33),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_208),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_232),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_271),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_235),
.B(n_259),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_208),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_229),
.B1(n_220),
.B2(n_225),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_240),
.B(n_223),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_219),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_274),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_224),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_184),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_279),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_237),
.B(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_283),
.B1(n_287),
.B2(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_217),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_217),
.C(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_257),
.C(n_242),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_208),
.B1(n_226),
.B2(n_174),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_245),
.A2(n_226),
.B1(n_177),
.B2(n_162),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_257),
.B1(n_256),
.B2(n_235),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_309),
.B1(n_296),
.B2(n_305),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_289),
.Y(n_332)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_269),
.B(n_309),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_244),
.B(n_190),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_236),
.B1(n_248),
.B2(n_105),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_288),
.B1(n_264),
.B2(n_270),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_182),
.C(n_155),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_314),
.C(n_282),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_312),
.Y(n_336)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_146),
.C(n_152),
.Y(n_314)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_318),
.Y(n_333)
);

NOR4xp25_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_15),
.C(n_14),
.D(n_11),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_307),
.CI(n_286),
.CON(n_321),
.SN(n_321)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_292),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_321),
.B(n_341),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_323),
.A2(n_335),
.B1(n_293),
.B2(n_302),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_267),
.Y(n_325)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_331),
.C(n_342),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_263),
.Y(n_329)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_262),
.C(n_271),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_294),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_313),
.B1(n_304),
.B2(n_301),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_310),
.A2(n_289),
.B1(n_236),
.B2(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_119),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_340),
.B(n_316),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_15),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_199),
.C(n_119),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_343),
.B(n_318),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_297),
.C(n_317),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_365),
.C(n_367),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_354),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_351),
.A2(n_334),
.B1(n_349),
.B2(n_346),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_329),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_352),
.B(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_331),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_292),
.C(n_298),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_358),
.A2(n_344),
.B(n_320),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_339),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_295),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_361),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_324),
.A2(n_319),
.B1(n_304),
.B2(n_301),
.Y(n_363)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_199),
.C(n_111),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_9),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_138),
.C(n_129),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_369),
.A2(n_346),
.B1(n_372),
.B2(n_381),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_347),
.B(n_321),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_1),
.Y(n_400)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_321),
.C(n_344),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_374),
.A2(n_135),
.B1(n_124),
.B2(n_2),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_335),
.C(n_323),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_378),
.C(n_382),
.Y(n_391)
);

AO221x1_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_337),
.B1(n_326),
.B2(n_324),
.C(n_322),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_377),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_330),
.C(n_333),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_381),
.B(n_112),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_333),
.C(n_336),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_129),
.C(n_138),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_124),
.C(n_42),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_SL g384 ( 
.A(n_351),
.B(n_14),
.C(n_112),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_384),
.A2(n_0),
.B(n_1),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_385),
.B(n_362),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_357),
.B1(n_350),
.B2(n_355),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_389),
.A2(n_390),
.B1(n_386),
.B2(n_368),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_359),
.B1(n_367),
.B2(n_365),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_393),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_135),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_394),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_399),
.Y(n_414)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_398),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_1),
.Y(n_399)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_400),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_373),
.A2(n_1),
.B(n_2),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_401),
.B(n_371),
.Y(n_407)
);

INVx6_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_378),
.C(n_376),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_409),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_368),
.C(n_375),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_8),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_379),
.C(n_383),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_390),
.Y(n_418)
);

OA22x2_ASAP7_75t_L g412 ( 
.A1(n_387),
.A2(n_374),
.B1(n_380),
.B2(n_386),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_392),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_397),
.B1(n_401),
.B2(n_393),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_418),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_410),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_420),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_404),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_421),
.A2(n_422),
.B(n_425),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_396),
.C(n_4),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_3),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_424),
.C(n_414),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_3),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_421),
.B(n_413),
.Y(n_427)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_427),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_405),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_412),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_430),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_403),
.C(n_412),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_426),
.C(n_428),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_405),
.C(n_4),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_3),
.B(n_4),
.Y(n_434)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_434),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_438),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_430),
.A2(n_5),
.B(n_7),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_432),
.C(n_7),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_441),
.Y(n_444)
);

AO21x2_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_435),
.B(n_437),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_443),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_444),
.B(n_442),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_446),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_8),
.Y(n_448)
);


endmodule