module real_jpeg_25020_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_0),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_0),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_0),
.B(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_0),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_0),
.B(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_3),
.B(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_3),
.B(n_83),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_97),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_3),
.B(n_159),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_5),
.B(n_41),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_50),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_5),
.B(n_47),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_5),
.B(n_83),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_5),
.B(n_97),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_5),
.B(n_128),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_5),
.B(n_201),
.Y(n_371)
);

INVx8_ASAP7_75t_SL g129 ( 
.A(n_6),
.Y(n_129)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_50),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_7),
.B(n_83),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_7),
.B(n_97),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_7),
.B(n_201),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_8),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_9),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_9),
.B(n_47),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_83),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_97),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_9),
.B(n_222),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_74),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_11),
.B(n_50),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_47),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_11),
.B(n_83),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_11),
.B(n_97),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_11),
.B(n_128),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_11),
.B(n_201),
.Y(n_358)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_13),
.B(n_50),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_13),
.B(n_97),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_128),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_13),
.B(n_222),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_15),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_41),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_15),
.B(n_50),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_15),
.B(n_83),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_15),
.B(n_97),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_15),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_16),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_17),
.Y(n_116)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_376),
.B(n_377),
.C(n_381),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_367),
.C(n_375),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_352),
.C(n_353),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_329),
.C(n_330),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_299),
.C(n_300),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_274),
.C(n_275),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_243),
.C(n_244),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_205),
.C(n_206),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_166),
.C(n_167),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_133),
.C(n_134),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_109),
.C(n_110),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_88),
.C(n_89),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_66),
.C(n_67),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_52),
.C(n_57),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_46),
.C(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_41),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_60),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_65),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_72),
.C(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_74),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_77),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_87),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.C(n_87),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.C(n_100),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_95),
.C(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_103),
.C(n_104),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_108),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_125),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_126),
.C(n_132),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_120),
.C(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_119),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_121),
.Y(n_385)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.CI(n_124),
.CON(n_121),
.SN(n_121)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.CI(n_131),
.CON(n_126),
.SN(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_128),
.Y(n_217)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_149),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_138),
.C(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_145),
.C(n_148),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_140),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.CI(n_143),
.CON(n_140),
.SN(n_140)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_142),
.C(n_143),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_156),
.C(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B1(n_164),
.B2(n_165),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_192),
.C(n_193),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_162),
.C(n_163),
.Y(n_187)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_160),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_188),
.B2(n_204),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_189),
.C(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_172),
.C(n_181),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_181),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_177),
.C(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_175),
.B(n_228),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_186),
.C(n_187),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_228),
.Y(n_253)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_241),
.B2(n_242),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_232),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_232),
.C(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_219),
.C(n_220),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_210),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.CI(n_215),
.CON(n_210),
.SN(n_210)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_212),
.B(n_217),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_217),
.B(n_228),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_231),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_226),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_230),
.C(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_250),
.C(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_239),
.C(n_240),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_247),
.C(n_273),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_261),
.B2(n_273),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_256),
.C(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_254),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_SL g314 ( 
.A(n_253),
.B(n_279),
.C(n_282),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_257),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.CI(n_260),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_261),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.CI(n_264),
.CON(n_261),
.SN(n_261)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_272),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_269),
.A2(n_270),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_296),
.C(n_297),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_298),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_289),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_289),
.C(n_298),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_284),
.C(n_285),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_281),
.A2(n_282),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_SL g340 ( 
.A(n_282),
.B(n_307),
.C(n_309),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_285),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.CI(n_288),
.CON(n_285),
.SN(n_285)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_303),
.C(n_316),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_315),
.B2(n_316),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_311),
.B2(n_312),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_313),
.C(n_314),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_309),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_309),
.A2(n_310),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_346),
.C(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_319),
.C(n_322),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_325),
.C(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_327),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_330)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_333),
.C(n_351),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_340),
.C(n_341),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_354),
.C(n_356),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.CI(n_338),
.CON(n_335),
.SN(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_344),
.B1(n_347),
.B2(n_348),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_342),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_346),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_363),
.C(n_366),
.Y(n_369)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_369),
.C(n_370),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_359),
.CI(n_360),
.CON(n_357),
.SN(n_357)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_365),
.B2(n_366),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_364),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_SL g382 ( 
.A(n_364),
.B(n_371),
.C(n_374),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_365),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_373),
.A2(n_374),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_380),
.Y(n_381)
);


endmodule