module fake_ariane_1178_n_1697 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1697);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1697;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_15),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_25),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_119),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_96),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_3),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_49),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_88),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_29),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_99),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_18),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_35),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_23),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_69),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_67),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_27),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_42),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_58),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_27),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_133),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_55),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_59),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_77),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_56),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_14),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_40),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_141),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_60),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_53),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_80),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_5),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_75),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_48),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_13),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_15),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_45),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_18),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_52),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_36),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

INVx4_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_137),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_45),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_100),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_105),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_19),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_85),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_95),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_28),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_51),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_126),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_4),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_32),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_148),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_97),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_54),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_46),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_34),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_68),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_34),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_61),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_11),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_63),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_35),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_125),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_71),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_121),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_26),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_140),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_101),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_113),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_73),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_41),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_112),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_83),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_37),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_3),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_130),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_144),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_50),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_41),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_8),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_114),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_196),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_223),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_168),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_164),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_205),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_164),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_271),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_216),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_225),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_216),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_176),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_187),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_153),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_153),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_197),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_152),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_200),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_192),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_169),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_201),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_236),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_236),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_220),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_213),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_229),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_233),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_159),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_226),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_240),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_159),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_197),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_247),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_242),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_166),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_254),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_171),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_260),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_215),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_218),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_266),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_156),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_286),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_167),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_256),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_174),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_219),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_180),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_191),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_193),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_206),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_242),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_208),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_242),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_334),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_306),
.B(n_256),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_305),
.A2(n_243),
.B(n_228),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_157),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_307),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_326),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_341),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_224),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_340),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_188),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_310),
.A2(n_304),
.B(n_258),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_306),
.B(n_207),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_354),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_321),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_313),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_349),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_359),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_329),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_340),
.B(n_227),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_314),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_R g416 ( 
.A(n_323),
.B(n_171),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_341),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_338),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_261),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_344),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_154),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_368),
.B(n_154),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_337),
.B(n_151),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_182),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_361),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_337),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_322),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_377),
.B(n_294),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_315),
.B(n_246),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_325),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_362),
.B(n_182),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_371),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_327),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_375),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_327),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_368),
.B(n_210),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_316),
.B1(n_365),
.B2(n_324),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_R g456 ( 
.A(n_389),
.B(n_331),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_397),
.B(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_385),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_447),
.B(n_393),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_381),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_403),
.B(n_358),
.Y(n_461)
);

BUFx4f_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

CKINVDCx6p67_ASAP7_75t_R g464 ( 
.A(n_436),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_414),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_427),
.A2(n_378),
.B1(n_372),
.B2(n_376),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_410),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_377),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_373),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_410),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_312),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_380),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_418),
.B(n_332),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_406),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_379),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_427),
.B(n_373),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_SL g493 ( 
.A1(n_399),
.A2(n_320),
.B(n_318),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_424),
.B(n_277),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_438),
.A2(n_348),
.B1(n_351),
.B2(n_301),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_413),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_374),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_398),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_433),
.B(n_376),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_425),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_SL g505 ( 
.A1(n_420),
.A2(n_350),
.B(n_346),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_449),
.A2(n_378),
.B1(n_366),
.B2(n_352),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_386),
.A2(n_301),
.B1(n_172),
.B2(n_283),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_386),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_433),
.A2(n_303),
.B1(n_283),
.B2(n_172),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_442),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_424),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

AND3x2_ASAP7_75t_L g515 ( 
.A(n_433),
.B(n_352),
.C(n_333),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_422),
.B(n_434),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_388),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_424),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_422),
.B(n_151),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

CKINVDCx6p67_ASAP7_75t_R g525 ( 
.A(n_412),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_383),
.B(n_328),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_390),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_394),
.B(n_333),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_391),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_424),
.A2(n_367),
.B1(n_364),
.B2(n_363),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_383),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_417),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_383),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_405),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_417),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_434),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_444),
.B(n_328),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_405),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_444),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_425),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_429),
.B(n_330),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_404),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_416),
.A2(n_293),
.B1(n_185),
.B2(n_184),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_439),
.A2(n_281),
.B(n_279),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_425),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

AO21x2_ASAP7_75t_L g555 ( 
.A1(n_407),
.A2(n_297),
.B(n_288),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_384),
.A2(n_367),
.B1(n_364),
.B2(n_363),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_423),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_423),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_429),
.B(n_443),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_398),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_426),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_426),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_421),
.B(n_330),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_429),
.A2(n_178),
.B1(n_177),
.B2(n_184),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_SL g569 ( 
.A1(n_421),
.A2(n_360),
.B(n_357),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_425),
.Y(n_570)
);

AO22x2_ASAP7_75t_L g571 ( 
.A1(n_431),
.A2(n_437),
.B1(n_432),
.B2(n_440),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

AO21x2_ASAP7_75t_L g573 ( 
.A1(n_431),
.A2(n_298),
.B(n_357),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_446),
.B(n_155),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_395),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_435),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_435),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_446),
.B(n_155),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_446),
.B(n_160),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_446),
.B(n_160),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_392),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_448),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_409),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_419),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_419),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_419),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_384),
.A2(n_360),
.B(n_356),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_437),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_549),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_571),
.A2(n_384),
.B1(n_400),
.B2(n_441),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_505),
.A2(n_441),
.B1(n_440),
.B2(n_241),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_528),
.B(n_425),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_498),
.B(n_425),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_543),
.B(n_404),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_486),
.B(n_161),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_491),
.B(n_495),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_512),
.B(n_384),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_491),
.B(n_161),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_512),
.B(n_521),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_505),
.A2(n_241),
.B1(n_210),
.B2(n_300),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_495),
.B(n_162),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_479),
.B(n_237),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_585),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_502),
.B(n_536),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_585),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_513),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_513),
.B(n_162),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_490),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_566),
.A2(n_178),
.B1(n_293),
.B2(n_289),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_248),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_585),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_490),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_524),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_536),
.B(n_400),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_539),
.B(n_400),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_545),
.B(n_342),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_524),
.B(n_163),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_457),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_585),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_478),
.B(n_163),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_527),
.B(n_530),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_472),
.B(n_165),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_476),
.B(n_170),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_527),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_543),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_493),
.B(n_252),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_450),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_487),
.B(n_170),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_566),
.A2(n_285),
.B1(n_177),
.B2(n_185),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_453),
.B(n_259),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_530),
.B(n_175),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_450),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_500),
.B(n_179),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_461),
.B(n_289),
.C(n_291),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_532),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_474),
.B(n_262),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_550),
.B(n_291),
.C(n_285),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_571),
.A2(n_343),
.B1(n_356),
.B2(n_353),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_509),
.B(n_263),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_533),
.B(n_181),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_454),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_566),
.B(n_181),
.Y(n_657)
);

OR2x2_ASAP7_75t_SL g658 ( 
.A(n_492),
.B(n_411),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_509),
.B(n_265),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_566),
.B(n_183),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_566),
.B(n_183),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_533),
.B(n_186),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_545),
.B(n_303),
.C(n_275),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_549),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_550),
.B(n_295),
.C(n_278),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_571),
.A2(n_353),
.B1(n_347),
.B2(n_345),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_452),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_452),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_342),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_548),
.B(n_186),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_535),
.B(n_540),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_526),
.B(n_343),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_463),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_534),
.B(n_278),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_523),
.B(n_295),
.C(n_282),
.Y(n_675)
);

BUFx6f_ASAP7_75t_SL g676 ( 
.A(n_464),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_535),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_463),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_460),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_345),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_490),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_540),
.B(n_280),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_490),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_515),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_544),
.A2(n_280),
.B(n_300),
.Y(n_685)
);

BUFx8_ASAP7_75t_L g686 ( 
.A(n_525),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_468),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_282),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_460),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_544),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_587),
.B(n_588),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_587),
.B(n_284),
.Y(n_692)
);

BUFx8_ASAP7_75t_L g693 ( 
.A(n_525),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_547),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_468),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_586),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_588),
.B(n_589),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_589),
.B(n_284),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_586),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_547),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_569),
.B(n_287),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_526),
.B(n_459),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_569),
.B(n_490),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_542),
.B(n_456),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_451),
.B(n_317),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_590),
.B(n_287),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_542),
.B(n_317),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_455),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_526),
.B(n_0),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_590),
.B(n_296),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_591),
.B(n_296),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_484),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_560),
.B(n_1),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_1),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_506),
.B(n_189),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_594),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_594),
.B(n_5),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_571),
.A2(n_494),
.B1(n_573),
.B2(n_555),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_584),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_494),
.B(n_190),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_516),
.B(n_538),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_494),
.B(n_194),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_518),
.B(n_6),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_494),
.B(n_195),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_466),
.B(n_6),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_494),
.B(n_198),
.Y(n_728)
);

AOI21x1_ASAP7_75t_L g729 ( 
.A1(n_592),
.A2(n_231),
.B(n_274),
.Y(n_729)
);

INVxp33_ASAP7_75t_SL g730 ( 
.A(n_567),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_494),
.B(n_273),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_455),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_567),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_494),
.B(n_272),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_516),
.B(n_270),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_556),
.B(n_269),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_516),
.B(n_268),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_465),
.A2(n_267),
.B(n_264),
.C(n_255),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_516),
.B(n_538),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_465),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_516),
.B(n_253),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_593),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_573),
.A2(n_250),
.B1(n_249),
.B2(n_245),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_467),
.B(n_244),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_467),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_469),
.B(n_238),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_469),
.B(n_235),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_458),
.Y(n_748)
);

NAND2x1_ASAP7_75t_L g749 ( 
.A(n_466),
.B(n_81),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_538),
.B(n_232),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_462),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_458),
.B(n_480),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_497),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_573),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_508),
.B(n_230),
.C(n_221),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_748),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_679),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_699),
.B(n_592),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_604),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_751),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_612),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_613),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_650),
.B(n_510),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_680),
.B(n_538),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_751),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_617),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_730),
.A2(n_555),
.B1(n_552),
.B2(n_481),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_641),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_619),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_668),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_680),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_646),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_SL g773 ( 
.A(n_704),
.B(n_583),
.C(n_582),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_626),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_686),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_630),
.B(n_538),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_733),
.B(n_753),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_689),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_650),
.B(n_480),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_702),
.A2(n_581),
.B1(n_576),
.B2(n_496),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_639),
.B(n_466),
.Y(n_781)
);

AND2x6_ASAP7_75t_SL g782 ( 
.A(n_600),
.B(n_557),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_615),
.B(n_471),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_669),
.B(n_462),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_SL g785 ( 
.A(n_595),
.B(n_580),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_656),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_552),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_672),
.B(n_552),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_702),
.B(n_696),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_R g791 ( 
.A(n_676),
.B(n_473),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_621),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_686),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_632),
.B(n_555),
.Y(n_794)
);

BUFx4f_ASAP7_75t_L g795 ( 
.A(n_664),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_638),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_597),
.B(n_485),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_649),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_623),
.A2(n_580),
.B1(n_541),
.B2(n_537),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_707),
.B(n_499),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_634),
.B(n_485),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_712),
.B(n_485),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_653),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_668),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_693),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_677),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_729),
.A2(n_557),
.B(n_564),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_690),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_621),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_685),
.A2(n_496),
.B(n_475),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_609),
.A2(n_496),
.B1(n_578),
.B2(n_554),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_605),
.A2(n_470),
.B(n_475),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_694),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_693),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_623),
.A2(n_541),
.B1(n_507),
.B2(n_537),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_605),
.A2(n_470),
.B(n_482),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_640),
.A2(n_551),
.B1(n_519),
.B2(n_514),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_676),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_657),
.B(n_522),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_579),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_743),
.A2(n_719),
.B1(n_701),
.B2(n_705),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_621),
.B(n_501),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_708),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_732),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_700),
.B(n_579),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_611),
.B(n_499),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_611),
.B(n_499),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_740),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_551),
.B1(n_519),
.B2(n_514),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_625),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_732),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_673),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_625),
.B(n_501),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_R g836 ( 
.A(n_684),
.B(n_473),
.Y(n_836)
);

NOR2x2_ASAP7_75t_L g837 ( 
.A(n_709),
.B(n_482),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_658),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_SL g839 ( 
.A(n_723),
.B(n_483),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_644),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_654),
.B(n_531),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_725),
.B(n_477),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_601),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_678),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_603),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_651),
.B(n_665),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_SL g847 ( 
.A(n_622),
.B(n_199),
.C(n_202),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_675),
.B(n_554),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_654),
.B(n_578),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_745),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_687),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_602),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_695),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_660),
.B(n_522),
.Y(n_854)
);

AND2x6_ASAP7_75t_L g855 ( 
.A(n_606),
.B(n_483),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_644),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_742),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_659),
.B(n_554),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_659),
.B(n_563),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_714),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_602),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_716),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_607),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_718),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_652),
.B(n_578),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_607),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_652),
.B(n_666),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_625),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_720),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_614),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_477),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_625),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_616),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_666),
.B(n_563),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_635),
.A2(n_488),
.B(n_489),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_608),
.B(n_563),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_714),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_637),
.B(n_488),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_489),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_681),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_719),
.A2(n_529),
.B1(n_558),
.B2(n_572),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_681),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_SL g883 ( 
.A(n_643),
.B(n_631),
.C(n_662),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_635),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_642),
.B(n_562),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_671),
.A2(n_522),
.B(n_574),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_647),
.B(n_575),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_713),
.B(n_610),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_610),
.B(n_575),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_681),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_683),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_648),
.B(n_558),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_683),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_620),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_701),
.A2(n_529),
.B1(n_572),
.B2(n_507),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_683),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_661),
.B(n_501),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_671),
.Y(n_898)
);

INVx3_ASAP7_75t_SL g899 ( 
.A(n_618),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_663),
.B(n_568),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_624),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_633),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_691),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_697),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_752),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_628),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_717),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_717),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_703),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_599),
.A2(n_574),
.B(n_565),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_618),
.B(n_570),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_645),
.B(n_568),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_688),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_629),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_749),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_754),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_SL g917 ( 
.A(n_645),
.B(n_570),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_655),
.B(n_561),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_655),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_662),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_670),
.B(n_501),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_715),
.B(n_561),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_722),
.Y(n_923)
);

OAI22xp33_ASAP7_75t_L g924 ( 
.A1(n_636),
.A2(n_559),
.B1(n_501),
.B2(n_214),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_727),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_682),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_738),
.B(n_204),
.C(n_209),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_727),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_674),
.B(n_692),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_667),
.B(n_559),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_734),
.A2(n_546),
.B1(n_501),
.B2(n_217),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_779),
.A2(n_722),
.B(n_739),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_757),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_SL g934 ( 
.A(n_775),
.B(n_724),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_763),
.A2(n_736),
.B1(n_747),
.B2(n_746),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_812),
.A2(n_596),
.B(n_739),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_756),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_856),
.B(n_711),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_759),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_925),
.A2(n_596),
.B1(n_706),
.B2(n_698),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_777),
.B(n_710),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_805),
.B(n_726),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_795),
.B(n_721),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_903),
.B(n_598),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_795),
.B(n_728),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_819),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_777),
.A2(n_744),
.B1(n_731),
.B2(n_741),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_910),
.A2(n_750),
.B(n_737),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_840),
.A2(n_750),
.B(n_737),
.C(n_735),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_840),
.A2(n_735),
.B1(n_546),
.B2(n_212),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_862),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_926),
.B(n_211),
.Y(n_952)
);

O2A1O1Ixp5_ASAP7_75t_L g953 ( 
.A1(n_921),
.A2(n_553),
.B(n_503),
.C(n_11),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_910),
.A2(n_553),
.B(n_503),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_768),
.Y(n_955)
);

INVx3_ASAP7_75t_SL g956 ( 
.A(n_815),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_926),
.B(n_919),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_SL g958 ( 
.A1(n_907),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_819),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_793),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_771),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_761),
.Y(n_962)
);

OR2x6_ASAP7_75t_SL g963 ( 
.A(n_888),
.B(n_10),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_893),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_860),
.A2(n_877),
.B(n_907),
.C(n_908),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_790),
.B(n_13),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_772),
.Y(n_967)
);

AO32x2_ASAP7_75t_L g968 ( 
.A1(n_852),
.A2(n_863),
.A3(n_920),
.B1(n_866),
.B2(n_861),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_785),
.B(n_74),
.Y(n_969)
);

AO21x2_ASAP7_75t_L g970 ( 
.A1(n_807),
.A2(n_503),
.B(n_66),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_886),
.A2(n_62),
.B(n_138),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_771),
.B(n_14),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_928),
.A2(n_829),
.B(n_828),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_877),
.B(n_883),
.C(n_929),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_899),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_790),
.B(n_21),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_778),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_836),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_786),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_812),
.A2(n_22),
.B(n_24),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_762),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_891),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_SL g983 ( 
.A1(n_838),
.A2(n_899),
.B1(n_823),
.B2(n_846),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_841),
.A2(n_76),
.B(n_127),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_904),
.B(n_24),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_791),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_886),
.A2(n_57),
.B(n_118),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_849),
.A2(n_858),
.B(n_887),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_800),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_891),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_843),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_836),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_929),
.A2(n_28),
.B(n_30),
.C(n_33),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_R g994 ( 
.A(n_791),
.B(n_90),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_905),
.B(n_30),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_766),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_846),
.B(n_36),
.C(n_37),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_769),
.Y(n_998)
);

CKINVDCx11_ASAP7_75t_R g999 ( 
.A(n_782),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_774),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_867),
.B(n_884),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_913),
.B(n_38),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_898),
.B(n_47),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_813),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_822),
.B(n_47),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_845),
.B(n_98),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_813),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_883),
.A2(n_823),
.B1(n_802),
.B2(n_781),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_834),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_906),
.A2(n_885),
.B(n_878),
.Y(n_1010)
);

AOI33xp33_ASAP7_75t_L g1011 ( 
.A1(n_789),
.A2(n_803),
.A3(n_798),
.B1(n_796),
.B2(n_808),
.B3(n_806),
.Y(n_1011)
);

OAI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_842),
.A2(n_814),
.B1(n_850),
.B2(n_830),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_927),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_844),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_851),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_783),
.A2(n_784),
.B(n_820),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_914),
.B(n_909),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_787),
.B(n_788),
.Y(n_1018)
);

CKINVDCx10_ASAP7_75t_R g1019 ( 
.A(n_842),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_802),
.A2(n_781),
.B1(n_892),
.B2(n_900),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_770),
.B(n_804),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_792),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_760),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_794),
.B(n_865),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_892),
.A2(n_842),
.B1(n_764),
.B2(n_839),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_843),
.B(n_792),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_SL g1027 ( 
.A(n_847),
.B(n_773),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_927),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_889),
.A2(n_918),
.B(n_821),
.C(n_773),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_854),
.A2(n_801),
.B(n_875),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_874),
.B(n_864),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_817),
.A2(n_875),
.B(n_876),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_817),
.A2(n_810),
.B(n_911),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

NOR2xp67_ASAP7_75t_SL g1035 ( 
.A(n_792),
.B(n_832),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_897),
.A2(n_859),
.B(n_879),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_758),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_826),
.B(n_833),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_869),
.B(n_770),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_853),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_857),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_792),
.B(n_896),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_917),
.A2(n_827),
.B(n_824),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_824),
.A2(n_835),
.B(n_776),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_760),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_813),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_L g1047 ( 
.A(n_804),
.B(n_825),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_767),
.A2(n_811),
.B1(n_780),
.B2(n_931),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_767),
.B(n_833),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_835),
.A2(n_912),
.B(n_797),
.C(n_765),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_826),
.B(n_901),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_811),
.A2(n_879),
.B1(n_799),
.B2(n_918),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_923),
.A2(n_848),
.B(n_765),
.C(n_895),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_871),
.B(n_894),
.Y(n_1054)
);

CKINVDCx8_ASAP7_75t_R g1055 ( 
.A(n_880),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_879),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_870),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_809),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_895),
.A2(n_915),
.B(n_799),
.C(n_816),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_871),
.A2(n_924),
.B(n_873),
.C(n_902),
.Y(n_1060)
);

BUFx8_ASAP7_75t_SL g1061 ( 
.A(n_813),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_930),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_816),
.A2(n_818),
.B(n_831),
.C(n_930),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_831),
.B(n_922),
.C(n_881),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_868),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_868),
.A2(n_872),
.B(n_882),
.Y(n_1066)
);

BUFx10_ASAP7_75t_L g1067 ( 
.A(n_946),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_941),
.B(n_832),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_973),
.A2(n_896),
.B(n_890),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1032),
.A2(n_881),
.B(n_916),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1029),
.A2(n_855),
.B(n_922),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1011),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_938),
.B(n_890),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_940),
.A2(n_974),
.B(n_1008),
.Y(n_1074)
);

AOI221xp5_ASAP7_75t_L g1075 ( 
.A1(n_940),
.A2(n_837),
.B1(n_868),
.B2(n_872),
.C(n_882),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_982),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1020),
.B(n_890),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_939),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1030),
.A2(n_855),
.B(n_896),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_948),
.A2(n_855),
.B(n_872),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_962),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_959),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_961),
.B(n_882),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1010),
.A2(n_1018),
.B(n_932),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_SL g1085 ( 
.A(n_997),
.B(n_1028),
.C(n_1013),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1012),
.B(n_965),
.Y(n_1086)
);

INVx8_ASAP7_75t_L g1087 ( 
.A(n_1061),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_1018),
.A2(n_1048),
.A3(n_1024),
.B(n_1052),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1052),
.A2(n_985),
.B1(n_1048),
.B2(n_963),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_933),
.B(n_989),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_993),
.B(n_1027),
.C(n_986),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_989),
.B(n_1001),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_985),
.A2(n_1063),
.B1(n_980),
.B2(n_976),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1001),
.B(n_966),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_1005),
.B(n_1056),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_999),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_981),
.B(n_996),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_971),
.A2(n_987),
.B(n_1016),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1043),
.A2(n_936),
.B(n_1036),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_982),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_983),
.A2(n_1064),
.B1(n_937),
.B2(n_1062),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_998),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_954),
.A2(n_1044),
.B(n_1066),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1000),
.B(n_1031),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_978),
.B(n_992),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1055),
.B(n_990),
.Y(n_1106)
);

NAND3x1_ASAP7_75t_L g1107 ( 
.A(n_1025),
.B(n_980),
.C(n_972),
.Y(n_1107)
);

AO32x2_ASAP7_75t_L g1108 ( 
.A1(n_968),
.A2(n_1049),
.A3(n_1058),
.B1(n_1022),
.B2(n_958),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_1024),
.A2(n_1049),
.A3(n_1059),
.B(n_1053),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_949),
.A2(n_935),
.B(n_1060),
.C(n_947),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_957),
.A2(n_1002),
.B1(n_975),
.B2(n_995),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_977),
.B(n_1034),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_951),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1050),
.A2(n_944),
.B(n_984),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1031),
.B(n_1017),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_955),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_952),
.A2(n_1003),
.B(n_995),
.C(n_943),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1017),
.B(n_1051),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_944),
.A2(n_1003),
.B(n_953),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1039),
.B(n_1038),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1037),
.A2(n_945),
.B(n_1042),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1041),
.B(n_1054),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_967),
.B(n_1014),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_990),
.B(n_1021),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_979),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1009),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1015),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1006),
.A2(n_950),
.B(n_934),
.C(n_1047),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_990),
.B(n_1026),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1057),
.A2(n_1040),
.A3(n_970),
.B(n_968),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_964),
.B(n_960),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_968),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_964),
.B(n_942),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_964),
.B(n_1023),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_970),
.A2(n_1065),
.A3(n_1046),
.B(n_1004),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1004),
.A2(n_1065),
.A3(n_1046),
.B(n_1007),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1045),
.B(n_1065),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1004),
.B(n_1007),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_994),
.B(n_1035),
.C(n_1007),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1046),
.B(n_969),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1019),
.A2(n_763),
.B(n_650),
.C(n_974),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_R g1142 ( 
.A(n_969),
.B(n_542),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1018),
.A2(n_1059),
.B(n_779),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_938),
.B(n_730),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1032),
.A2(n_1030),
.B(n_807),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1029),
.A2(n_763),
.B(n_940),
.Y(n_1146)
);

NOR2xp67_ASAP7_75t_L g1147 ( 
.A(n_933),
.B(n_689),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_941),
.A2(n_925),
.B1(n_763),
.B2(n_877),
.Y(n_1148)
);

INVx4_ASAP7_75t_SL g1149 ( 
.A(n_956),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1048),
.A2(n_1052),
.B1(n_940),
.B2(n_1018),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_974),
.A2(n_763),
.B(n_650),
.C(n_840),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_982),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1033),
.A2(n_807),
.B(n_1032),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1032),
.A2(n_1030),
.B(n_807),
.Y(n_1154)
);

NOR2x1_ASAP7_75t_L g1155 ( 
.A(n_991),
.B(n_775),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_938),
.B(n_777),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1033),
.A2(n_807),
.B(n_1032),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1029),
.A2(n_763),
.B(n_940),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_1030),
.B(n_807),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1029),
.A2(n_763),
.B(n_940),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_938),
.B(n_730),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_974),
.A2(n_763),
.B(n_650),
.C(n_840),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_938),
.B(n_730),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1032),
.A2(n_1033),
.B(n_1030),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1018),
.A2(n_1059),
.B(n_779),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_1022),
.B(n_1058),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1018),
.B(n_867),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_991),
.B(n_771),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1029),
.A2(n_763),
.B(n_940),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1011),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_938),
.B(n_777),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1022),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_951),
.Y(n_1173)
);

AOI221x1_ASAP7_75t_L g1174 ( 
.A1(n_997),
.A2(n_980),
.B1(n_1048),
.B2(n_940),
.C(n_1029),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1048),
.B(n_730),
.Y(n_1175)
);

AOI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1048),
.A2(n_763),
.B(n_1052),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_938),
.B(n_777),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_938),
.B(n_777),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1018),
.A2(n_1059),
.B(n_779),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_933),
.Y(n_1180)
);

AO21x1_ASAP7_75t_L g1181 ( 
.A1(n_1048),
.A2(n_940),
.B(n_1052),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_938),
.B(n_777),
.Y(n_1182)
);

CKINVDCx14_ASAP7_75t_R g1183 ( 
.A(n_959),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_933),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_941),
.B(n_856),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_946),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1018),
.A2(n_1048),
.A3(n_1024),
.B(n_1010),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_988),
.A2(n_973),
.B(n_779),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1032),
.A2(n_1030),
.B(n_807),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1097),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1090),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1167),
.B(n_1115),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1078),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1130),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1189),
.A2(n_1098),
.B(n_1103),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1156),
.A2(n_1182),
.B1(n_1177),
.B2(n_1171),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1081),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1086),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1186),
.Y(n_1200)
);

NAND3x1_ASAP7_75t_L g1201 ( 
.A(n_1144),
.B(n_1163),
.C(n_1161),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1167),
.B(n_1088),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1178),
.A2(n_1151),
.B1(n_1162),
.B2(n_1141),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1102),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1176),
.A2(n_1146),
.B(n_1158),
.C(n_1169),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1181),
.A2(n_1174),
.A3(n_1089),
.B(n_1084),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1105),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1130),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1113),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1087),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1080),
.A2(n_1114),
.B(n_1079),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1099),
.A2(n_1070),
.B(n_1188),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_1087),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1130),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1175),
.A2(n_1089),
.B1(n_1176),
.B2(n_1160),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1148),
.A2(n_1074),
.B1(n_1160),
.B2(n_1146),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1095),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1126),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1158),
.A2(n_1169),
.B(n_1148),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1127),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1074),
.A2(n_1175),
.B(n_1119),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1164),
.Y(n_1222)
);

AOI332xp33_ASAP7_75t_L g1223 ( 
.A1(n_1111),
.A2(n_1170),
.A3(n_1072),
.B1(n_1112),
.B2(n_1094),
.B3(n_1120),
.C1(n_1118),
.C2(n_1132),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1136),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1119),
.A2(n_1117),
.B(n_1165),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1092),
.B(n_1104),
.Y(n_1226)
);

NAND2x1_ASAP7_75t_L g1227 ( 
.A(n_1143),
.B(n_1179),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1173),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1093),
.A2(n_1110),
.B(n_1111),
.C(n_1075),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1093),
.A2(n_1185),
.B1(n_1150),
.B2(n_1073),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1123),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1088),
.B(n_1150),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1168),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1121),
.A2(n_1128),
.B(n_1068),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1100),
.B(n_1129),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_1096),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1082),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1129),
.B(n_1139),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1139),
.B(n_1083),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1124),
.B(n_1106),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1085),
.B(n_1133),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1142),
.B(n_1184),
.C(n_1180),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1137),
.A2(n_1138),
.B(n_1166),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1107),
.A2(n_1172),
.B(n_1101),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1116),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1172),
.A2(n_1140),
.B(n_1122),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1125),
.A2(n_1109),
.A3(n_1187),
.B(n_1088),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1091),
.A2(n_1147),
.B(n_1187),
.C(n_1134),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1187),
.A2(n_1152),
.B(n_1076),
.C(n_1155),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1152),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1183),
.A2(n_1108),
.B(n_1135),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_L g1252 ( 
.A(n_1149),
.B(n_1136),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1067),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1067),
.B(n_730),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1077),
.B(n_1089),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1151),
.A2(n_650),
.B(n_1162),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1077),
.B(n_1089),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1097),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1086),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1167),
.B(n_1115),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1130),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1082),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1145),
.A2(n_1159),
.B(n_1154),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1100),
.B(n_1035),
.Y(n_1265)
);

AOI322xp5_ASAP7_75t_L g1266 ( 
.A1(n_1176),
.A2(n_497),
.A3(n_763),
.B1(n_753),
.B2(n_354),
.C1(n_386),
.C2(n_777),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1090),
.B(n_1094),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1156),
.A2(n_1171),
.B1(n_1178),
.B2(n_1177),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1151),
.A2(n_1162),
.B(n_763),
.C(n_1141),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1176),
.A2(n_1175),
.B1(n_1089),
.B2(n_1181),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1131),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1087),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1100),
.B(n_1035),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1090),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1130),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1151),
.A2(n_650),
.B(n_1162),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1175),
.B(n_1089),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1100),
.B(n_1035),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1151),
.A2(n_1162),
.B(n_763),
.C(n_1141),
.Y(n_1284)
);

AO22x2_ASAP7_75t_L g1285 ( 
.A1(n_1089),
.A2(n_1174),
.B1(n_1093),
.B2(n_1158),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1097),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1136),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1167),
.B(n_1115),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1131),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1130),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1131),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1153),
.A2(n_1157),
.B(n_1154),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1130),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1097),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1076),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1145),
.A2(n_1159),
.B(n_1154),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1181),
.A2(n_1174),
.A3(n_1089),
.B(n_1048),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1077),
.B(n_1089),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1191),
.B(n_1276),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1197),
.B(n_1268),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1227),
.A2(n_1216),
.B(n_1205),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1285),
.B(n_1219),
.Y(n_1303)
);

OAI31xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1215),
.A2(n_1203),
.A3(n_1282),
.B(n_1221),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1226),
.B(n_1193),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1252),
.B(n_1251),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1256),
.A2(n_1280),
.B(n_1284),
.C(n_1269),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1193),
.B(n_1260),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1260),
.B(n_1289),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1289),
.B(n_1267),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1285),
.B(n_1232),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1190),
.B(n_1258),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1285),
.B(n_1232),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1229),
.A2(n_1205),
.B(n_1284),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1298),
.B(n_1202),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1194),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1262),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1298),
.B(n_1202),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1298),
.B(n_1198),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1204),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1270),
.A2(n_1229),
.B1(n_1215),
.B2(n_1201),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1286),
.B(n_1295),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1199),
.B(n_1259),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1298),
.B(n_1206),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1199),
.B(n_1259),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1282),
.A2(n_1225),
.B(n_1230),
.C(n_1248),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1248),
.A2(n_1249),
.B(n_1283),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1206),
.B(n_1247),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1206),
.B(n_1247),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1206),
.B(n_1247),
.Y(n_1330)
);

BUFx2_ASAP7_75t_R g1331 ( 
.A(n_1237),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1270),
.B(n_1233),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1210),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1239),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1249),
.A2(n_1265),
.B(n_1273),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1210),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1209),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1210),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1195),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1233),
.B(n_1271),
.Y(n_1341)
);

NAND2x1_ASAP7_75t_L g1342 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1299),
.A2(n_1242),
.B1(n_1254),
.B2(n_1241),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1218),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1220),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1290),
.B(n_1292),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1224),
.B(n_1288),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1262),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1208),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1243),
.A2(n_1211),
.B(n_1222),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1231),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1254),
.A2(n_1217),
.B1(n_1238),
.B2(n_1244),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1228),
.Y(n_1353)
);

O2A1O1Ixp5_ASAP7_75t_L g1354 ( 
.A1(n_1243),
.A2(n_1250),
.B(n_1253),
.C(n_1238),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1213),
.A2(n_1240),
.B1(n_1253),
.B2(n_1272),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1200),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_L g1357 ( 
.A1(n_1250),
.A2(n_1223),
.B(n_1272),
.C(n_1235),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1246),
.B(n_1297),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1266),
.B(n_1245),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1264),
.B(n_1297),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1264),
.B(n_1297),
.Y(n_1361)
);

BUFx4f_ASAP7_75t_SL g1362 ( 
.A(n_1236),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1192),
.A2(n_1281),
.B(n_1275),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1263),
.A2(n_1287),
.B(n_1274),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1278),
.A2(n_1279),
.B(n_1293),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1296),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1234),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1296),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1212),
.A2(n_1196),
.B(n_1277),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1214),
.A2(n_1261),
.B1(n_1277),
.B2(n_1291),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1291),
.A2(n_1227),
.B(n_1216),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1294),
.B(n_1197),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1294),
.B(n_1197),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1262),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1191),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1207),
.Y(n_1376)
);

AND2x2_ASAP7_75t_SL g1377 ( 
.A(n_1270),
.B(n_1175),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1191),
.B(n_1276),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1360),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1328),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1337),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1303),
.B(n_1324),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1360),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1367),
.A2(n_1324),
.B(n_1302),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1314),
.A2(n_1307),
.B(n_1304),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_1375),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1328),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1361),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1358),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1329),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1321),
.A2(n_1301),
.B(n_1377),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1371),
.A2(n_1350),
.B(n_1303),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1377),
.A2(n_1326),
.B(n_1357),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1358),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1315),
.B(n_1318),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1327),
.B(n_1335),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1315),
.B(n_1318),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1344),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1330),
.A2(n_1332),
.B(n_1313),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1345),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1319),
.B(n_1330),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1316),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1311),
.A2(n_1313),
.B(n_1370),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1319),
.B(n_1311),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1333),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1320),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1308),
.B(n_1309),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_1310),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1343),
.A2(n_1355),
.B(n_1338),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1369),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1351),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1363),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1353),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1363),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1364),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1300),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1364),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1312),
.A2(n_1352),
.B(n_1339),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1306),
.B(n_1347),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1322),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1365),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1365),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1379),
.B(n_1383),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1383),
.B(n_1365),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1411),
.Y(n_1429)
);

OAI211xp5_ASAP7_75t_L g1430 ( 
.A1(n_1385),
.A2(n_1342),
.B(n_1376),
.C(n_1340),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1388),
.B(n_1378),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1388),
.B(n_1423),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1389),
.B(n_1341),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1416),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1419),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1389),
.B(n_1306),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1423),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1389),
.B(n_1306),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1381),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1394),
.B(n_1346),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.B(n_1347),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1368),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1397),
.B(n_1366),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1397),
.B(n_1349),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1431),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_R g1449 ( 
.A(n_1445),
.B(n_1317),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1437),
.A2(n_1385),
.B1(n_1391),
.B2(n_1393),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1431),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1430),
.A2(n_1391),
.B1(n_1393),
.B2(n_1414),
.C(n_1408),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1445),
.B(n_1414),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1429),
.A2(n_1382),
.B1(n_1405),
.B2(n_1404),
.C(n_1392),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1406),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1429),
.A2(n_1382),
.B1(n_1405),
.B2(n_1404),
.C(n_1392),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1443),
.B(n_1420),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1435),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1442),
.A2(n_1404),
.B1(n_1400),
.B2(n_1382),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1430),
.A2(n_1396),
.B(n_1410),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1443),
.B(n_1418),
.C(n_1425),
.Y(n_1461)
);

AOI222xp33_ASAP7_75t_L g1462 ( 
.A1(n_1447),
.A2(n_1359),
.B1(n_1405),
.B2(n_1390),
.C1(n_1387),
.C2(n_1380),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1443),
.Y(n_1463)
);

OAI33xp33_ASAP7_75t_L g1464 ( 
.A1(n_1442),
.A2(n_1408),
.A3(n_1424),
.B1(n_1409),
.B2(n_1413),
.B3(n_1380),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1428),
.A2(n_1404),
.B1(n_1392),
.B2(n_1380),
.C(n_1390),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1436),
.A2(n_1426),
.B(n_1421),
.Y(n_1466)
);

AOI33xp33_ASAP7_75t_L g1467 ( 
.A1(n_1439),
.A2(n_1399),
.A3(n_1401),
.B1(n_1407),
.B2(n_1403),
.B3(n_1413),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1442),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1437),
.A2(n_1404),
.B1(n_1400),
.B2(n_1392),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1438),
.B(n_1396),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1437),
.A2(n_1400),
.B1(n_1392),
.B2(n_1387),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1436),
.A2(n_1426),
.B(n_1421),
.Y(n_1472)
);

OAI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1440),
.A2(n_1396),
.B1(n_1424),
.B2(n_1387),
.C(n_1390),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1420),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1435),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1434),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1439),
.B(n_1394),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1440),
.A2(n_1386),
.B(n_1425),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.B(n_1386),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1446),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1447),
.A2(n_1400),
.B1(n_1422),
.B2(n_1384),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1446),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1466),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

INVx4_ASAP7_75t_SL g1488 ( 
.A(n_1470),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1455),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1466),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1465),
.A2(n_1418),
.B(n_1425),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1466),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1448),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1441),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1460),
.A2(n_1396),
.B(n_1384),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1449),
.B(n_1434),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_SL g1498 ( 
.A(n_1454),
.B(n_1317),
.C(n_1374),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1451),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1452),
.B(n_1362),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1470),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1456),
.B(n_1433),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1458),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1475),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1472),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1472),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1455),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1469),
.A2(n_1418),
.B(n_1415),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1482),
.A2(n_1415),
.B(n_1426),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1472),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1450),
.B(n_1417),
.C(n_1412),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1427),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1516)
);

BUFx8_ASAP7_75t_L g1517 ( 
.A(n_1468),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1463),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1497),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1494),
.B(n_1468),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1502),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1514),
.B(n_1461),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1494),
.B(n_1457),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1331),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1502),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1504),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1457),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1498),
.B(n_1464),
.C(n_1461),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1512),
.B(n_1513),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1519),
.B(n_1476),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1490),
.Y(n_1535)
);

NAND4xp75_ASAP7_75t_L g1536 ( 
.A(n_1491),
.B(n_1354),
.C(n_1336),
.D(n_1402),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1504),
.Y(n_1537)
);

NOR2x1p5_ASAP7_75t_L g1538 ( 
.A(n_1498),
.B(n_1348),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1487),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1518),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1493),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1493),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1514),
.A2(n_1374),
.B1(n_1348),
.B2(n_1356),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1491),
.A2(n_1462),
.B(n_1471),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1488),
.B(n_1484),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1488),
.B(n_1438),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1519),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1490),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1491),
.B(n_1462),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1480),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1503),
.A2(n_1459),
.B1(n_1478),
.B2(n_1495),
.C(n_1516),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1517),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1490),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1515),
.B(n_1485),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1489),
.B(n_1485),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1496),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1496),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1491),
.B(n_1478),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1489),
.B(n_1508),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1540),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1491),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1560),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1560),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1539),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1568)
);

NOR2xp67_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1508),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_SL g1571 ( 
.A(n_1532),
.B(n_1495),
.C(n_1473),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1541),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1499),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1554),
.B(n_1488),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1523),
.B(n_1508),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1541),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1517),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.B(n_1544),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1531),
.B(n_1505),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1520),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1488),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1542),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1542),
.Y(n_1584)
);

NAND2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1545),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1522),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1520),
.B(n_1517),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1545),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1528),
.B(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1543),
.Y(n_1591)
);

AOI31xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1553),
.A2(n_1474),
.A3(n_1481),
.B(n_1432),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1543),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.B(n_1479),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_SL g1596 ( 
.A(n_1536),
.B(n_1501),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1551),
.A2(n_1509),
.B(n_1510),
.C(n_1507),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1572),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1580),
.B(n_1546),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1580),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1591),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1591),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1546),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1578),
.B(n_1524),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1588),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1570),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1577),
.B(n_1356),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1574),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1576),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1564),
.B(n_1524),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1590),
.B(n_1552),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1583),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1568),
.B(n_1531),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1589),
.A2(n_1557),
.B(n_1561),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1579),
.B(n_1529),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1574),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1590),
.B(n_1556),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1564),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_L g1623 ( 
.A1(n_1599),
.A2(n_1604),
.B1(n_1571),
.B2(n_1563),
.C1(n_1565),
.C2(n_1600),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1610),
.B(n_1596),
.Y(n_1624)
);

OAI211xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1619),
.A2(n_1586),
.B(n_1565),
.C(n_1582),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1618),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1568),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1613),
.A2(n_1597),
.B1(n_1595),
.B2(n_1585),
.C(n_1592),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1621),
.A2(n_1593),
.B(n_1585),
.Y(n_1629)
);

AOI211xp5_ASAP7_75t_L g1630 ( 
.A1(n_1617),
.A2(n_1574),
.B(n_1569),
.C(n_1581),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1618),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1611),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1610),
.B(n_1581),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1611),
.B(n_1594),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1621),
.A2(n_1585),
.B(n_1587),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1605),
.A2(n_1581),
.B1(n_1573),
.B2(n_1501),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1606),
.B(n_1529),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.B(n_1620),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1608),
.B(n_1530),
.Y(n_1639)
);

OAI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1614),
.A2(n_1573),
.B(n_1567),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1598),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1638),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1632),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1627),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1634),
.B(n_1640),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1633),
.B(n_1620),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1630),
.B(n_1609),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1625),
.B(n_1607),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1626),
.B(n_1594),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1623),
.B(n_1607),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1624),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1631),
.B(n_1612),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1637),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1650),
.A2(n_1628),
.B(n_1629),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1648),
.B(n_1629),
.C(n_1639),
.D(n_1637),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1650),
.A2(n_1509),
.B1(n_1510),
.B2(n_1639),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1648),
.A2(n_1636),
.B(n_1609),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1653),
.A2(n_1635),
.B(n_1641),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1642),
.B(n_1615),
.Y(n_1659)
);

NOR4xp25_ASAP7_75t_L g1660 ( 
.A(n_1651),
.B(n_1642),
.C(n_1644),
.D(n_1652),
.Y(n_1660)
);

AOI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1643),
.A2(n_1602),
.B(n_1601),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_1645),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1663)
);

NOR4xp25_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1646),
.C(n_1647),
.D(n_1603),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1656),
.A2(n_1587),
.B1(n_1555),
.B2(n_1550),
.C(n_1535),
.Y(n_1665)
);

AO21x1_ASAP7_75t_L g1666 ( 
.A1(n_1658),
.A2(n_1537),
.B(n_1530),
.Y(n_1666)
);

O2A1O1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1660),
.A2(n_1555),
.B(n_1550),
.C(n_1522),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1662),
.Y(n_1668)
);

AOI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1655),
.A2(n_1575),
.B(n_1567),
.C(n_1579),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1664),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_SL g1672 ( 
.A(n_1666),
.B(n_1659),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1669),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1667),
.B(n_1663),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1665),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1672),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1671),
.B(n_1657),
.C(n_1661),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1674),
.A2(n_1537),
.B(n_1575),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1670),
.A2(n_1536),
.B(n_1535),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

NAND2x1p5_ASAP7_75t_L g1681 ( 
.A(n_1680),
.B(n_1675),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_SL g1682 ( 
.A(n_1677),
.B(n_1535),
.C(n_1522),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1676),
.A2(n_1538),
.B1(n_1550),
.B2(n_1555),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1681),
.B(n_1678),
.C(n_1679),
.Y(n_1684)
);

OAI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1682),
.B(n_1683),
.C(n_1561),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1685),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1685),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1686),
.B(n_1492),
.C(n_1486),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1687),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1689),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1688),
.B(n_1558),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1690),
.Y(n_1692)
);

AO221x2_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1691),
.B1(n_1559),
.B2(n_1558),
.C(n_1538),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1693),
.B(n_1547),
.Y(n_1694)
);

AOI322xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1547),
.A3(n_1548),
.B1(n_1486),
.B2(n_1511),
.C1(n_1506),
.C2(n_1507),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1695),
.A2(n_1547),
.B1(n_1548),
.B2(n_1507),
.Y(n_1696)
);

AOI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1559),
.B(n_1557),
.C(n_1486),
.Y(n_1697)
);


endmodule