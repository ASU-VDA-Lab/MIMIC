module fake_jpeg_108_n_120 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_40),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_16),
.B1(n_22),
.B2(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_4),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_24),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_20),
.B1(n_33),
.B2(n_35),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_26),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_26),
.Y(n_53)
);

AO21x1_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_56),
.B(n_59),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_29),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_27),
.B(n_16),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_38),
.B1(n_27),
.B2(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_7),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_10),
.C(n_11),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_47),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_8),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_10),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_57),
.Y(n_73)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_45),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_53),
.CI(n_60),
.CON(n_77),
.SN(n_77)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_56),
.C(n_54),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_74),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_69),
.B1(n_62),
.B2(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_95),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_72),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_74),
.A3(n_65),
.B1(n_86),
.B2(n_77),
.C1(n_69),
.C2(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_79),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_77),
.C(n_76),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_78),
.C(n_63),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.C(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_58),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_92),
.B1(n_50),
.B2(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_68),
.C(n_27),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_67),
.C(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_97),
.B1(n_107),
.B2(n_11),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_112),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_97),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_111),
.B(n_13),
.C(n_43),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_43),
.Y(n_120)
);


endmodule