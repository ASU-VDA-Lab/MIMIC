module real_jpeg_23528_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_79),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_1),
.A2(n_64),
.B1(n_66),
.B2(n_79),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_1),
.A2(n_53),
.B1(n_59),
.B2(n_79),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_63),
.B1(n_85),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_2),
.A2(n_53),
.B1(n_59),
.B2(n_63),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_84),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_84),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_6),
.A2(n_53),
.B1(n_59),
.B2(n_84),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_30),
.B1(n_141),
.B2(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_168),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_7),
.A2(n_64),
.B1(n_66),
.B2(n_168),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_7),
.A2(n_53),
.B1(n_59),
.B2(n_168),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_41),
.B1(n_64),
.B2(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_41),
.B1(n_53),
.B2(n_59),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_41),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_36),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_21),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_64),
.C(n_91),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_221),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_11),
.B(n_132),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_11),
.A2(n_64),
.B1(n_66),
.B2(n_221),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_11),
.B(n_53),
.C(n_69),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_11),
.A2(n_52),
.B(n_282),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_22),
.B1(n_27),
.B2(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_13),
.A2(n_64),
.B1(n_66),
.B2(n_117),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_13),
.A2(n_53),
.B1(n_59),
.B2(n_117),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_22),
.B1(n_27),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_14),
.A2(n_64),
.B1(n_66),
.B2(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_30),
.B1(n_95),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_14),
.A2(n_53),
.B1(n_59),
.B2(n_95),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_34),
.B1(n_53),
.B2(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_34),
.B1(n_64),
.B2(n_66),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_34),
.Y(n_156)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_16),
.A2(n_190),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_42),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_28),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_21),
.A2(n_28),
.B1(n_116),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_21),
.A2(n_28),
.B1(n_40),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_27),
.B1(n_91),
.B2(n_92),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_22),
.B(n_26),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_22),
.B(n_245),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_25),
.A2(n_27),
.A3(n_31),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_28),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_28),
.A2(n_120),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_30),
.Y(n_141)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_32),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_32),
.B(n_82),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_32),
.A2(n_78),
.B1(n_118),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_32),
.A2(n_118),
.B1(n_140),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_32),
.A2(n_80),
.B(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_39),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_39),
.B(n_354),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_353),
.B(n_355),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_341),
.B(n_352),
.Y(n_45)
);

OAI31xp33_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_143),
.A3(n_158),
.B(n_338),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_121),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_48),
.B(n_121),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_86),
.C(n_102),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_49),
.A2(n_86),
.B1(n_87),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_49),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_74),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_51),
.B(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_51),
.A2(n_60),
.B1(n_61),
.B2(n_75),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_58),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_55),
.B1(n_58),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_52),
.A2(n_55),
.B1(n_107),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_52),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_52),
.A2(n_192),
.B1(n_194),
.B2(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_52),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_52),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_54),
.Y(n_250)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_57),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_57),
.B(n_221),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_59),
.B(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_67),
.B1(n_73),
.B2(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_66),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_64),
.B(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_73),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_67),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_67),
.A2(n_73),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_71),
.A2(n_98),
.B1(n_111),
.B2(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_71),
.A2(n_178),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_71),
.A2(n_217),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_71),
.B(n_221),
.Y(n_301)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_73),
.B(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_85),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_89),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_89),
.A2(n_90),
.B1(n_134),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_89),
.A2(n_185),
.B(n_187),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_89),
.A2(n_187),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_90),
.A2(n_113),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_90),
.A2(n_171),
.B(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_96),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_98),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_98),
.A2(n_270),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_102),
.A2(n_103),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.C(n_114),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_104),
.A2(n_105),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_112),
.B(n_114),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_124),
.C(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_139),
.B2(n_142),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_136),
.C(n_139),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_131),
.A2(n_132),
.B1(n_186),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_131),
.A2(n_132),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_132),
.B(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_136),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_136),
.B(n_150),
.C(n_155),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_142),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_139),
.B(n_146),
.C(n_149),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_144),
.A2(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_145),
.B(n_157),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_151),
.Y(n_348)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_156),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_331),
.B(n_337),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_206),
.B(n_330),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_199),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_161),
.B(n_199),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_179),
.C(n_181),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_162),
.A2(n_163),
.B1(n_179),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_173),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_169),
.C(n_173),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_179),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_181),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_188),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_184),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_196),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_194),
.A2(n_295),
.B(n_303),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_336)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_237),
.B(n_324),
.C(n_329),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_231),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_231),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_223),
.C(n_224),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_209),
.A2(n_210),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_215),
.C(n_219),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_223),
.B(n_224),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_229),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_318),
.B(n_323),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_271),
.B(n_317),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_260),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_260),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.C(n_257),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_246),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B(n_251),
.Y(n_246)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_267),
.C(n_268),
.Y(n_322)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_311),
.B(n_316),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_291),
.B(n_310),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_285),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_285),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_315)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_289),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_299),
.B(n_309),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_297),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_304),
.B(n_308),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_336),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_336),
.Y(n_337)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_343),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_351),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_345),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_347),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_349),
.C(n_351),
.Y(n_354)
);


endmodule