module fake_jpeg_30122_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_39),
.C(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_2),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_12),
.A2(n_3),
.B(n_4),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_18),
.B1(n_16),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_43),
.B1(n_38),
.B2(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_27),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_37),
.B1(n_20),
.B2(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_67),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_45),
.C(n_54),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_46),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_48),
.B1(n_53),
.B2(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_49),
.B1(n_45),
.B2(n_40),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_38),
.B1(n_46),
.B2(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_73),
.B(n_38),
.Y(n_79)
);

BUFx24_ASAP7_75t_SL g77 ( 
.A(n_71),
.Y(n_77)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_44),
.B(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_80),
.C(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_40),
.B1(n_51),
.B2(n_47),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_70),
.B1(n_59),
.B2(n_71),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_38),
.B(n_41),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_46),
.B1(n_68),
.B2(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_91),
.B1(n_82),
.B2(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_70),
.C(n_63),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_95),
.C(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_61),
.B1(n_69),
.B2(n_62),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_59),
.B(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_70),
.C(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_82),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_103),
.C(n_95),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_77),
.B(n_58),
.C(n_73),
.D(n_60),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_84),
.B(n_32),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_31),
.B(n_29),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_107),
.C(n_99),
.Y(n_111)
);

AO221x1_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_6),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_90),
.C(n_89),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_32),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_104),
.C(n_102),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_108),
.B(n_97),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_100),
.B(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_97),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_118),
.B(n_116),
.C(n_9),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_8),
.B(n_9),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_56),
.Y(n_121)
);


endmodule