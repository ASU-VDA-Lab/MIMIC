module fake_jpeg_11466_n_41 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_18),
.B(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.C(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_25),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_25),
.B(n_16),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_36),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_41)
);


endmodule