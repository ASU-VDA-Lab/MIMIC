module fake_netlist_1_5195_n_38 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_4), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_6), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_15), .B(n_1), .Y(n_22) );
INVxp67_ASAP7_75t_SL g23 ( .A(n_17), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
BUFx12f_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_14), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_25), .Y(n_28) );
AOI32xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_18), .A3(n_20), .B1(n_25), .B2(n_19), .Y(n_29) );
NAND3xp33_ASAP7_75t_L g30 ( .A(n_27), .B(n_19), .C(n_16), .Y(n_30) );
XOR2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_20), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_18), .B1(n_19), .B2(n_16), .Y(n_32) );
NOR2x1_ASAP7_75t_SL g33 ( .A(n_31), .B(n_16), .Y(n_33) );
AND4x1_ASAP7_75t_L g34 ( .A(n_32), .B(n_19), .C(n_7), .D(n_8), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
NOR3xp33_ASAP7_75t_L g36 ( .A(n_33), .B(n_16), .C(n_9), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
AOI322xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_36), .A3(n_34), .B1(n_11), .B2(n_12), .C1(n_13), .C2(n_10), .Y(n_38) );
endmodule