module fake_jpeg_19312_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_65),
.B1(n_51),
.B2(n_59),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_63),
.B1(n_35),
.B2(n_18),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_44),
.B1(n_38),
.B2(n_35),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_71),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_73),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_39),
.B1(n_44),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_87),
.B1(n_92),
.B2(n_104),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_86),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_57),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_76),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_44),
.B1(n_35),
.B2(n_38),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_95),
.B1(n_96),
.B2(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_82),
.B1(n_93),
.B2(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_37),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_44),
.B1(n_43),
.B2(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_89),
.Y(n_138)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_33),
.B1(n_18),
.B2(n_16),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_30),
.B1(n_26),
.B2(n_16),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_27),
.B1(n_32),
.B2(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_108),
.Y(n_137)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_42),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_42),
.Y(n_109)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_41),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_27),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.C(n_127),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_23),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_131),
.B1(n_106),
.B2(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_11),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_41),
.B1(n_40),
.B2(n_36),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_91),
.B1(n_67),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_126),
.B1(n_135),
.B2(n_137),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_24),
.C(n_31),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.C(n_36),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_31),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_134),
.B1(n_119),
.B2(n_118),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_67),
.A3(n_106),
.B1(n_90),
.B2(n_99),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_101),
.B1(n_89),
.B2(n_78),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_147),
.B1(n_159),
.B2(n_113),
.Y(n_179)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_152),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_70),
.B1(n_94),
.B2(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_41),
.B(n_40),
.C(n_36),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_113),
.B1(n_110),
.B2(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_70),
.B1(n_85),
.B2(n_104),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_158),
.B1(n_165),
.B2(n_131),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_98),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_107),
.B1(n_80),
.B2(n_40),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_118),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_105),
.C(n_36),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_168),
.C(n_0),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_112),
.B(n_114),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_36),
.B1(n_105),
.B2(n_32),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_24),
.B(n_22),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_4),
.B(n_5),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_109),
.C(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_32),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_0),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_173),
.B(n_190),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_176),
.B1(n_191),
.B2(n_193),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_113),
.B1(n_116),
.B2(n_110),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_187),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_144),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_22),
.B(n_1),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_183),
.B(n_184),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_22),
.B1(n_14),
.B2(n_13),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_142),
.B1(n_149),
.B2(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_150),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_203),
.B1(n_187),
.B2(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_182),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_170),
.B1(n_156),
.B2(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_140),
.A2(n_157),
.B1(n_161),
.B2(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_206),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_209),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_207),
.B(n_210),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_150),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_219),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_188),
.C(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_221),
.C(n_223),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_227),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_151),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_220),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_153),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_146),
.C(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_171),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_225),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_231),
.B1(n_199),
.B2(n_185),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_12),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_197),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_5),
.B(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_173),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_241),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_203),
.B1(n_172),
.B2(n_179),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_238),
.B1(n_252),
.B2(n_254),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_189),
.B1(n_196),
.B2(n_174),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_231),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_177),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_177),
.B1(n_201),
.B2(n_200),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_190),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_208),
.B1(n_211),
.B2(n_215),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_261),
.A2(n_270),
.B1(n_275),
.B2(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_209),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_239),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_223),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_240),
.Y(n_276)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_212),
.C(n_205),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_271),
.C(n_272),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_213),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_218),
.B1(n_226),
.B2(n_177),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_228),
.C(n_198),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_255),
.C(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_183),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_254),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_229),
.C(n_185),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_233),
.C(n_246),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_5),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_280),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_258),
.B(n_237),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_249),
.C(n_234),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_257),
.B1(n_259),
.B2(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_229),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_249),
.C(n_234),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_263),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_296),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_269),
.B1(n_244),
.B2(n_265),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_280),
.B1(n_283),
.B2(n_277),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_270),
.B(n_7),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_7),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_309),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_287),
.C(n_285),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_285),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_277),
.B(n_276),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_299),
.B(n_292),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_307),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_298),
.B(n_296),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_298),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_318),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_314),
.B(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_310),
.C(n_320),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_324),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_306),
.Y(n_327)
);

AOI311xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_304),
.A3(n_9),
.B(n_10),
.C(n_8),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_8),
.B(n_10),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_8),
.B(n_10),
.Y(n_330)
);


endmodule