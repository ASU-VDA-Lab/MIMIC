module fake_jpeg_29141_n_513 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_513);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_513;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_60),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_28),
.B(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_73),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_70),
.Y(n_123)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_29),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_43),
.Y(n_105)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_44),
.B(n_7),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_119),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_129),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_113),
.B(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_83),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_71),
.B(n_50),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_94),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_148),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_56),
.B(n_0),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_95),
.C(n_49),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

CKINVDCx12_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_162),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_182),
.B1(n_184),
.B2(n_196),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_168),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_78),
.B1(n_59),
.B2(n_58),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_134),
.B1(n_155),
.B2(n_149),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_117),
.A2(n_52),
.B1(n_53),
.B2(n_99),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_173),
.A2(n_180),
.B1(n_190),
.B2(n_197),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_36),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_211),
.Y(n_232)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_36),
.Y(n_178)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_74),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_215),
.C(n_127),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_97),
.B1(n_100),
.B2(n_93),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_181),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_26),
.B1(n_42),
.B2(n_32),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_105),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_189),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_108),
.A2(n_133),
.B1(n_103),
.B2(n_132),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_103),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_118),
.A2(n_92),
.B1(n_88),
.B2(n_91),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

BUFx24_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_32),
.B1(n_101),
.B2(n_49),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_49),
.B1(n_33),
.B2(n_25),
.Y(n_197)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

AO22x2_ASAP7_75t_L g201 ( 
.A1(n_124),
.A2(n_55),
.B1(n_94),
.B2(n_96),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_201),
.A2(n_153),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_155),
.B1(n_159),
.B2(n_130),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_140),
.B1(n_123),
.B2(n_96),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_141),
.B(n_41),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_107),
.B(n_25),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_115),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_123),
.Y(n_224)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_49),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_11),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_218),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_104),
.B(n_33),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_221),
.A2(n_222),
.B1(n_242),
.B2(n_188),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_149),
.B1(n_126),
.B2(n_128),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_240),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_167),
.A2(n_160),
.B(n_131),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_197),
.B(n_180),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_33),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_137),
.B1(n_122),
.B2(n_140),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_258),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_246),
.A2(n_198),
.B1(n_169),
.B2(n_202),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_171),
.A2(n_135),
.B(n_148),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_260),
.B(n_264),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_201),
.A2(n_0),
.B(n_1),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_1),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_187),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_201),
.A2(n_165),
.B(n_203),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_266),
.B(n_268),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_279),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_273),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_181),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_168),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_209),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_277),
.B(n_290),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_191),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_173),
.B(n_216),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_280),
.B(n_283),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_166),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_199),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_293),
.Y(n_325)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_193),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_285),
.B(n_286),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_300),
.B1(n_251),
.B2(n_261),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_193),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_292),
.B(n_294),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_207),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_234),
.B(n_15),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_253),
.B1(n_219),
.B2(n_230),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_198),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_304),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_169),
.C(n_185),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_249),
.C(n_243),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_336)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_225),
.C(n_223),
.D(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_254),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_220),
.B(n_12),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_307),
.A2(n_315),
.B1(n_330),
.B2(n_337),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_259),
.B(n_251),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_321),
.B(n_295),
.Y(n_358)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_319),
.C(n_342),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_293),
.A2(n_253),
.B1(n_262),
.B2(n_248),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_286),
.A2(n_261),
.B1(n_219),
.B2(n_259),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_227),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_320),
.A2(n_338),
.B1(n_304),
.B2(n_268),
.Y(n_343)
);

OAI22x1_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_223),
.B1(n_195),
.B2(n_210),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_328),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_288),
.A2(n_174),
.B1(n_164),
.B2(n_236),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_281),
.A2(n_236),
.B1(n_230),
.B2(n_223),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_279),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_296),
.A2(n_11),
.B1(n_13),
.B2(n_7),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_275),
.A2(n_8),
.B1(n_12),
.B2(n_15),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_15),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_362),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_312),
.B(n_280),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_344),
.B(n_346),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_294),
.Y(n_346)
);

INVx13_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_348),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_306),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_353),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_323),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_369),
.C(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_266),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_276),
.Y(n_354)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_275),
.B1(n_281),
.B2(n_285),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_356),
.A2(n_364),
.B1(n_320),
.B2(n_315),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_370),
.B(n_366),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_273),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_361),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_270),
.Y(n_360)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_274),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_332),
.A2(n_296),
.B1(n_300),
.B2(n_279),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_334),
.B(n_274),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_316),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_279),
.B1(n_284),
.B2(n_283),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_366),
.A2(n_367),
.B(n_311),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_297),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_306),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_371),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_298),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_324),
.A2(n_272),
.B(n_269),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_292),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_265),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_337),
.Y(n_388)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

OR2x2_ASAP7_75t_SL g375 ( 
.A(n_340),
.B(n_265),
.Y(n_375)
);

XOR2x2_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_297),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_380),
.C(n_396),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_342),
.C(n_316),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_364),
.Y(n_408)
);

XOR2x2_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_327),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_384),
.B(n_405),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_404),
.Y(n_407)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_389),
.B(n_391),
.Y(n_423)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_325),
.B(n_331),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_335),
.C(n_333),
.Y(n_396)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_399),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_401),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_362),
.B1(n_343),
.B2(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_403),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_366),
.A2(n_326),
.B(n_322),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_408),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_412),
.A2(n_415),
.B1(n_416),
.B2(n_421),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_356),
.B1(n_355),
.B2(n_345),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_376),
.A2(n_355),
.B1(n_358),
.B2(n_373),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_349),
.C(n_374),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_424),
.C(n_428),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_402),
.A2(n_367),
.B1(n_373),
.B2(n_357),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_339),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_386),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_357),
.C(n_339),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_394),
.B(n_348),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_425),
.B(n_429),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_291),
.Y(n_426)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_326),
.C(n_347),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_395),
.B(n_313),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_287),
.Y(n_430)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_379),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_431),
.B(n_435),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_427),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_433),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_393),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_439),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_410),
.B(n_389),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_405),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_443),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_410),
.B(n_412),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_450),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_382),
.C(n_404),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_408),
.C(n_429),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_383),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_449),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_391),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_451),
.B(n_460),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_452),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_423),
.C(n_415),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_455),
.C(n_456),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_447),
.C(n_449),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_421),
.C(n_407),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_398),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_433),
.B(n_385),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_462),
.B(n_465),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_388),
.Y(n_465)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_445),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_469),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_453),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_463),
.A2(n_413),
.B1(n_387),
.B2(n_381),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_472),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_414),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_451),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_480),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_459),
.B(n_387),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_477),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_457),
.A2(n_416),
.B1(n_417),
.B2(n_381),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_475),
.A2(n_471),
.B1(n_464),
.B2(n_397),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_443),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_478),
.B(n_438),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_438),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_468),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_392),
.Y(n_498)
);

INVx6_ASAP7_75t_L g482 ( 
.A(n_476),
.Y(n_482)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_482),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_488),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_397),
.B1(n_403),
.B2(n_401),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_484),
.B(n_491),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_480),
.A2(n_425),
.B(n_377),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_479),
.A2(n_420),
.B(n_392),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_467),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_496),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_479),
.C(n_469),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_481),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_482),
.C(n_485),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_499),
.B(n_501),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_489),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_502),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_377),
.Y(n_502)
);

AOI21xp33_ASAP7_75t_L g505 ( 
.A1(n_503),
.A2(n_492),
.B(n_490),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g508 ( 
.A1(n_505),
.A2(n_492),
.A3(n_399),
.B1(n_265),
.B2(n_297),
.C1(n_301),
.C2(n_5),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_500),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_508),
.C(n_504),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_4),
.C(n_5),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_4),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_511),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_4),
.Y(n_513)
);


endmodule