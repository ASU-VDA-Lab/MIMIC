module fake_jpeg_26300_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_58),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_22),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_51),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_32),
.B1(n_42),
.B2(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_43),
.B1(n_26),
.B2(n_24),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_34),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_25),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_30),
.C(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_21),
.B1(n_23),
.B2(n_40),
.Y(n_75)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_30),
.B1(n_27),
.B2(n_19),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_31),
.B1(n_20),
.B2(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_67),
.Y(n_120)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_75),
.B1(n_88),
.B2(n_96),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_84),
.B1(n_93),
.B2(n_59),
.Y(n_125)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_98),
.Y(n_106)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_R g115 ( 
.A(n_83),
.B(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_41),
.B1(n_37),
.B2(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_89),
.Y(n_123)
);

HB1xp67_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_41),
.B1(n_30),
.B2(n_27),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_31),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_57),
.B1(n_55),
.B2(n_64),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_93),
.B1(n_109),
.B2(n_118),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_74),
.Y(n_127)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_104),
.B1(n_111),
.B2(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_0),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_129),
.B(n_17),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_74),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_132),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_98),
.B(n_82),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_140),
.B1(n_144),
.B2(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_77),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_87),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_107),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_146),
.B1(n_39),
.B2(n_4),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_99),
.B1(n_85),
.B2(n_91),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_58),
.C(n_71),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_149),
.C(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_72),
.B1(n_78),
.B2(n_49),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_52),
.B1(n_49),
.B2(n_45),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_52),
.C(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_52),
.B1(n_45),
.B2(n_27),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.C(n_101),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_158),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_152),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_102),
.B(n_105),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_159),
.B(n_169),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_122),
.B(n_108),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_165),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_17),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_173),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_110),
.B1(n_17),
.B2(n_121),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_142),
.B1(n_148),
.B2(n_145),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_16),
.A3(n_15),
.B1(n_39),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_126),
.B(n_15),
.C(n_7),
.D(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_133),
.B1(n_151),
.B2(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_149),
.C(n_143),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_174),
.C(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_156),
.B1(n_173),
.B2(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_187),
.Y(n_200)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_130),
.B1(n_128),
.B2(n_141),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_128),
.B(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_134),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_192),
.A3(n_194),
.B1(n_170),
.B2(n_157),
.C(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_147),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_199),
.B1(n_209),
.B2(n_188),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_162),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_202),
.C(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_169),
.B(n_159),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_158),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_190),
.C(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_179),
.C(n_160),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_182),
.B1(n_187),
.B2(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_186),
.B1(n_179),
.B2(n_185),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_217),
.B1(n_205),
.B2(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_153),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_190),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_202),
.C(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_199),
.B(n_160),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_150),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_224),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_206),
.B(n_198),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_10),
.C(n_11),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_215),
.B(n_5),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_192),
.B(n_5),
.C(n_9),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_223),
.B1(n_215),
.B2(n_9),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_228),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_231),
.B(n_225),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_12),
.B(n_13),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_234),
.C(n_239),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_238),
.C(n_230),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_14),
.B(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_252),
.A2(n_251),
.B(n_14),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_14),
.Y(n_254)
);


endmodule