module fake_jpeg_19862_n_85 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx24_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_10),
.B(n_14),
.C(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2x1_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_19),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_18),
.B1(n_17),
.B2(n_11),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_19),
.C(n_22),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_24),
.B1(n_11),
.B2(n_8),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_13),
.B1(n_9),
.B2(n_14),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_9),
.B1(n_19),
.B2(n_15),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_36),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_30),
.B(n_32),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_31),
.B1(n_34),
.B2(n_3),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_47),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_45),
.C(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_58),
.B1(n_44),
.B2(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_45),
.C(n_31),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_34),
.C(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AOI21x1_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_59),
.B(n_2),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_1),
.B(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_66),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_70),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_75),
.C(n_74),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_68),
.C(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_7),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_4),
.B(n_5),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_4),
.C(n_5),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_5),
.Y(n_85)
);


endmodule