module real_jpeg_23694_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_1),
.A2(n_70),
.B1(n_73),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_1),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_60),
.B1(n_65),
.B2(n_109),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_1),
.A2(n_27),
.B1(n_33),
.B2(n_109),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_27),
.B1(n_33),
.B2(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_3),
.A2(n_47),
.B1(n_60),
.B2(n_65),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_3),
.A2(n_47),
.B1(n_143),
.B2(n_210),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_70),
.B1(n_73),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_5),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_60),
.B1(n_65),
.B2(n_160),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_160),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_5),
.A2(n_27),
.B1(n_33),
.B2(n_160),
.Y(n_285)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_57),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_7),
.A2(n_27),
.B1(n_33),
.B2(n_57),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_8),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_34),
.B1(n_60),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_8),
.A2(n_34),
.B1(n_143),
.B2(n_210),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_38),
.B1(n_60),
.B2(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_38),
.B1(n_55),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_27),
.B1(n_33),
.B2(n_38),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_12),
.B(n_70),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_59),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_12),
.B(n_39),
.C(n_81),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_12),
.A2(n_60),
.B1(n_65),
.B2(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_12),
.B(n_124),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_211),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_27),
.C(n_43),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_12),
.A2(n_26),
.B(n_273),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_60),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_70),
.B1(n_71),
.B2(n_85),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_27),
.B1(n_33),
.B2(n_85),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_15),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_15),
.A2(n_60),
.B1(n_65),
.B2(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_72),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_15),
.A2(n_27),
.B1(n_33),
.B2(n_72),
.Y(n_243)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_350),
.B(n_353),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_345),
.B(n_349),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_332),
.B(n_344),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_134),
.A3(n_150),
.B(n_329),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_113),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_22),
.B(n_113),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_92),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_23),
.A2(n_76),
.B1(n_77),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_23),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_24),
.A2(n_25),
.B(n_51),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_25),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_25),
.A2(n_35),
.B1(n_36),
.B2(n_50),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_26),
.A2(n_32),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_26),
.A2(n_29),
.B1(n_97),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_26),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_26),
.A2(n_184),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_26),
.B(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_26),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_29),
.B(n_211),
.Y(n_297)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_33),
.B(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_37),
.A2(n_41),
.B1(n_48),
.B2(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_39),
.A2(n_40),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_39),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_41),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_41),
.A2(n_48),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_41),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_41),
.A2(n_48),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_45),
.A2(n_88),
.B1(n_103),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_45),
.A2(n_170),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_45),
.A2(n_206),
.B(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_45),
.B(n_211),
.Y(n_292)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_48),
.B(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_53),
.A2(n_58),
.B1(n_110),
.B2(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_73),
.Y(n_75)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_56),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_58),
.A2(n_110),
.B1(n_132),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_58),
.A2(n_67),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_74),
.B1(n_108),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_59),
.A2(n_74),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_59),
.A2(n_74),
.B1(n_340),
.B2(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_59),
.A2(n_74),
.B(n_347),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_65),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_60),
.B(n_66),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_60),
.B(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_63),
.A2(n_65),
.A3(n_73),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_74),
.A2(n_112),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_87),
.B(n_91),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_79),
.A2(n_80),
.B1(n_126),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_79),
.A2(n_177),
.B(n_179),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_79),
.A2(n_179),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_80),
.A2(n_105),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_80),
.A2(n_163),
.B(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_88),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_88),
.A2(n_261),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_92),
.A2(n_93),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.C(n_106),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_94),
.A2(n_95),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_99),
.A2(n_168),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_99),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_104),
.B(n_106),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B(n_111),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_116),
.C(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_131),
.B2(n_133),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_128),
.C(n_131),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_123),
.A2(n_124),
.B1(n_178),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_123),
.A2(n_124),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_164),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_128),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_128),
.B(n_141),
.C(n_147),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_131),
.B(n_137),
.C(n_140),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_135),
.A2(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_149),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_136),
.B(n_149),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_142),
.Y(n_339)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_148),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_322),
.B(n_328),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_195),
.B(n_321),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_188),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_153),
.B(n_188),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_171),
.C(n_173),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_154),
.A2(n_155),
.B1(n_171),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_171),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_173),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_176),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_180),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_182),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_190),
.B(n_191),
.C(n_194),
.Y(n_327)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_228),
.B(n_315),
.C(n_320),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_222),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_222),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_213),
.C(n_214),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_198),
.A2(n_199),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_204),
.C(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B(n_212),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_213),
.B(n_214),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_309),
.B(n_314),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_262),
.B(n_308),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_251),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_233),
.B(n_251),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.C(n_248),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_237),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B(n_242),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_241),
.A2(n_285),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_244),
.A2(n_248),
.B1(n_249),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_302),
.B(n_307),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_281),
.B(n_301),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_275),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_290),
.B(n_300),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_288),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_295),
.B(n_299),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_306),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_334),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_341),
.C(n_343),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_348),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_355),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);


endmodule