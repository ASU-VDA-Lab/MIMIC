module fake_jpeg_31575_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_265;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_156;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_34),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_63),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_35),
.B1(n_41),
.B2(n_29),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_72),
.B1(n_81),
.B2(n_88),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_31),
.C(n_20),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_82),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_71),
.B(n_85),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_35),
.B1(n_29),
.B2(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_29),
.B1(n_17),
.B2(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_78),
.B1(n_87),
.B2(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_77),
.B(n_79),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_18),
.B1(n_37),
.B2(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_28),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_18),
.B1(n_40),
.B2(n_36),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_0),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_90),
.B(n_92),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_19),
.B1(n_23),
.B2(n_37),
.Y(n_98)
);

NOR2x1_ASAP7_75t_R g103 ( 
.A(n_51),
.B(n_28),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_15),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_42),
.A2(n_23),
.B1(n_28),
.B2(n_3),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_115),
.B1(n_1),
.B2(n_15),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_42),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_11),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_11),
.B1(n_14),
.B2(n_3),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_114),
.B1(n_105),
.B2(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_9),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_12),
.B1(n_14),
.B2(n_3),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_126),
.B1(n_105),
.B2(n_106),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_127),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_135),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_107),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_75),
.Y(n_148)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_143),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_106),
.B1(n_109),
.B2(n_101),
.Y(n_167)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_82),
.B(n_89),
.C(n_84),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_93),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_89),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_160),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_70),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_105),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_129),
.B1(n_107),
.B2(n_127),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_96),
.B1(n_109),
.B2(n_101),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_122),
.B1(n_66),
.B2(n_130),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_140),
.B1(n_135),
.B2(n_143),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_171),
.B(n_179),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_91),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_93),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_102),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_102),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_91),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_66),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_126),
.B(n_66),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_100),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_121),
.B1(n_134),
.B2(n_128),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_185),
.B1(n_198),
.B2(n_164),
.Y(n_209)
);

NAND2x1_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_128),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_201),
.B(n_203),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_116),
.B1(n_74),
.B2(n_131),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_74),
.B1(n_123),
.B2(n_118),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_176),
.B1(n_151),
.B2(n_161),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_R g203 ( 
.A(n_150),
.B(n_75),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_133),
.B(n_139),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_178),
.B(n_177),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_212),
.B1(n_196),
.B2(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_149),
.B1(n_154),
.B2(n_151),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_152),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_153),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_160),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_225),
.C(n_193),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_224),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_149),
.C(n_157),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_189),
.C(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_233),
.C(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_235),
.B1(n_240),
.B2(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_182),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_191),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_195),
.C(n_194),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_190),
.C(n_181),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_203),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_242),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_183),
.B1(n_185),
.B2(n_149),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_190),
.C(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_198),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_213),
.B1(n_222),
.B2(n_211),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_248),
.B1(n_159),
.B2(n_169),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_244),
.B(n_231),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_249),
.B(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_243),
.B1(n_241),
.B2(n_237),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_223),
.B(n_225),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_223),
.A3(n_216),
.B1(n_227),
.B2(n_212),
.C1(n_221),
.C2(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_211),
.B(n_183),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_215),
.B(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_257),
.B1(n_192),
.B2(n_197),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_254),
.C(n_256),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_263),
.C(n_251),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_252),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_232),
.B1(n_233),
.B2(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_215),
.C(n_217),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_217),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_159),
.B(n_166),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_265),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_263),
.C(n_260),
.Y(n_279)
);

OAI21x1_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_248),
.B(n_169),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_278),
.B(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_280),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_259),
.C(n_262),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_272),
.B(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_264),
.C(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_271),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_279),
.C(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_271),
.B(n_169),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_202),
.C(n_156),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_292),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_202),
.Y(n_296)
);


endmodule