module fake_jpeg_18312_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_31),
.B1(n_20),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_54),
.B1(n_38),
.B2(n_44),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_41),
.B1(n_43),
.B2(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_44),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_31),
.B1(n_20),
.B2(n_24),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_22),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_54),
.C(n_47),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_60),
.B1(n_22),
.B2(n_37),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_65),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_63),
.A2(n_96),
.B(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_33),
.B1(n_41),
.B2(n_16),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_74),
.B1(n_76),
.B2(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_71),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_41),
.B1(n_27),
.B2(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_21),
.B1(n_27),
.B2(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_42),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_81),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_21),
.B1(n_30),
.B2(n_35),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_18),
.B1(n_38),
.B2(n_43),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_93),
.B1(n_44),
.B2(n_40),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_91),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_101),
.B1(n_102),
.B2(n_37),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_38),
.B1(n_30),
.B2(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_23),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_97),
.Y(n_128)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_40),
.B1(n_44),
.B2(n_29),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_42),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_100),
.Y(n_129)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_42),
.B1(n_40),
.B2(n_44),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_37),
.B(n_22),
.C(n_40),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_132),
.B(n_89),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_126),
.B1(n_95),
.B2(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_32),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_40),
.C(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_102),
.B1(n_101),
.B2(n_62),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_64),
.A2(n_44),
.B1(n_34),
.B2(n_17),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_89),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_71),
.Y(n_138)
);

AND2x4_ASAP7_75t_SL g132 ( 
.A(n_63),
.B(n_29),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_137),
.B1(n_143),
.B2(n_147),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_99),
.B1(n_86),
.B2(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_142),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_63),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_144),
.B(n_145),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_63),
.A3(n_93),
.B1(n_83),
.B2(n_23),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_23),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_109),
.A2(n_81),
.B1(n_79),
.B2(n_26),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_92),
.B(n_87),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_148),
.A2(n_108),
.B(n_128),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_32),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_153),
.Y(n_162)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_157),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_32),
.Y(n_153)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_104),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_89),
.B1(n_34),
.B2(n_17),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_126),
.B1(n_112),
.B2(n_125),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_34),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_111),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_163),
.B(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_114),
.B1(n_125),
.B2(n_122),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_188),
.B1(n_145),
.B2(n_140),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_103),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_131),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_120),
.C(n_133),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_105),
.C(n_34),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_104),
.B(n_108),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_130),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_105),
.B1(n_17),
.B2(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_148),
.B1(n_145),
.B2(n_113),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_114),
.B1(n_121),
.B2(n_115),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_118),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_119),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_127),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_106),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_0),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_205),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_202),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_212),
.B1(n_214),
.B2(n_179),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_140),
.B1(n_110),
.B2(n_141),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_204),
.B1(n_218),
.B2(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_144),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_209),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_159),
.B1(n_123),
.B2(n_113),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_193),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_202),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_170),
.C(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_217),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_225),
.Y(n_258)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_197),
.B(n_175),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_235),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_165),
.B(n_182),
.C(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_227),
.B1(n_213),
.B2(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_238),
.C(n_211),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_173),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_220),
.A2(n_173),
.B1(n_176),
.B2(n_164),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_166),
.C(n_164),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_218),
.B(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_199),
.B1(n_200),
.B2(n_220),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_179),
.B(n_189),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_219),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_259),
.B1(n_0),
.B2(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_230),
.B1(n_226),
.B2(n_237),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_228),
.C(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_260),
.C(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_192),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_221),
.B1(n_198),
.B2(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_206),
.C(n_203),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_194),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_226),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_269),
.C(n_276),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_226),
.B(n_230),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_252),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_201),
.B1(n_174),
.B2(n_192),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_201),
.B(n_229),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_275),
.B1(n_260),
.B2(n_261),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_174),
.B(n_6),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_248),
.B(n_259),
.C(n_11),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_262),
.CI(n_250),
.CON(n_283),
.SN(n_283)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_244),
.A2(n_5),
.B(n_12),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_263),
.B1(n_268),
.B2(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_257),
.C(n_10),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.C(n_3),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_281),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_266),
.C(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_278),
.C(n_279),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_273),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_293),
.B(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_294),
.C(n_295),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_278),
.B(n_288),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_280),
.B(n_284),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_306),
.B(n_301),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_280),
.B1(n_275),
.B2(n_11),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_302),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_307),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_1),
.Y(n_312)
);


endmodule