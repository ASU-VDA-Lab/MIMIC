module fake_jpeg_24029_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_59;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_22),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_4),
.B(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_5),
.B1(n_8),
.B2(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_39),
.B(n_13),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_44),
.B1(n_34),
.B2(n_39),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_10),
.B1(n_16),
.B2(n_19),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_16),
.B(n_19),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_49),
.B(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_33),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_14),
.B(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_33),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_56),
.C(n_38),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_30),
.C(n_29),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

AOI22x1_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_47),
.B1(n_38),
.B2(n_43),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_41),
.B1(n_43),
.B2(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_54),
.B1(n_52),
.B2(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_66),
.B1(n_62),
.B2(n_67),
.Y(n_69)
);

AO221x1_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_41),
.B1(n_35),
.B2(n_52),
.C(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_65),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_64),
.B(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_59),
.B(n_35),
.Y(n_74)
);


endmodule