module fake_jpeg_25715_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_20),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_29),
.B(n_26),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_15),
.C(n_14),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_64),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_46),
.B1(n_27),
.B2(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_16),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_27),
.B1(n_25),
.B2(n_33),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_46),
.B1(n_25),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_86),
.B1(n_48),
.B2(n_63),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_80),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_76),
.B1(n_78),
.B2(n_97),
.Y(n_109)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_73),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_28),
.B(n_26),
.C(n_21),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_87),
.B(n_24),
.C(n_33),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_79),
.Y(n_105)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_63),
.B1(n_43),
.B2(n_37),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_29),
.B1(n_30),
.B2(n_16),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_48),
.C(n_38),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_17),
.B(n_36),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_36),
.B(n_34),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_36),
.B(n_40),
.Y(n_102)
);

OR2x2_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_38),
.C(n_42),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_45),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_71),
.B1(n_68),
.B2(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_124),
.B1(n_92),
.B2(n_17),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_43),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_83),
.B(n_36),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_42),
.C(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_23),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_37),
.B1(n_41),
.B2(n_45),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_128),
.Y(n_158)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_33),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_30),
.B(n_24),
.C(n_31),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_136),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_137),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_91),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_73),
.B1(n_80),
.B2(n_76),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_151),
.B1(n_154),
.B2(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_93),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_174)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_88),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_9),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_106),
.B1(n_110),
.B2(n_115),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_168),
.B1(n_172),
.B2(n_40),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_114),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_164),
.B(n_173),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_117),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_98),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_119),
.B1(n_103),
.B2(n_108),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_115),
.B1(n_104),
.B2(n_103),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_181),
.B1(n_129),
.B2(n_146),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_118),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_120),
.B1(n_99),
.B2(n_126),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_99),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_182),
.B(n_31),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_183),
.B(n_186),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_90),
.B(n_94),
.C(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_90),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_134),
.B(n_45),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_128),
.B(n_45),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_144),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_138),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_204),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_138),
.C(n_31),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_200),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_45),
.B1(n_41),
.B2(n_42),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_168),
.B1(n_184),
.B2(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_218),
.B1(n_160),
.B2(n_157),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_23),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_40),
.C(n_18),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_207),
.C(n_213),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_18),
.C(n_35),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_23),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_163),
.B(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_22),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_31),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_22),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_159),
.B(n_22),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_162),
.A2(n_35),
.B1(n_22),
.B2(n_34),
.Y(n_218)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_162),
.B(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_162),
.B(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_190),
.B1(n_194),
.B2(n_203),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_200),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_238),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_167),
.B1(n_158),
.B2(n_181),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_239),
.B1(n_197),
.B2(n_219),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_166),
.B(n_165),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_166),
.B(n_164),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_235),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_164),
.B(n_186),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_164),
.C(n_180),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_157),
.C(n_159),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_8),
.B(n_15),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_10),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_207),
.C(n_191),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_253),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_197),
.CI(n_194),
.CON(n_250),
.SN(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_205),
.C(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_252),
.C(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_209),
.C(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_201),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_231),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_259),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_265),
.B1(n_241),
.B2(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_35),
.C(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_237),
.C(n_226),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_276),
.C(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_228),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_256),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_32),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_222),
.B1(n_221),
.B2(n_243),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_257),
.B1(n_262),
.B2(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_226),
.C(n_230),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_232),
.C(n_234),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_259),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_247),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_266),
.C(n_248),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_278),
.C(n_270),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

BUFx12f_ASAP7_75t_SL g287 ( 
.A(n_283),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_250),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.C(n_274),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_233),
.C(n_250),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_288),
.C(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_14),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_304),
.C(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_282),
.C(n_279),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_310),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_277),
.B(n_273),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_294),
.B(n_13),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_271),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_32),
.C(n_34),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_286),
.B1(n_295),
.B2(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_13),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_321),
.B(n_308),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_32),
.C(n_13),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_312),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_11),
.B(n_10),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_0),
.B(n_1),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_307),
.B1(n_303),
.B2(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_327),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_0),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_1),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_319),
.B(n_3),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_328),
.B(n_326),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_324),
.A3(n_329),
.B1(n_331),
.B2(n_5),
.C1(n_2),
.C2(n_7),
.Y(n_333)
);

AO21x2_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_2),
.B(n_3),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_317),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_4),
.B(n_5),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_4),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_6),
.B1(n_7),
.B2(n_317),
.Y(n_338)
);


endmodule