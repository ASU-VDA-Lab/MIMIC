module fake_jpeg_12946_n_393 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_51),
.B(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_58),
.Y(n_96)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_56),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_19),
.A2(n_12),
.B(n_8),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_63),
.Y(n_87)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_0),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_8),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_79),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_1),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_84),
.Y(n_130)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_26),
.B1(n_39),
.B2(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_86),
.A2(n_93),
.B1(n_131),
.B2(n_132),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_26),
.B1(n_41),
.B2(n_39),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_92),
.A2(n_97),
.B1(n_103),
.B2(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_39),
.B1(n_35),
.B2(n_38),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_35),
.B1(n_42),
.B2(n_32),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_95),
.A2(n_110),
.B1(n_113),
.B2(n_127),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_33),
.B1(n_38),
.B2(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_36),
.B1(n_34),
.B2(n_42),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_24),
.CON(n_106),
.SN(n_106)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_120),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_55),
.A2(n_32),
.B1(n_28),
.B2(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_34),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_28),
.B1(n_20),
.B2(n_24),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_1),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_84),
.B1(n_67),
.B2(n_54),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_5),
.B1(n_6),
.B2(n_88),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_3),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_89),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_45),
.B(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_72),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_48),
.A2(n_5),
.B1(n_6),
.B2(n_78),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_52),
.A2(n_75),
.B1(n_77),
.B2(n_73),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_47),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_136),
.B(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_69),
.B1(n_68),
.B2(n_49),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_140),
.A2(n_143),
.B1(n_145),
.B2(n_144),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_157),
.Y(n_220)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_56),
.B1(n_62),
.B2(n_70),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_6),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_106),
.B1(n_111),
.B2(n_120),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_93),
.B1(n_121),
.B2(n_86),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_151),
.A2(n_165),
.B(n_156),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_107),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_115),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_94),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_109),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_117),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_89),
.Y(n_173)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_108),
.Y(n_175)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_108),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_179),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_89),
.A2(n_100),
.B1(n_118),
.B2(n_98),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_91),
.B1(n_173),
.B2(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_117),
.B(n_109),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_144),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_195),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_99),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_189),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_99),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_158),
.B1(n_180),
.B2(n_150),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_156),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_140),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_167),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_91),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_151),
.A2(n_135),
.B1(n_139),
.B2(n_158),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_138),
.B1(n_174),
.B2(n_163),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_138),
.B(n_137),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_135),
.B(n_166),
.C(n_143),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_222),
.A2(n_212),
.B(n_218),
.C(n_181),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_157),
.B(n_170),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_225),
.A2(n_253),
.B(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_229),
.A2(n_251),
.B(n_253),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_248),
.Y(n_271)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_192),
.B(n_162),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_171),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_181),
.C(n_189),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_142),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_168),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_194),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_247),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_169),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_164),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_207),
.B(n_163),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_252),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_163),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_200),
.B(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_238),
.Y(n_302)
);

AOI22x1_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_222),
.B1(n_226),
.B2(n_205),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_206),
.A3(n_214),
.B1(n_198),
.B2(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_181),
.B1(n_195),
.B2(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_238),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_222),
.A2(n_199),
.B1(n_196),
.B2(n_186),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_282),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_191),
.B(n_201),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_248),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_199),
.C(n_203),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_286),
.C(n_253),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_223),
.A2(n_191),
.B(n_202),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_203),
.C(n_201),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_245),
.C(n_240),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_302),
.C(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_299),
.B(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_242),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_301),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_251),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_303),
.B(n_308),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_222),
.B1(n_252),
.B2(n_239),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_306),
.A2(n_271),
.B1(n_282),
.B2(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_254),
.C(n_197),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_188),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_262),
.C(n_257),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_311),
.Y(n_330)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_268),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_328),
.C(n_289),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_283),
.B1(n_262),
.B2(n_273),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_319),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_297),
.A2(n_274),
.B(n_284),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_271),
.B(n_290),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_293),
.B1(n_297),
.B2(n_307),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_262),
.B1(n_285),
.B2(n_257),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_277),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_260),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_333),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_260),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_SL g334 ( 
.A1(n_331),
.A2(n_295),
.A3(n_288),
.B1(n_264),
.B2(n_301),
.C1(n_292),
.C2(n_306),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_337),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_302),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_340),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_SL g337 ( 
.A(n_328),
.B(n_288),
.C(n_303),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_342),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_323),
.A2(n_307),
.B1(n_262),
.B2(n_294),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_309),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_314),
.B(n_284),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_326),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_263),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_345),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_327),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_308),
.C(n_300),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_349),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_267),
.C(n_275),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_320),
.C(n_332),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_313),
.B(n_277),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_322),
.B1(n_317),
.B2(n_318),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_357),
.C(n_335),
.Y(n_364)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_359),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_315),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_358),
.B(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_362),
.A2(n_315),
.B(n_275),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_325),
.B1(n_316),
.B2(n_321),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_363),
.A2(n_259),
.B(n_250),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_371),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_351),
.A2(n_339),
.B(n_329),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_365),
.A2(n_366),
.B(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_368),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_336),
.C(n_340),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_352),
.A2(n_341),
.B(n_296),
.Y(n_369)
);

OAI32xp33_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_325),
.A3(n_269),
.B1(n_256),
.B2(n_231),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_269),
.C(n_259),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_356),
.C(n_362),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_358),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_379),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_354),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_355),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_380),
.B(n_357),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_355),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_383),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_375),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_235),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_377),
.B(n_380),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_386),
.A2(n_388),
.B1(n_381),
.B2(n_382),
.Y(n_389)
);

AOI321xp33_ASAP7_75t_SL g391 ( 
.A1(n_389),
.A2(n_390),
.A3(n_205),
.B1(n_193),
.B2(n_202),
.C(n_210),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_210),
.B1(n_183),
.B2(n_188),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_193),
.C(n_209),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_209),
.Y(n_393)
);


endmodule