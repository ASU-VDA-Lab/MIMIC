module fake_netlist_6_4725_n_1751 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1751);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1751;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_85),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_46),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_60),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_50),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_79),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_28),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_149),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_67),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_139),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_46),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_44),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_125),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_101),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_40),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_13),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_0),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_120),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_164),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_113),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_84),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_47),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_37),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_32),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_89),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_29),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_12),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_94),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_53),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_23),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_91),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_61),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_82),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_37),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_51),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_45),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_119),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_159),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_137),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_70),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_77),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_27),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_166),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_124),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_136),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_152),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_80),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_5),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_74),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_155),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_54),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_76),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_3),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_48),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_0),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_68),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_133),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_81),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_160),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_58),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_7),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_35),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_27),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_112),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_47),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_147),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_23),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_20),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_162),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_168),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_59),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_123),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_172),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_95),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_48),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_56),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_154),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_50),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_65),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_78),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_45),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_170),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_161),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_40),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_39),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_42),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_43),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_104),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_26),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_158),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_2),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_52),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_96),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_54),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_22),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_102),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_42),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_64),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_156),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_17),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_14),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_51),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_49),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_31),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_49),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_141),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_13),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_17),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_148),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_100),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_15),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_41),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_6),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_97),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_16),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_140),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_114),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_11),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_179),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_240),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_240),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_240),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_240),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_240),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_213),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_333),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_246),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_246),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_246),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_246),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_246),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_219),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_222),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_228),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_267),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_294),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_182),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_231),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_234),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_237),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_203),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_193),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_220),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_238),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_175),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_241),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_248),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_224),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_193),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_195),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_267),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_175),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_183),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_278),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_249),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_205),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_206),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_183),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_214),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_229),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_269),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_189),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_278),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_250),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_252),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_284),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_254),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_243),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_245),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_271),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_272),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_287),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_298),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_299),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_305),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_189),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_313),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_325),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_255),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_225),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_312),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_197),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_197),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_211),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_225),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_317),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_211),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_256),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_312),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_353),
.B(n_186),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

BUFx8_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_431),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_201),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_358),
.B(n_201),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_361),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_173),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_417),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_359),
.B(n_186),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_355),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_226),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_173),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_367),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_351),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_357),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_362),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_362),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_364),
.B(n_226),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_397),
.B(n_198),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_374),
.B(n_230),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

AOI22x1_ASAP7_75t_SL g474 ( 
.A1(n_384),
.A2(n_273),
.B1(n_264),
.B2(n_332),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_366),
.B(n_174),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_359),
.B(n_317),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_366),
.B(n_230),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_370),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_360),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_368),
.B(n_259),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_371),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_380),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_372),
.B(n_277),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_373),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_374),
.B(n_174),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_396),
.B(n_176),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_369),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

NAND2x1_ASAP7_75t_L g498 ( 
.A(n_400),
.B(n_277),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_401),
.A2(n_301),
.B(n_289),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_356),
.A2(n_244),
.B1(n_347),
.B2(n_321),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_375),
.B(n_178),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_403),
.A2(n_301),
.B(n_289),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_386),
.A2(n_321),
.B1(n_331),
.B2(n_332),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_378),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_363),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_334),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_376),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_411),
.Y(n_515)
);

AND3x2_ASAP7_75t_L g516 ( 
.A(n_470),
.B(n_394),
.C(n_377),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_470),
.B(n_381),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_499),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_439),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_440),
.A2(n_437),
.B1(n_402),
.B2(n_423),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_464),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_455),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_457),
.B(n_382),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_442),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_499),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_439),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_456),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_457),
.B(n_383),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_387),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_456),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_457),
.B(n_389),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_453),
.B(n_390),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_481),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_440),
.A2(n_434),
.B1(n_414),
.B2(n_375),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_480),
.B(n_399),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_453),
.B(n_409),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_462),
.B(n_410),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_440),
.A2(n_411),
.B1(n_415),
.B2(n_416),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_447),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_452),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_460),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_460),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_462),
.B(n_413),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_448),
.B(n_428),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_454),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_449),
.B(n_438),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_454),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_R g561 ( 
.A(n_463),
.B(n_514),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_476),
.B(n_406),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_476),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_448),
.B(n_239),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_446),
.B(n_483),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_508),
.A2(n_335),
.B1(n_339),
.B2(n_341),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_472),
.B(n_416),
.C(n_415),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_445),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_300),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_459),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_499),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_459),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_472),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_509),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_430),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

AND2x2_ASAP7_75t_SL g585 ( 
.A(n_500),
.B(n_177),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_446),
.B(n_483),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_446),
.B(n_194),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

NOR3xp33_ASAP7_75t_L g589 ( 
.A(n_502),
.B(n_320),
.C(n_223),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_467),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_463),
.B(n_391),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_472),
.B(n_430),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_247),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_467),
.Y(n_599)
);

BUFx4f_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_473),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_445),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_471),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_507),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_513),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_473),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_493),
.B(n_339),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_473),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_469),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_446),
.B(n_194),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_475),
.B(n_260),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_507),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_451),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

AO21x2_ASAP7_75t_L g618 ( 
.A1(n_493),
.A2(n_188),
.B(n_187),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_486),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_412),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_486),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_509),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_435),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_498),
.B(n_207),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_510),
.B(n_435),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

BUFx8_ASAP7_75t_SL g627 ( 
.A(n_474),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_510),
.B(n_515),
.Y(n_628)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_500),
.A2(n_216),
.B(n_215),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_515),
.B(n_261),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_SL g631 ( 
.A1(n_484),
.A2(n_436),
.B(n_419),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_498),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_486),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_486),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_505),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_505),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_469),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_466),
.B(n_266),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_505),
.A2(n_257),
.B(n_253),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_469),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_461),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_469),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_477),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_451),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_466),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_466),
.B(n_279),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_477),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_466),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_494),
.B(n_281),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_499),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_499),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_494),
.B(n_282),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_451),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_484),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_511),
.B(n_436),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_503),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_640),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_546),
.B(n_503),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_555),
.B(n_503),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_571),
.B(n_503),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_664),
.B(n_178),
.Y(n_672)
);

NOR2x1p5_ASAP7_75t_L g673 ( 
.A(n_541),
.B(n_579),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_563),
.B(n_511),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_556),
.B(n_503),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_L g676 ( 
.A(n_559),
.B(n_502),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_503),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_563),
.B(n_180),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_520),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_598),
.B(n_503),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_622),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_598),
.B(n_505),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_598),
.B(n_505),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_598),
.B(n_443),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_585),
.B(n_272),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_623),
.A2(n_640),
.B(n_645),
.C(n_643),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_527),
.B(n_532),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_614),
.B(n_443),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_624),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_664),
.B(n_180),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_538),
.B(n_181),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_533),
.B(n_451),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_520),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_181),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_594),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_530),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_664),
.B(n_184),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_530),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_537),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_643),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_600),
.A2(n_490),
.B(n_497),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_585),
.B(n_272),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_585),
.B(n_600),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_634),
.B(n_272),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_570),
.B(n_485),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_517),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_645),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_600),
.B(n_272),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_639),
.B(n_490),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_485),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_606),
.B(n_488),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_647),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_517),
.B(n_488),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_647),
.B(n_497),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_648),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_569),
.B(n_489),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_664),
.B(n_184),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_648),
.B(n_512),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_649),
.B(n_512),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_523),
.B(n_185),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_649),
.B(n_512),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_620),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_554),
.B(n_185),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_581),
.B(n_190),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_554),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_548),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_544),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_542),
.B(n_227),
.C(n_217),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_597),
.B(n_272),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_540),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_549),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_581),
.B(n_190),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_653),
.B(n_497),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_665),
.B(n_191),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_653),
.B(n_506),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_656),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_557),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_597),
.A2(n_295),
.B1(n_297),
.B2(n_283),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_618),
.A2(n_342),
.B1(n_349),
.B2(n_263),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_549),
.B(n_506),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_631),
.A2(n_501),
.B(n_489),
.C(n_492),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_492),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_552),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_536),
.B(n_501),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_268),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_558),
.B(n_309),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_558),
.B(n_329),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_597),
.B(n_272),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_539),
.B(n_191),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_625),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_560),
.B(n_330),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_589),
.B(n_242),
.C(n_236),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_625),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_560),
.B(n_478),
.Y(n_755)
);

AOI221xp5_ASAP7_75t_L g756 ( 
.A1(n_651),
.A2(n_341),
.B1(n_343),
.B2(n_345),
.C(n_258),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_272),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_618),
.A2(n_461),
.B1(n_221),
.B2(n_262),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_565),
.B(n_478),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_547),
.B(n_192),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_633),
.B(n_291),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_543),
.B(n_192),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_565),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_573),
.B(n_478),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_573),
.B(n_479),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_583),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_633),
.B(n_292),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_583),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_544),
.B(n_196),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_584),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_595),
.B(n_418),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_609),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_603),
.B(n_420),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_584),
.B(n_479),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_593),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_544),
.B(n_421),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_593),
.B(n_479),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_561),
.B(n_567),
.C(n_569),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_599),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_630),
.A2(n_308),
.B1(n_296),
.B2(n_303),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_611),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_618),
.A2(n_306),
.B1(n_311),
.B2(n_348),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_544),
.B(n_196),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_601),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_611),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_601),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_562),
.A2(n_323),
.B1(n_200),
.B2(n_202),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_604),
.Y(n_788)
);

BUFx5_ASAP7_75t_L g789 ( 
.A(n_633),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_604),
.B(n_199),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_605),
.B(n_482),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_608),
.B(n_613),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_611),
.B(n_199),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_658),
.B(n_662),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_587),
.B(n_200),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_521),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_608),
.B(n_482),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_622),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_522),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_631),
.A2(n_421),
.B(n_422),
.C(n_424),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_612),
.B(n_202),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_613),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_615),
.B(n_487),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_615),
.B(n_487),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_617),
.B(n_626),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_516),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_641),
.A2(n_340),
.B1(n_204),
.B2(n_208),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_522),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_638),
.A2(n_461),
.B1(n_221),
.B2(n_262),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_617),
.B(n_487),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_626),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_635),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_635),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_638),
.B(n_491),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_628),
.B(n_655),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_638),
.B(n_204),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_524),
.B(n_491),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_528),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_624),
.A2(n_348),
.B1(n_208),
.B2(n_327),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_528),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_624),
.A2(n_318),
.B1(n_209),
.B2(n_210),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_524),
.B(n_496),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_624),
.A2(n_461),
.B1(n_221),
.B2(n_194),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_524),
.B(n_535),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_590),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_624),
.A2(n_209),
.B1(n_210),
.B2(n_340),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_524),
.B(n_535),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_654),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_525),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_697),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_798),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_668),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_SL g833 ( 
.A1(n_735),
.A2(n_474),
.B1(n_345),
.B2(n_262),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_697),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_735),
.B(n_535),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_687),
.A2(n_566),
.B1(n_586),
.B2(n_579),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_679),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_789),
.B(n_654),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_751),
.B(n_535),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_687),
.A2(n_661),
.B1(n_660),
.B2(n_659),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_754),
.B(n_576),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_SL g843 ( 
.A(n_694),
.B(n_723),
.C(n_801),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_785),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_798),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_728),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_704),
.A2(n_661),
.B1(n_660),
.B2(n_659),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_708),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_785),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_713),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_785),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_679),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_SL g853 ( 
.A1(n_695),
.A2(n_288),
.B1(n_232),
.B2(n_233),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_789),
.B(n_657),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_816),
.B(n_576),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_816),
.B(n_576),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_723),
.B(n_674),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_763),
.B(n_576),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_SL g859 ( 
.A1(n_750),
.A2(n_669),
.B(n_670),
.C(n_666),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_693),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_728),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_745),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_766),
.B(n_657),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_716),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_681),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_776),
.B(n_567),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_801),
.A2(n_286),
.B1(n_251),
.B2(n_265),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_789),
.B(n_619),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_696),
.Y(n_869)
);

OR2x2_ASAP7_75t_SL g870 ( 
.A(n_778),
.B(n_729),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_829),
.B(n_689),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_737),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_699),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_768),
.B(n_526),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_674),
.B(n_519),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_727),
.B(n_425),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_770),
.B(n_526),
.Y(n_877)
);

NOR2x2_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_627),
.Y(n_878)
);

AO22x1_ASAP7_75t_L g879 ( 
.A1(n_694),
.A2(n_290),
.B1(n_270),
.B2(n_274),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_711),
.B(n_577),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_682),
.A2(n_683),
.B(n_680),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_727),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_784),
.B(n_526),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_700),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_773),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_712),
.B(n_425),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_789),
.B(n_529),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_789),
.B(n_619),
.Y(n_888)
);

AND2x4_ASAP7_75t_SL g889 ( 
.A(n_726),
.B(n_663),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_738),
.Y(n_890)
);

INVx6_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_704),
.A2(n_621),
.B1(n_652),
.B2(n_632),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_676),
.B(n_725),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_725),
.B(n_733),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_731),
.B(n_568),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_691),
.A2(n_621),
.B1(n_652),
.B2(n_632),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_707),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_732),
.B(n_568),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_753),
.B(n_337),
.C(n_318),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_707),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_685),
.A2(n_534),
.B1(n_531),
.B2(n_550),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_673),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_732),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_714),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_785),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_689),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_744),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_744),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_714),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_775),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_691),
.A2(n_636),
.B1(n_637),
.B2(n_646),
.Y(n_911)
);

AND2x6_ASAP7_75t_SL g912 ( 
.A(n_762),
.B(n_426),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_775),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_667),
.B(n_519),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_733),
.B(n_519),
.Y(n_915)
);

AO22x1_ASAP7_75t_L g916 ( 
.A1(n_762),
.A2(n_750),
.B1(n_772),
.B2(n_806),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_779),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_786),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_786),
.B(n_572),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_689),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_761),
.A2(n_767),
.B1(n_743),
.B2(n_714),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_678),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_743),
.B(n_771),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_743),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_771),
.Y(n_925)
);

AND2x6_ASAP7_75t_L g926 ( 
.A(n_667),
.B(n_663),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_789),
.B(n_636),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

AND2x2_ASAP7_75t_SL g929 ( 
.A(n_758),
.B(n_519),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_771),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_717),
.B(n_574),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_790),
.B(n_574),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_706),
.B(n_426),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_724),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_688),
.B(n_637),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_802),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_825),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_675),
.B(n_646),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_678),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_781),
.B(n_427),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_811),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_781),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_SL g943 ( 
.A1(n_787),
.A2(n_285),
.B1(n_275),
.B2(n_316),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_686),
.A2(n_642),
.B1(n_629),
.B2(n_346),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_814),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_742),
.B(n_427),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_685),
.A2(n_703),
.B1(n_740),
.B2(n_730),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_790),
.B(n_574),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_812),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_684),
.B(n_529),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_813),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_746),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_671),
.B(n_529),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_761),
.A2(n_588),
.B1(n_575),
.B2(n_650),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_677),
.B(n_578),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_710),
.B(n_578),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_824),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_828),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_703),
.A2(n_730),
.B1(n_749),
.B2(n_739),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_749),
.A2(n_551),
.B1(n_531),
.B2(n_534),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_692),
.B(n_578),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_702),
.B(n_529),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_747),
.B(n_578),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_792),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_741),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_819),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_756),
.A2(n_551),
.B1(n_550),
.B2(n_553),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_815),
.A2(n_588),
.B(n_575),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_705),
.B(n_629),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_796),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_805),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_755),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_809),
.A2(n_346),
.B1(n_323),
.B2(n_337),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_826),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_782),
.A2(n_575),
.B1(n_588),
.B2(n_616),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_748),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_794),
.A2(n_529),
.B(n_616),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_752),
.B(n_580),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_715),
.B(n_580),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_799),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_719),
.B(n_580),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_800),
.A2(n_590),
.B(n_602),
.C(n_610),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_808),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_709),
.B(n_580),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_769),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_720),
.B(n_722),
.Y(n_987)
);

INVx5_ASAP7_75t_L g988 ( 
.A(n_808),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_734),
.A2(n_591),
.B1(n_553),
.B2(n_592),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_818),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_736),
.Y(n_991)
);

AND2x6_ASAP7_75t_SL g992 ( 
.A(n_759),
.B(n_429),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_820),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_721),
.B(n_276),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_820),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_SL g996 ( 
.A(n_793),
.B(n_644),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_764),
.B(n_582),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_807),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_817),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_795),
.B(n_582),
.Y(n_1000)
);

AO22x1_ASAP7_75t_L g1001 ( 
.A1(n_821),
.A2(n_293),
.B1(n_280),
.B2(n_304),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_822),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_873),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_843),
.A2(n_718),
.B(n_672),
.C(n_690),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_857),
.B(n_698),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_857),
.B(n_765),
.Y(n_1006)
);

AOI33xp33_ASAP7_75t_L g1007 ( 
.A1(n_833),
.A2(n_823),
.A3(n_780),
.B1(n_496),
.B2(n_315),
.B3(n_310),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_906),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_906),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_894),
.B(n_774),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_937),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_884),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_881),
.A2(n_945),
.B(n_856),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_906),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_893),
.B(n_777),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_882),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_947),
.A2(n_827),
.B1(n_760),
.B2(n_804),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_890),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_971),
.B(n_783),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_947),
.A2(n_810),
.B1(n_803),
.B2(n_797),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_843),
.A2(n_327),
.B1(n_791),
.B2(n_307),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_968),
.A2(n_650),
.B(n_582),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_945),
.A2(n_757),
.B(n_644),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_922),
.B(n_616),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_855),
.A2(n_644),
.B(n_650),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_922),
.B(n_616),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_875),
.A2(n_461),
.B1(n_610),
.B2(n_607),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_939),
.B(n_923),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_961),
.A2(n_644),
.B(n_602),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_890),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_907),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_902),
.B(n_2),
.C(n_4),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_923),
.B(n_591),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_865),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_962),
.A2(n_644),
.B(n_602),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_939),
.B(n_596),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_838),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_925),
.B(n_644),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_866),
.B(n_4),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_845),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_906),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_925),
.B(n_169),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_852),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_991),
.B(n_880),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_849),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_910),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_886),
.B(n_5),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_966),
.A2(n_461),
.B1(n_8),
.B2(n_9),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_930),
.B(n_165),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_862),
.B(n_6),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_899),
.A2(n_9),
.B(n_12),
.C(n_15),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_952),
.B(n_461),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_959),
.A2(n_62),
.B1(n_157),
.B2(n_153),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_831),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_861),
.B(n_145),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_913),
.Y(n_1058)
);

OAI22x1_ASAP7_75t_L g1059 ( 
.A1(n_837),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_885),
.B(n_18),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_846),
.B(n_143),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_917),
.Y(n_1062)
);

BUFx4f_ASAP7_75t_L g1063 ( 
.A(n_861),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_976),
.B(n_461),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_998),
.B(n_19),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_928),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_930),
.B(n_130),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_915),
.B(n_21),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_915),
.B(n_21),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_25),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_921),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_832),
.B(n_30),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_836),
.B(n_31),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_951),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_860),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_861),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_848),
.B(n_33),
.Y(n_1077)
);

INVx6_ASAP7_75t_L g1078 ( 
.A(n_876),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_912),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_924),
.B(n_86),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_924),
.B(n_871),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_849),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_869),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_850),
.A2(n_73),
.B1(n_117),
.B2(n_116),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_920),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_903),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_899),
.A2(n_973),
.B(n_986),
.C(n_994),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_987),
.A2(n_108),
.B(n_105),
.Y(n_1088)
);

AOI222xp33_ASAP7_75t_L g1089 ( 
.A1(n_974),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.C1(n_43),
.C2(n_52),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_920),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_864),
.A2(n_93),
.B1(n_53),
.B2(n_55),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_918),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_859),
.A2(n_38),
.B(n_55),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_951),
.B(n_56),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_959),
.A2(n_57),
.B1(n_870),
.B2(n_835),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_849),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_872),
.A2(n_946),
.B1(n_964),
.B2(n_904),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_965),
.B(n_972),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_SL g1099 ( 
.A1(n_929),
.A2(n_948),
.B(n_932),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_981),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_871),
.B(n_920),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_940),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_934),
.B(n_904),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_955),
.A2(n_956),
.B(n_914),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_940),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_946),
.A2(n_909),
.B(n_935),
.C(n_933),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_933),
.B(n_853),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_867),
.A2(n_941),
.B(n_949),
.C(n_936),
.Y(n_1108)
);

OAI22x1_ASAP7_75t_L g1109 ( 
.A1(n_830),
.A2(n_834),
.B1(n_900),
.B2(n_897),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_935),
.B(n_953),
.Y(n_1110)
);

AO21x1_ASAP7_75t_L g1111 ( 
.A1(n_950),
.A2(n_953),
.B(n_944),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_992),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_891),
.B(n_830),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_943),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_970),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_891),
.B(n_834),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_979),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_946),
.A2(n_958),
.B(n_840),
.C(n_842),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_914),
.A2(n_888),
.B(n_927),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_965),
.B(n_972),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_858),
.A2(n_863),
.B(n_936),
.C(n_941),
.Y(n_1121)
);

INVxp67_ASAP7_75t_R g1122 ( 
.A(n_984),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_949),
.A2(n_883),
.B(n_877),
.C(n_874),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_916),
.B(n_879),
.C(n_964),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_871),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_851),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_964),
.B(n_1002),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_990),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_999),
.B(n_900),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_851),
.B(n_905),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_929),
.A2(n_1000),
.B(n_841),
.C(n_983),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1000),
.A2(n_983),
.B(n_847),
.C(n_931),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_997),
.A2(n_985),
.B(n_938),
.C(n_963),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_851),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_851),
.B(n_905),
.Y(n_1135)
);

CKINVDCx11_ASAP7_75t_R g1136 ( 
.A(n_878),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_891),
.B(n_905),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_897),
.A2(n_905),
.B1(n_975),
.B2(n_957),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1001),
.B(n_889),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_957),
.A2(n_844),
.B1(n_988),
.B2(n_942),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_868),
.A2(n_839),
.B(n_854),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_997),
.A2(n_985),
.B(n_938),
.C(n_978),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_957),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_993),
.B(n_995),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1006),
.B(n_1010),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1016),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_SL g1147 ( 
.A(n_1089),
.B(n_967),
.C(n_896),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1013),
.A2(n_982),
.B(n_980),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1046),
.B(n_967),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1111),
.A2(n_1131),
.A3(n_1132),
.B(n_1095),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1040),
.B(n_911),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_1034),
.B(n_977),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1114),
.A2(n_996),
.B1(n_942),
.B2(n_926),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1099),
.A2(n_892),
.B(n_901),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1022),
.A2(n_1119),
.B(n_1141),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1015),
.A2(n_988),
.B(n_895),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1068),
.A2(n_898),
.B(n_919),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1005),
.B(n_989),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1100),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1110),
.A2(n_969),
.B(n_954),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1041),
.B(n_960),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1127),
.B(n_1098),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1020),
.A2(n_926),
.A3(n_960),
.B(n_989),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1008),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1019),
.B(n_926),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1069),
.A2(n_926),
.B(n_1118),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1128),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1097),
.A2(n_1091),
.B1(n_1065),
.B2(n_1143),
.Y(n_1168)
);

CKINVDCx8_ASAP7_75t_R g1169 ( 
.A(n_1112),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1003),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1035),
.A2(n_1025),
.B(n_1133),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1041),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1120),
.B(n_1037),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1012),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1123),
.A2(n_1142),
.B(n_1017),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1029),
.A2(n_1138),
.B(n_1121),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1018),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1023),
.A2(n_1140),
.B(n_1106),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1097),
.A2(n_1091),
.B1(n_1108),
.B2(n_1050),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1049),
.B(n_1102),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1093),
.A2(n_1027),
.B(n_1124),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1136),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1129),
.B(n_1024),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1088),
.A2(n_1027),
.B(n_1135),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1036),
.B(n_1048),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1058),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1030),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1062),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1130),
.A2(n_1055),
.B(n_1066),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1137),
.A2(n_1004),
.B(n_1087),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1144),
.B(n_1038),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1045),
.B(n_1075),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_1125),
.B(n_1107),
.Y(n_1195)
);

NOR4xp25_ASAP7_75t_L g1196 ( 
.A(n_1053),
.B(n_1071),
.C(n_1074),
.D(n_1007),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1137),
.A2(n_1080),
.B(n_1028),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1083),
.B(n_1092),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1105),
.B(n_1070),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1086),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1078),
.A2(n_1094),
.B1(n_1139),
.B2(n_1103),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1137),
.A2(n_1057),
.B(n_1084),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1063),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1109),
.A2(n_1059),
.A3(n_1077),
.B(n_1073),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1008),
.Y(n_1206)
);

NOR4xp25_ASAP7_75t_L g1207 ( 
.A(n_1021),
.B(n_1089),
.C(n_1072),
.D(n_1067),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1039),
.A2(n_1084),
.B(n_1054),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1079),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1115),
.A2(n_1117),
.B(n_1082),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1033),
.B(n_1096),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1033),
.B(n_1096),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1044),
.A2(n_1051),
.B1(n_1060),
.B2(n_1052),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1032),
.B(n_1064),
.C(n_1057),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1122),
.B(n_1078),
.Y(n_1215)
);

CKINVDCx8_ASAP7_75t_R g1216 ( 
.A(n_1009),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1047),
.B(n_1082),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1047),
.A2(n_1134),
.B(n_1126),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1126),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1134),
.A2(n_1126),
.B(n_1057),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1009),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1014),
.C(n_1042),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1014),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1009),
.A2(n_1090),
.B1(n_1042),
.B2(n_1043),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1076),
.B(n_1014),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1042),
.A2(n_1043),
.B(n_1085),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1043),
.B(n_1085),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1085),
.A2(n_1090),
.B(n_1061),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1004),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1005),
.B(n_544),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1008),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1136),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1022),
.A2(n_1119),
.B(n_1141),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1040),
.B(n_866),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1004),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1100),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1013),
.A2(n_887),
.B(n_859),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1004),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1013),
.A2(n_1111),
.B(n_1131),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_R g1242 ( 
.A(n_1016),
.B(n_464),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1013),
.A2(n_887),
.B(n_1104),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1022),
.A2(n_1119),
.B(n_1141),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1013),
.A2(n_1111),
.B(n_1131),
.Y(n_1245)
);

BUFx2_ASAP7_75t_SL g1246 ( 
.A(n_1008),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1006),
.A2(n_857),
.B1(n_735),
.B2(n_894),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1004),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_R g1249 ( 
.A(n_1016),
.B(n_464),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1016),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1034),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1016),
.Y(n_1252)
);

O2A1O1Ixp5_ASAP7_75t_L g1253 ( 
.A1(n_1068),
.A2(n_894),
.B(n_857),
.C(n_916),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1008),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_857),
.B(n_893),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1013),
.A2(n_887),
.B(n_1104),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1013),
.A2(n_1111),
.B(n_1131),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1100),
.Y(n_1258)
);

NOR2x1_ASAP7_75t_SL g1259 ( 
.A(n_1137),
.B(n_849),
.Y(n_1259)
);

NAND2x1p5_ASAP7_75t_L g1260 ( 
.A(n_1134),
.B(n_844),
.Y(n_1260)
);

NAND3x1_ASAP7_75t_L g1261 ( 
.A(n_1065),
.B(n_567),
.C(n_1040),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1005),
.B(n_857),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1004),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1006),
.B(n_857),
.Y(n_1264)
);

O2A1O1Ixp5_ASAP7_75t_L g1265 ( 
.A1(n_1068),
.A2(n_894),
.B(n_857),
.C(n_916),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1100),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1006),
.B(n_857),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1011),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1006),
.B(n_857),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1013),
.A2(n_887),
.B(n_1104),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1046),
.B(n_525),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1111),
.A2(n_1131),
.A3(n_1013),
.B(n_1132),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1041),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1016),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1006),
.B(n_857),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1013),
.A2(n_887),
.B(n_859),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1006),
.A2(n_857),
.B1(n_735),
.B2(n_894),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1013),
.A2(n_1111),
.B(n_1131),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1008),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1184),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1235),
.B(n_1151),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1247),
.A2(n_1279),
.B(n_1236),
.C(n_1248),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1184),
.B(n_1200),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1262),
.B(n_1145),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1231),
.A2(n_1278),
.B(n_1239),
.Y(n_1287)
);

NAND2x1_ASAP7_75t_L g1288 ( 
.A(n_1203),
.B(n_1219),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1187),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1187),
.Y(n_1290)
);

AO21x1_ASAP7_75t_L g1291 ( 
.A1(n_1247),
.A2(n_1279),
.B(n_1179),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1252),
.B(n_1273),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1199),
.B(n_1180),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1278),
.A2(n_1176),
.B(n_1171),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1251),
.Y(n_1295)
);

BUFx4_ASAP7_75t_SL g1296 ( 
.A(n_1146),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1167),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1255),
.A2(n_1272),
.B(n_1154),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1261),
.A2(n_1240),
.B(n_1230),
.Y(n_1299)
);

OAI21xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1145),
.A2(n_1269),
.B(n_1264),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1200),
.B(n_1238),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1255),
.A2(n_1178),
.B(n_1154),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1207),
.A2(n_1147),
.B1(n_1196),
.B2(n_1179),
.C(n_1263),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1217),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1170),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1238),
.B(n_1266),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1192),
.A2(n_1148),
.B(n_1166),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1162),
.B(n_1173),
.Y(n_1308)
);

NAND2x1_ASAP7_75t_L g1309 ( 
.A(n_1219),
.B(n_1197),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1310)
);

BUFx8_ASAP7_75t_SL g1311 ( 
.A(n_1233),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1253),
.A2(n_1265),
.B(n_1157),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1174),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1207),
.B(n_1168),
.C(n_1214),
.Y(n_1314)
);

AOI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_1221),
.B1(n_1156),
.B2(n_1229),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1210),
.A2(n_1191),
.B(n_1241),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1268),
.B(n_1259),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1241),
.A2(n_1280),
.B(n_1245),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1271),
.B(n_1277),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1172),
.B(n_1275),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_1177),
.Y(n_1321)
);

AOI221x1_ASAP7_75t_L g1322 ( 
.A1(n_1168),
.A2(n_1271),
.B1(n_1277),
.B2(n_1165),
.C(n_1149),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1245),
.A2(n_1257),
.B(n_1280),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1217),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1188),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1196),
.A2(n_1152),
.B(n_1149),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1158),
.A2(n_1183),
.A3(n_1185),
.B(n_1257),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_1183),
.A3(n_1185),
.B(n_1274),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1181),
.A2(n_1218),
.B(n_1227),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1193),
.B(n_1215),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1195),
.B(n_1189),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1190),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1193),
.B(n_1198),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1201),
.A2(n_1237),
.B1(n_1258),
.B2(n_1267),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1194),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1211),
.B(n_1212),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1161),
.A2(n_1260),
.B(n_1224),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1202),
.A2(n_1153),
.B1(n_1204),
.B2(n_1223),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1160),
.A2(n_1208),
.B(n_1225),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1211),
.A2(n_1212),
.B(n_1226),
.C(n_1270),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1228),
.A2(n_1226),
.B(n_1220),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1242),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1164),
.B(n_1206),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1222),
.A2(n_1205),
.B(n_1150),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1274),
.A2(n_1163),
.B(n_1246),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1169),
.A2(n_1216),
.B1(n_1182),
.B2(n_1209),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1232),
.Y(n_1347)
);

NAND2xp33_ASAP7_75t_SL g1348 ( 
.A(n_1249),
.B(n_1232),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1254),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1250),
.A2(n_1276),
.B1(n_1254),
.B2(n_1281),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1254),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1163),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1281),
.B(n_1250),
.Y(n_1353)
);

AND2x2_ASAP7_75t_SL g1354 ( 
.A(n_1281),
.B(n_1276),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1247),
.A2(n_1059),
.B1(n_857),
.B2(n_735),
.C(n_1114),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1187),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1261),
.A2(n_384),
.B1(n_386),
.B2(n_351),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1262),
.B(n_843),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1147),
.A2(n_857),
.B1(n_843),
.B2(n_1089),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1207),
.A2(n_833),
.B1(n_1114),
.B2(n_1065),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1235),
.B(n_1151),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1187),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1251),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1264),
.A2(n_837),
.B1(n_1114),
.B2(n_843),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1247),
.B(n_1279),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1186),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1251),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1159),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1187),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1187),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1230),
.A2(n_1071),
.B(n_1240),
.C(n_1236),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1187),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1247),
.A2(n_894),
.B(n_843),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1187),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1172),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1159),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1175),
.A2(n_1256),
.B(n_1243),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1187),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1235),
.B(n_1151),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1159),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1182),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1159),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1172),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1159),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1247),
.B(n_894),
.C(n_857),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_L g1391 ( 
.A(n_1247),
.B(n_894),
.C(n_857),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1155),
.A2(n_1244),
.B(n_1234),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1184),
.B(n_1200),
.Y(n_1393)
);

NOR2xp67_ASAP7_75t_L g1394 ( 
.A(n_1342),
.B(n_1368),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1342),
.B(n_1330),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1329),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1353),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1296),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1329),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1283),
.B(n_1361),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1288),
.B(n_1284),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1359),
.A2(n_1360),
.B1(n_1314),
.B2(n_1358),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1382),
.B(n_1293),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1318),
.A2(n_1323),
.B(n_1316),
.Y(n_1404)
);

O2A1O1Ixp5_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1291),
.B(n_1299),
.C(n_1339),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1384),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1382),
.B(n_1301),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1340),
.A2(n_1391),
.B(n_1389),
.Y(n_1409)
);

O2A1O1Ixp5_ASAP7_75t_L g1410 ( 
.A1(n_1365),
.A2(n_1374),
.B(n_1287),
.C(n_1309),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1364),
.A2(n_1358),
.B(n_1372),
.C(n_1359),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1303),
.A2(n_1338),
.B(n_1322),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1372),
.A2(n_1319),
.B(n_1300),
.C(n_1326),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1319),
.B(n_1333),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1376),
.A2(n_1387),
.B(n_1321),
.C(n_1344),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1357),
.A2(n_1350),
.B1(n_1292),
.B2(n_1363),
.Y(n_1416)
);

OA22x2_ASAP7_75t_L g1417 ( 
.A1(n_1331),
.A2(n_1341),
.B1(n_1373),
.B2(n_1371),
.Y(n_1417)
);

OA22x2_ASAP7_75t_L g1418 ( 
.A1(n_1289),
.A2(n_1362),
.B1(n_1375),
.B2(n_1370),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1350),
.A2(n_1354),
.B1(n_1295),
.B2(n_1334),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1304),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1290),
.B(n_1356),
.Y(n_1421)
);

AND2x2_ASAP7_75t_SL g1422 ( 
.A(n_1354),
.B(n_1317),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1381),
.B(n_1336),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1345),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1311),
.Y(n_1425)
);

O2A1O1Ixp5_ASAP7_75t_L g1426 ( 
.A1(n_1366),
.A2(n_1352),
.B(n_1369),
.C(n_1379),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1311),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1304),
.Y(n_1428)
);

AOI211xp5_ASAP7_75t_L g1429 ( 
.A1(n_1355),
.A2(n_1346),
.B(n_1348),
.C(n_1320),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1297),
.A2(n_1332),
.B(n_1325),
.C(n_1313),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1298),
.A2(n_1302),
.B(n_1310),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1305),
.A2(n_1385),
.B(n_1383),
.C(n_1388),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1298),
.A2(n_1302),
.B(n_1285),
.Y(n_1433)
);

AOI31xp33_ASAP7_75t_L g1434 ( 
.A1(n_1348),
.A2(n_1393),
.A3(n_1334),
.B(n_1335),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1298),
.A2(n_1393),
.B(n_1343),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1383),
.A2(n_1385),
.B1(n_1352),
.B2(n_1324),
.C(n_1307),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1282),
.A2(n_1315),
.B1(n_1349),
.B2(n_1351),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1282),
.A2(n_1347),
.B1(n_1384),
.B2(n_1343),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1307),
.A2(n_1337),
.B1(n_1380),
.B2(n_1312),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1328),
.Y(n_1440)
);

AOI21x1_ASAP7_75t_SL g1441 ( 
.A1(n_1327),
.A2(n_1328),
.B(n_1294),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1367),
.B(n_1377),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1378),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1386),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1390),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1392),
.B(n_1317),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1283),
.B(n_1361),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1359),
.A2(n_1261),
.B1(n_1360),
.B2(n_857),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1359),
.A2(n_1261),
.B1(n_1360),
.B2(n_857),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1320),
.B(n_1283),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1342),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1303),
.A2(n_857),
.B(n_893),
.C(n_894),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1286),
.B(n_1308),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1359),
.A2(n_1261),
.B1(n_1360),
.B2(n_857),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_L g1456 ( 
.A(n_1354),
.Y(n_1456)
);

CKINVDCx6p67_ASAP7_75t_R g1457 ( 
.A(n_1384),
.Y(n_1457)
);

O2A1O1Ixp5_ASAP7_75t_L g1458 ( 
.A1(n_1365),
.A2(n_1291),
.B(n_1299),
.C(n_1175),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1296),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1432),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1424),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1442),
.B(n_1440),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1402),
.A2(n_1455),
.B1(n_1450),
.B2(n_1449),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1431),
.B(n_1433),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1404),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1414),
.B(n_1423),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1445),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1447),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1426),
.A2(n_1405),
.B(n_1439),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1446),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1447),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1421),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1435),
.B(n_1401),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1396),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1415),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1418),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1418),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1430),
.Y(n_1480)
);

INVx4_ASAP7_75t_SL g1481 ( 
.A(n_1401),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1401),
.B(n_1409),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1430),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1444),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1405),
.A2(n_1410),
.B(n_1458),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1417),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1417),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1443),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1443),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1415),
.A2(n_1411),
.B(n_1437),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1397),
.Y(n_1492)
);

OAI21xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1434),
.A2(n_1422),
.B(n_1413),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1458),
.B(n_1453),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1400),
.B(n_1448),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1468),
.B(n_1474),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1467),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1475),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1479),
.B(n_1425),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1451),
.Y(n_1501)
);

INVx5_ASAP7_75t_L g1502 ( 
.A(n_1464),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1480),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1468),
.B(n_1403),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1474),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1492),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1476),
.B(n_1413),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1470),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_1408),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1479),
.A2(n_1419),
.B1(n_1456),
.B2(n_1416),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1470),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1465),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1465),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1438),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1474),
.B(n_1488),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1463),
.A2(n_1456),
.B1(n_1395),
.B2(n_1407),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1499),
.B(n_1493),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1496),
.B(n_1515),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1498),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1508),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1509),
.Y(n_1523)
);

NAND4xp25_ASAP7_75t_L g1524 ( 
.A(n_1507),
.B(n_1463),
.C(n_1429),
.D(n_1480),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1510),
.A2(n_1482),
.B1(n_1486),
.B2(n_1487),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1498),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1508),
.Y(n_1527)
);

OAI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1510),
.A2(n_1490),
.B(n_1493),
.C(n_1486),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1511),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1507),
.A2(n_1482),
.B1(n_1490),
.B2(n_1491),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1503),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1517),
.A2(n_1482),
.B1(n_1487),
.B2(n_1473),
.C(n_1466),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1514),
.A2(n_1482),
.B1(n_1491),
.B2(n_1494),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1514),
.A2(n_1482),
.B(n_1494),
.Y(n_1534)
);

AOI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1503),
.A2(n_1477),
.B1(n_1478),
.B2(n_1483),
.C(n_1472),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1497),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1514),
.A2(n_1482),
.B1(n_1491),
.B2(n_1494),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1517),
.A2(n_1473),
.B1(n_1484),
.B2(n_1494),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1499),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1506),
.Y(n_1541)
);

OAI211xp5_ASAP7_75t_L g1542 ( 
.A1(n_1516),
.A2(n_1494),
.B(n_1485),
.C(n_1483),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1496),
.B(n_1471),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1514),
.A2(n_1491),
.B1(n_1485),
.B2(n_1473),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1485),
.C(n_1477),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1502),
.B(n_1489),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1514),
.A2(n_1485),
.B1(n_1473),
.B2(n_1464),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1500),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1502),
.B(n_1489),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1514),
.A2(n_1473),
.B1(n_1484),
.B2(n_1478),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1502),
.A2(n_1485),
.B1(n_1464),
.B2(n_1469),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1502),
.B(n_1489),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1522),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1521),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1550),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1522),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1527),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1526),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1519),
.Y(n_1561)
);

NOR2xp67_ASAP7_75t_L g1562 ( 
.A(n_1545),
.B(n_1502),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1546),
.B(n_1502),
.Y(n_1564)
);

AOI21xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1540),
.A2(n_1427),
.B(n_1459),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1539),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1546),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1528),
.B(n_1502),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1518),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1524),
.B(n_1469),
.C(n_1460),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1523),
.B(n_1515),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1530),
.B(n_1481),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1505),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1559),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1561),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1555),
.B(n_1543),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1561),
.Y(n_1581)
);

OAI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1571),
.A2(n_1524),
.B(n_1544),
.C(n_1542),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1572),
.B(n_1501),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1555),
.B(n_1547),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1555),
.B(n_1549),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1572),
.B(n_1535),
.Y(n_1586)
);

O2A1O1Ixp5_ASAP7_75t_L g1587 ( 
.A1(n_1571),
.A2(n_1525),
.B(n_1534),
.C(n_1538),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1559),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1567),
.B(n_1536),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1556),
.B(n_1501),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1556),
.B(n_1501),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1573),
.B(n_1505),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1570),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1563),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1554),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1573),
.B(n_1504),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1574),
.B(n_1504),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1577),
.B(n_1541),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1554),
.Y(n_1605)
);

OAI31xp33_ASAP7_75t_L g1606 ( 
.A1(n_1575),
.A2(n_1532),
.A3(n_1533),
.B(n_1537),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1560),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1558),
.B(n_1566),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1558),
.B(n_1548),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1610)
);

AND4x1_ASAP7_75t_L g1611 ( 
.A(n_1577),
.B(n_1544),
.C(n_1545),
.D(n_1551),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1569),
.B(n_1553),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1577),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1558),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1588),
.B(n_1560),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.B(n_1560),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1598),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1584),
.B(n_1570),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1611),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1570),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1598),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1602),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

AOI21xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1604),
.A2(n_1575),
.B(n_1398),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1605),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1583),
.B(n_1566),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1613),
.B(n_1577),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1607),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1579),
.B(n_1566),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1581),
.B(n_1577),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1586),
.B(n_1577),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1576),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1605),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1582),
.B(n_1576),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1614),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1614),
.Y(n_1637)
);

AOI211x1_ASAP7_75t_SL g1638 ( 
.A1(n_1599),
.A2(n_1562),
.B(n_1394),
.C(n_1557),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1578),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1611),
.B(n_1587),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1595),
.B(n_1562),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1608),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1606),
.B(n_1564),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1591),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1593),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1578),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1596),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1601),
.B(n_1495),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1629),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1619),
.A2(n_1606),
.B1(n_1595),
.B2(n_1552),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1639),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1646),
.B(n_1633),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1641),
.B(n_1585),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1641),
.B(n_1600),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1629),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1640),
.A2(n_1592),
.B(n_1589),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1641),
.B(n_1600),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1648),
.B(n_1603),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1615),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1640),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1648),
.B(n_1603),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1565),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1622),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1622),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1592),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1615),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1644),
.A2(n_1464),
.B1(n_1597),
.B2(n_1457),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1565),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1630),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1654),
.A2(n_1644),
.B(n_1635),
.Y(n_1677)
);

OAI32xp33_ASAP7_75t_L g1678 ( 
.A1(n_1654),
.A2(n_1638),
.A3(n_1631),
.B1(n_1630),
.B2(n_1620),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1653),
.B(n_1618),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1653),
.B(n_1620),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1665),
.A2(n_1623),
.B(n_1649),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1650),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1665),
.B(n_1649),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1659),
.B(n_1642),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1652),
.A2(n_1625),
.B(n_1643),
.C(n_1597),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1660),
.A2(n_1626),
.B1(n_1637),
.B2(n_1624),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1652),
.A2(n_1452),
.B1(n_1428),
.B2(n_1420),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1674),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1660),
.A2(n_1623),
.B1(n_1617),
.B2(n_1621),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1634),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1673),
.B(n_1564),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1674),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1676),
.Y(n_1693)
);

AND3x2_ASAP7_75t_L g1694 ( 
.A(n_1651),
.B(n_1636),
.C(n_1645),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1676),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1652),
.A2(n_1627),
.B(n_1590),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1688),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1694),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1679),
.B(n_1653),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1692),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1677),
.B(n_1651),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1667),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1693),
.B(n_1651),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1695),
.Y(n_1706)
);

AND2x4_ASAP7_75t_SL g1707 ( 
.A(n_1686),
.B(n_1672),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1681),
.B(n_1672),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1702),
.A2(n_1689),
.B1(n_1686),
.B2(n_1673),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1707),
.A2(n_1678),
.B1(n_1689),
.B2(n_1696),
.C(n_1655),
.Y(n_1711)
);

AOI22x1_ASAP7_75t_L g1712 ( 
.A1(n_1699),
.A2(n_1672),
.B1(n_1656),
.B2(n_1664),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1707),
.A2(n_1685),
.B(n_1675),
.C(n_1691),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1703),
.B(n_1684),
.C(n_1690),
.D(n_1655),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1700),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1698),
.B(n_1657),
.Y(n_1716)
);

OAI321xp33_ASAP7_75t_L g1717 ( 
.A1(n_1708),
.A2(n_1658),
.A3(n_1661),
.B1(n_1657),
.B2(n_1687),
.C(n_1663),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1705),
.A2(n_1661),
.B(n_1658),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1699),
.A2(n_1658),
.B(n_1661),
.C(n_1670),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1716),
.Y(n_1720)
);

AOI31xp33_ASAP7_75t_L g1721 ( 
.A1(n_1711),
.A2(n_1709),
.A3(n_1704),
.B(n_1697),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1715),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1710),
.A2(n_1709),
.B(n_1706),
.C(n_1701),
.Y(n_1723)
);

AOI211x1_ASAP7_75t_SL g1724 ( 
.A1(n_1713),
.A2(n_1670),
.B(n_1660),
.C(n_1645),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1722),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1720),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1721),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1723),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1724),
.B(n_1714),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_L g1730 ( 
.A(n_1720),
.B(n_1664),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1726),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1730),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1727),
.B(n_1712),
.C(n_1719),
.Y(n_1733)
);

AOI222xp33_ASAP7_75t_L g1734 ( 
.A1(n_1728),
.A2(n_1717),
.B1(n_1700),
.B2(n_1718),
.C1(n_1664),
.C2(n_1660),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1725),
.B(n_1664),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1735),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1731),
.B(n_1662),
.Y(n_1737)
);

NAND4xp25_ASAP7_75t_L g1738 ( 
.A(n_1733),
.B(n_1729),
.C(n_1664),
.D(n_1663),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1737),
.A2(n_1734),
.B(n_1738),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1739),
.Y(n_1740)
);

OR5x1_ASAP7_75t_L g1741 ( 
.A(n_1740),
.B(n_1736),
.C(n_1732),
.D(n_1669),
.E(n_1668),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1740),
.A2(n_1663),
.B1(n_1669),
.B2(n_1668),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1671),
.B1(n_1666),
.B2(n_1662),
.Y(n_1743)
);

OAI22x1_ASAP7_75t_L g1744 ( 
.A1(n_1741),
.A2(n_1671),
.B1(n_1666),
.B2(n_1662),
.Y(n_1744)
);

AOI22x1_ASAP7_75t_L g1745 ( 
.A1(n_1744),
.A2(n_1671),
.B1(n_1666),
.B2(n_1406),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1745),
.Y(n_1746)
);

AO22x2_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1743),
.B1(n_1591),
.B2(n_1627),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1747),
.B(n_1591),
.Y(n_1748)
);

OAI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1590),
.B1(n_1594),
.B2(n_1593),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1612),
.B1(n_1610),
.B2(n_1570),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1612),
.B(n_1594),
.C(n_1609),
.Y(n_1751)
);


endmodule