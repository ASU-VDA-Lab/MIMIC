module fake_jpeg_19429_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_12),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_29),
.B1(n_28),
.B2(n_14),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_56),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_16),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_28),
.B1(n_14),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_20),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_17),
.B1(n_25),
.B2(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_68),
.Y(n_135)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_75),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_43),
.B1(n_42),
.B2(n_33),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_74),
.A2(n_90),
.B1(n_97),
.B2(n_106),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_83),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_37),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_85),
.B(n_86),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_82),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_79),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_30),
.B1(n_22),
.B2(n_17),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_53),
.CI(n_51),
.CON(n_81),
.SN(n_81)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_87),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_43),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_30),
.B1(n_22),
.B2(n_17),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_100),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_18),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_93),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_18),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_46),
.B1(n_45),
.B2(n_19),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_110),
.B1(n_1),
.B2(n_3),
.Y(n_130)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_19),
.C(n_20),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_104),
.Y(n_116)
);

INVx11_ASAP7_75t_SL g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_103),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_15),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_66),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_15),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_105),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_66),
.B1(n_49),
.B2(n_20),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_12),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_108),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_49),
.A2(n_20),
.B1(n_12),
.B2(n_15),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_130),
.B1(n_137),
.B2(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_141),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_94),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_5),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_69),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_134),
.B(n_128),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_85),
.C(n_77),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_111),
.C(n_116),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_160),
.B(n_115),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_73),
.B1(n_67),
.B2(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_159),
.Y(n_182)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_125),
.B1(n_127),
.B2(n_135),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_69),
.B1(n_90),
.B2(n_92),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_171),
.B1(n_135),
.B2(n_91),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_114),
.A2(n_101),
.B1(n_104),
.B2(n_100),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_95),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_77),
.B(n_87),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_121),
.B(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_93),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_93),
.Y(n_166)
);

OR2x2_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_102),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_131),
.C(n_126),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_79),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_169),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_76),
.B1(n_107),
.B2(n_68),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_111),
.B1(n_122),
.B2(n_102),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_95),
.B1(n_83),
.B2(n_70),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_177),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_84),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_84),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_180),
.C(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_116),
.C(n_174),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_183),
.A2(n_188),
.B1(n_165),
.B2(n_154),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_140),
.B1(n_138),
.B2(n_118),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_199),
.B(n_204),
.Y(n_219)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_126),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_163),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_166),
.B(n_173),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_202),
.Y(n_210)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_117),
.B(n_134),
.C(n_130),
.D(n_137),
.Y(n_196)
);

OA21x2_ASAP7_75t_SL g231 ( 
.A1(n_196),
.A2(n_149),
.B(n_152),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_205),
.B1(n_159),
.B2(n_153),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_115),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_127),
.B(n_129),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_129),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_135),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_96),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_160),
.B(n_157),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_207),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_232),
.B(n_192),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_221),
.B1(n_233),
.B2(n_235),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_217),
.C(n_183),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_218),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_174),
.C(n_150),
.Y(n_217)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_184),
.A3(n_186),
.B1(n_203),
.B2(n_202),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_160),
.B1(n_152),
.B2(n_155),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_203),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_161),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_229),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_198),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_201),
.B(n_185),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_172),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_171),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_154),
.B1(n_125),
.B2(n_132),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_244),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_253),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_210),
.B(n_193),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_186),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_209),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_219),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_191),
.B1(n_196),
.B2(n_204),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_221),
.B1(n_224),
.B2(n_218),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_209),
.B1(n_200),
.B2(n_187),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_235),
.B1(n_233),
.B2(n_228),
.Y(n_260)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_211),
.B(n_208),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_232),
.B(n_219),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_261),
.B(n_266),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_258),
.A2(n_250),
.B1(n_254),
.B2(n_195),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_272),
.B1(n_239),
.B2(n_249),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_200),
.B(n_227),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_264),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_271),
.C(n_273),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_227),
.B1(n_210),
.B2(n_187),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_193),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_223),
.B1(n_222),
.B2(n_125),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_223),
.C(n_222),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_268),
.Y(n_275)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_279),
.B1(n_284),
.B2(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_239),
.B1(n_252),
.B2(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_273),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_195),
.B(n_189),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_132),
.B(n_262),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_189),
.B1(n_132),
.B2(n_9),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_132),
.C(n_72),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_264),
.C(n_263),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_269),
.B(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_286),
.Y(n_298)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_275),
.C(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_282),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_296),
.C(n_277),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_265),
.C(n_256),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_285),
.C(n_281),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_303),
.C(n_291),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_289),
.A3(n_292),
.B1(n_294),
.B2(n_10),
.C1(n_7),
.C2(n_9),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_287),
.B(n_290),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_300),
.B(n_304),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

OAI21x1_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_307),
.B(n_8),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_310),
.C(n_8),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_7),
.C(n_9),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_314),
.C(n_11),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_11),
.Y(n_318)
);


endmodule