module fake_jpeg_13892_n_442 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_53),
.B(n_62),
.Y(n_136)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_15),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_65),
.B(n_78),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_15),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_15),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_88),
.Y(n_98)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_0),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_27),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_22),
.B1(n_41),
.B2(n_40),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_42),
.B1(n_87),
.B2(n_86),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_22),
.B1(n_41),
.B2(n_21),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_96),
.B1(n_110),
.B2(n_115),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_30),
.B1(n_40),
.B2(n_22),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_84),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_137),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_123)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_61),
.B1(n_57),
.B2(n_56),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_24),
.B1(n_34),
.B2(n_37),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_43),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_163),
.B1(n_175),
.B2(n_95),
.Y(n_188)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_59),
.A3(n_85),
.B1(n_50),
.B2(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_152),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_153),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_165),
.B(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_33),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_155),
.B(n_156),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_33),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_90),
.Y(n_157)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_35),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_66),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_162),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_42),
.B1(n_70),
.B2(n_68),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_120),
.B1(n_114),
.B2(n_113),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_98),
.B(n_37),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_122),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_94),
.B(n_36),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_110),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_36),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_205)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_35),
.C(n_29),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_52),
.B1(n_48),
.B2(n_29),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_89),
.C(n_2),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.Y(n_186)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_133),
.B1(n_111),
.B2(n_119),
.Y(n_208)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_181),
.Y(n_202)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

NAND2x1_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_129),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_3),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_184),
.Y(n_207)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_189),
.B1(n_200),
.B2(n_179),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_96),
.B1(n_115),
.B2(n_135),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_111),
.B1(n_119),
.B2(n_112),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_91),
.B(n_117),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_154),
.B(n_117),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_158),
.B1(n_143),
.B2(n_99),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_145),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_219),
.B1(n_164),
.B2(n_157),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_131),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_144),
.A2(n_120),
.B1(n_114),
.B2(n_113),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_242),
.B1(n_244),
.B2(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_225),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_164),
.B1(n_180),
.B2(n_167),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_229),
.C(n_237),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_141),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_182),
.B(n_170),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_236),
.B(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_151),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_235),
.B(n_239),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_164),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_148),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_146),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_142),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_188),
.B1(n_198),
.B2(n_217),
.Y(n_252)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_246),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_184),
.B1(n_181),
.B2(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_166),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_187),
.Y(n_275)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_216),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_276),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_223),
.B1(n_233),
.B2(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_258),
.B(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_192),
.B1(n_212),
.B2(n_201),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_229),
.B(n_208),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_260),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_221),
.B(n_201),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_196),
.B(n_201),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_267),
.B(n_236),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_199),
.B(n_195),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_238),
.B(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_196),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_266),
.B(n_234),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_199),
.B(n_185),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_217),
.B1(n_190),
.B2(n_185),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_225),
.B1(n_254),
.B2(n_244),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_246),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_285),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_275),
.Y(n_282)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_283),
.A2(n_277),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_243),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_291),
.B1(n_298),
.B2(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_249),
.B(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_289),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_270),
.B(n_228),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_260),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_222),
.C(n_230),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_303),
.C(n_283),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_304),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_258),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_222),
.B1(n_239),
.B2(n_220),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_299),
.B1(n_302),
.B2(n_274),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_257),
.A2(n_253),
.B1(n_264),
.B2(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_241),
.B1(n_190),
.B2(n_226),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_300),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_265),
.B(n_227),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_187),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_256),
.A2(n_195),
.B(n_197),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_309),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_259),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_310),
.B(n_285),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_297),
.B1(n_284),
.B2(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_309),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_261),
.B1(n_250),
.B2(n_267),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_315),
.A2(n_325),
.B1(n_328),
.B2(n_299),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_261),
.B(n_262),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_277),
.B1(n_280),
.B2(n_300),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_261),
.C(n_263),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_321),
.C(n_327),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_273),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_323),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_269),
.C(n_161),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_269),
.B1(n_255),
.B2(n_268),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_271),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_298),
.A2(n_255),
.B1(n_268),
.B2(n_271),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_197),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_268),
.B1(n_190),
.B2(n_211),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_333),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_289),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_315),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_282),
.B1(n_292),
.B2(n_302),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_279),
.B1(n_303),
.B2(n_288),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_345),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_340),
.A2(n_343),
.B1(n_308),
.B2(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_311),
.A2(n_293),
.B1(n_295),
.B2(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_211),
.C(n_89),
.Y(n_346)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_91),
.B(n_193),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_149),
.B(n_131),
.Y(n_372)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_351),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_206),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_321),
.C(n_327),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_206),
.Y(n_353)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_355),
.A2(n_334),
.B1(n_336),
.B2(n_342),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_325),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_305),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_362),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_323),
.C(n_310),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_366),
.C(n_370),
.Y(n_374)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_340),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_319),
.C(n_313),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_173),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_313),
.C(n_318),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_328),
.C(n_160),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_371),
.B(n_350),
.C(n_348),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_149),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_386),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_345),
.C(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_379),
.A2(n_384),
.B1(n_360),
.B2(n_361),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_368),
.B(n_332),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_7),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_343),
.C(n_339),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_363),
.C(n_368),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_389),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_3),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_365),
.A2(n_4),
.B(n_5),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_388),
.B(n_390),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_358),
.A2(n_4),
.B(n_5),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_355),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_5),
.B(n_7),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_398),
.Y(n_417)
);

FAx1_ASAP7_75t_SL g392 ( 
.A(n_383),
.B(n_357),
.CI(n_369),
.CON(n_392),
.SN(n_392)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_397),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_403),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_359),
.B1(n_364),
.B2(n_367),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_385),
.A2(n_373),
.B1(n_354),
.B2(n_372),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_371),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_15),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_399),
.A2(n_379),
.B(n_11),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g400 ( 
.A(n_374),
.B(n_7),
.CI(n_9),
.CON(n_400),
.SN(n_400)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_386),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_10),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_374),
.C(n_404),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_407),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_391),
.A2(n_376),
.B(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_408),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_401),
.C(n_396),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_416),
.Y(n_419)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_412),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_380),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_405),
.A2(n_10),
.B(n_11),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_392),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_422),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_400),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_411),
.A2(n_402),
.B(n_393),
.C(n_394),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_413),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_403),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_418),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_410),
.C(n_414),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_427),
.A2(n_428),
.B(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_409),
.C(n_413),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_430),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_431),
.A2(n_432),
.B(n_419),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_433),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_434),
.A2(n_436),
.B(n_412),
.C(n_399),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_426),
.C(n_424),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_435),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_439),
.A2(n_437),
.B(n_12),
.C(n_13),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_440),
.A2(n_11),
.B(n_12),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_13),
.Y(n_442)
);


endmodule