module fake_jpeg_3859_n_157 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_157);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_13),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_35),
.B1(n_16),
.B2(n_12),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_42),
.B1(n_30),
.B2(n_36),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_16),
.B(n_19),
.C(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_60),
.Y(n_67)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_31),
.B1(n_30),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_40),
.B1(n_30),
.B2(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_62),
.B1(n_40),
.B2(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_45),
.B(n_43),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_72),
.B1(n_39),
.B2(n_24),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_44),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_26),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_51),
.A3(n_60),
.B1(n_54),
.B2(n_50),
.C1(n_56),
.C2(n_53),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_59),
.B1(n_49),
.B2(n_40),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_27),
.C(n_38),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_67),
.C(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_37),
.B1(n_44),
.B2(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_62),
.B1(n_70),
.B2(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_66),
.B1(n_65),
.B2(n_32),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_83),
.C(n_77),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_27),
.B(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_73),
.B1(n_86),
.B2(n_87),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_66),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_113),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_25),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_39),
.B1(n_26),
.B2(n_29),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_14),
.B1(n_18),
.B2(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_18),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_92),
.C(n_100),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_89),
.A3(n_96),
.B1(n_95),
.B2(n_91),
.C1(n_98),
.C2(n_27),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_121),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_25),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_114),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_107),
.Y(n_126)
);

OAI21x1_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_25),
.B(n_4),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_3),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_109),
.C(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.C(n_132),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_104),
.C(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_25),
.C(n_14),
.Y(n_132)
);

AOI31xp67_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_14),
.A3(n_1),
.B(n_2),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_3),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_116),
.B1(n_123),
.B2(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_141),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_4),
.B(n_5),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_144),
.B(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_145),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_131),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_138),
.B(n_140),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_138),
.B(n_6),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_6),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_7),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.C(n_7),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_147),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_9),
.Y(n_157)
);


endmodule