module fake_jpeg_11092_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_5),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_1),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_2),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_68),
.B(n_59),
.C(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_4),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_68),
.B(n_59),
.C(n_65),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_89),
.B(n_61),
.C(n_6),
.D(n_7),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_62),
.C(n_67),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_93),
.B(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_70),
.B1(n_72),
.B2(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_61),
.B1(n_10),
.B2(n_12),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_52),
.B1(n_70),
.B2(n_63),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_56),
.Y(n_101)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_13),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_51),
.B1(n_74),
.B2(n_60),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_103),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_74),
.B1(n_52),
.B2(n_71),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_111),
.B(n_99),
.C(n_100),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_119),
.B(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_5),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_8),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_15),
.C(n_21),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_9),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_13),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_117),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_14),
.B(n_61),
.C(n_17),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_38),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_138),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_91),
.B(n_87),
.C(n_19),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_35),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_14),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_23),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_110),
.C(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_46),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_50),
.B(n_25),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_24),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_149),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_153),
.B1(n_121),
.B2(n_127),
.C(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_118),
.B(n_30),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_155),
.B(n_156),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_122),
.C(n_128),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_47),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_49),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_160),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_164),
.Y(n_171)
);

AOI332xp33_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_166),
.A3(n_167),
.B1(n_159),
.B2(n_134),
.B3(n_153),
.C1(n_151),
.C2(n_161),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_152),
.C(n_155),
.Y(n_173)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_123),
.A3(n_145),
.B1(n_147),
.B2(n_161),
.C(n_170),
.Y(n_174)
);


endmodule