module fake_aes_2791_n_669 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_669);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_669;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_48), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_2), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_49), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_25), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_75), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_34), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_55), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_1), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_46), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_19), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_54), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_29), .Y(n_92) );
XNOR2xp5_ASAP7_75t_SL g93 ( .A(n_62), .B(n_18), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_20), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_56), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_22), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_10), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_50), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_3), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_28), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_16), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_42), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_58), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_44), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_5), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_60), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_67), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_20), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_21), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_74), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_79), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_94), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_89), .B(n_99), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_110), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_113), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_102), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVxp33_ASAP7_75t_SL g142 ( .A(n_99), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_86), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_78), .B(n_0), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_93), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_84), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_82), .Y(n_151) );
CKINVDCx6p67_ASAP7_75t_R g152 ( .A(n_91), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_123), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_98), .Y(n_155) );
OR2x2_ASAP7_75t_L g156 ( .A(n_85), .B(n_3), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_91), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_77), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_116), .B(n_4), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_88), .B(n_4), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_109), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_88), .B(n_5), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_97), .B(n_6), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_87), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
AO22x2_ASAP7_75t_L g169 ( .A1(n_159), .A2(n_124), .B1(n_95), .B2(n_120), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_149), .B(n_121), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_149), .B(n_115), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_159), .B(n_124), .Y(n_173) );
NAND2xp33_ASAP7_75t_L g174 ( .A(n_143), .B(n_95), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_159), .B(n_122), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_157), .B(n_106), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_125), .B(n_96), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
NOR3xp33_ASAP7_75t_L g182 ( .A(n_145), .B(n_111), .C(n_117), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx8_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_156), .A2(n_96), .B1(n_120), .B2(n_119), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_133), .A2(n_122), .B1(n_104), .B2(n_118), .C(n_105), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g190 ( .A(n_134), .B(n_105), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_142), .B(n_101), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_132), .B(n_107), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_131), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_132), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_125), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_126), .B(n_119), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_126), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_127), .B(n_108), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_150), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_133), .B(n_118), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_131), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_154), .B(n_127), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_136), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_128), .B(n_114), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_154), .B(n_104), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_128), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_136), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_129), .B(n_114), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_129), .B(n_103), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_135), .B(n_107), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_139), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_208), .B(n_156), .Y(n_228) );
CKINVDCx6p67_ASAP7_75t_R g229 ( .A(n_185), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_214), .A2(n_146), .B1(n_145), .B2(n_153), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_202), .B(n_146), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_211), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_206), .Y(n_233) );
NOR3xp33_ASAP7_75t_L g234 ( .A(n_189), .B(n_163), .C(n_160), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_214), .B(n_165), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_214), .B(n_165), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_214), .B(n_135), .Y(n_237) );
INVxp67_ASAP7_75t_L g238 ( .A(n_194), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_211), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_212), .B(n_163), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_202), .B(n_137), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_212), .B(n_218), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_180), .B(n_103), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_178), .B(n_164), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_191), .B(n_160), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_211), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_166), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_211), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_184), .B(n_144), .Y(n_252) );
NOR2xp67_ASAP7_75t_L g253 ( .A(n_210), .B(n_150), .Y(n_253) );
OR2x6_ASAP7_75t_L g254 ( .A(n_185), .B(n_144), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_212), .B(n_150), .Y(n_256) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_190), .B(n_112), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_212), .B(n_100), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_166), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_218), .B(n_90), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_180), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_170), .B(n_83), .C(n_130), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_180), .B(n_141), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_166), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_218), .B(n_6), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_205), .B(n_141), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_185), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_218), .B(n_141), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g273 ( .A(n_182), .B(n_140), .C(n_139), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_192), .B(n_140), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_192), .B(n_140), .Y(n_275) );
AO22x1_ASAP7_75t_L g276 ( .A1(n_208), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_185), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_216), .A2(n_8), .B(n_9), .C(n_10), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
AND3x1_ASAP7_75t_SL g280 ( .A(n_186), .B(n_11), .C(n_12), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_205), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_221), .B(n_36), .Y(n_283) );
BUFx8_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_203), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_210), .Y(n_286) );
AND2x6_ASAP7_75t_L g287 ( .A(n_203), .B(n_38), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
NOR3xp33_ASAP7_75t_SL g289 ( .A(n_172), .B(n_11), .C(n_12), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_186), .Y(n_290) );
NOR3xp33_ASAP7_75t_SL g291 ( .A(n_209), .B(n_13), .C(n_14), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_242), .B(n_224), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_252), .B(n_186), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_240), .B(n_186), .Y(n_295) );
INVx3_ASAP7_75t_SL g296 ( .A(n_229), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_240), .B(n_219), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_243), .B(n_219), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_237), .B(n_207), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_267), .B(n_208), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_247), .A2(n_221), .B(n_173), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_250), .B(n_224), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_249), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_247), .A2(n_204), .B(n_207), .C(n_175), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_267), .B(n_203), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_254), .B(n_175), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_290), .A2(n_169), .B1(n_166), .B2(n_175), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_279), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_256), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_169), .B1(n_174), .B2(n_173), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_275), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_237), .B(n_204), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_228), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_245), .A2(n_173), .B(n_169), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_244), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_284), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_234), .A2(n_223), .B(n_177), .C(n_198), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_233), .B(n_169), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_262), .B(n_175), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_235), .B(n_168), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_281), .A2(n_179), .B1(n_171), .B2(n_197), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_244), .B(n_196), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_228), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_246), .A2(n_179), .B(n_171), .C(n_197), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_277), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_269), .B(n_177), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_234), .A2(n_198), .B(n_188), .C(n_201), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_236), .B(n_188), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_254), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_236), .B(n_201), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_254), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_272), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_241), .Y(n_336) );
CKINVDCx14_ASAP7_75t_R g337 ( .A(n_260), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_244), .Y(n_339) );
NOR2xp33_ASAP7_75t_R g340 ( .A(n_285), .B(n_196), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_300), .A2(n_263), .B1(n_270), .B2(n_282), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_300), .A2(n_227), .B1(n_258), .B2(n_245), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_309), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_323), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_323), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_294), .B(n_246), .Y(n_346) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_316), .A2(n_283), .B(n_278), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_325), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_297), .B(n_261), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_295), .B(n_227), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_336), .A2(n_261), .B1(n_264), .B2(n_257), .C(n_230), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_315), .B(n_244), .Y(n_353) );
OAI222xp33_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_280), .B1(n_276), .B2(n_283), .C1(n_231), .C2(n_291), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_331), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_273), .B1(n_264), .B2(n_289), .C(n_291), .Y(n_357) );
INVx4_ASAP7_75t_SL g358 ( .A(n_300), .Y(n_358) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_316), .A2(n_268), .B(n_265), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_312), .A2(n_287), .B1(n_288), .B2(n_271), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_320), .A2(n_268), .B(n_265), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_313), .A2(n_287), .B1(n_271), .B2(n_266), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_306), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_297), .B(n_249), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_302), .B(n_259), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_302), .B(n_259), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_292), .B(n_279), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_306), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_346), .A2(n_352), .B1(n_350), .B2(n_345), .C(n_344), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_346), .A2(n_330), .B1(n_299), .B2(n_314), .C(n_303), .Y(n_373) );
INVx4_ASAP7_75t_L g374 ( .A(n_358), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_345), .B(n_326), .Y(n_375) );
AND2x4_ASAP7_75t_SL g376 ( .A(n_364), .B(n_307), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_370), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_352), .A2(n_330), .B1(n_299), .B2(n_314), .C(n_305), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_357), .A2(n_307), .B1(n_321), .B2(n_293), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_361), .A2(n_327), .B(n_193), .Y(n_380) );
OA21x2_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_167), .B(n_193), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_308), .B1(n_324), .B2(n_310), .C(n_298), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_370), .B(n_332), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_181), .B(n_167), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_364), .A2(n_334), .B1(n_328), .B2(n_280), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_350), .B(n_301), .C(n_253), .D(n_298), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_343), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_343), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_370), .B(n_329), .Y(n_389) );
AO22x1_ASAP7_75t_L g390 ( .A1(n_364), .A2(n_296), .B1(n_287), .B2(n_318), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_367), .A2(n_329), .B1(n_322), .B2(n_335), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_343), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_351), .B(n_329), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_333), .B(n_287), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_289), .B(n_340), .C(n_317), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_347), .A2(n_342), .B(n_359), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_375), .B(n_362), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_375), .B(n_351), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_385), .A2(n_363), .B(n_360), .Y(n_400) );
OAI33xp33_ASAP7_75t_L g401 ( .A1(n_386), .A2(n_342), .A3(n_341), .B1(n_356), .B2(n_366), .B3(n_349), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_391), .B1(n_372), .B2(n_393), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_374), .Y(n_403) );
INVx8_ASAP7_75t_L g404 ( .A(n_371), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
INVx6_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_372), .A2(n_341), .B1(n_364), .B2(n_363), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_371), .B(n_351), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_393), .B(n_367), .Y(n_409) );
OAI222xp33_ASAP7_75t_L g410 ( .A1(n_379), .A2(n_362), .B1(n_360), .B2(n_368), .C1(n_322), .C2(n_348), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_386), .A2(n_322), .B1(n_365), .B2(n_366), .C(n_349), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_396), .A2(n_347), .B(n_354), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_396), .A2(n_368), .B(n_369), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_387), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_395), .A2(n_347), .B(n_368), .Y(n_415) );
OR2x6_ASAP7_75t_L g416 ( .A(n_374), .B(n_355), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_373), .A2(n_356), .B1(n_358), .B2(n_347), .Y(n_417) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_395), .B(n_337), .C(n_348), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_382), .A2(n_353), .A3(n_355), .B(n_365), .Y(n_419) );
INVx5_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_389), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_383), .B(n_355), .Y(n_423) );
AO21x1_ASAP7_75t_SL g424 ( .A1(n_394), .A2(n_358), .B(n_287), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_373), .A2(n_348), .B1(n_304), .B2(n_317), .C(n_255), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_376), .B(n_358), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_358), .B1(n_353), .B2(n_348), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_376), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_378), .A2(n_358), .B1(n_353), .B2(n_359), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_389), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_394), .A2(n_359), .B(n_369), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_387), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_423), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_403), .Y(n_436) );
OAI31xp33_ASAP7_75t_L g437 ( .A1(n_402), .A2(n_376), .A3(n_353), .B(n_390), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_409), .B(n_392), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_409), .B(n_392), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_408), .B(n_392), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_414), .Y(n_441) );
INVx5_ASAP7_75t_SL g442 ( .A(n_427), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_408), .B(n_388), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_433), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
OAI33xp33_ASAP7_75t_L g446 ( .A1(n_405), .A2(n_181), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_15), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_415), .A2(n_388), .B(n_387), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_403), .B(n_378), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_421), .B(n_380), .Y(n_451) );
AO31x2_ASAP7_75t_L g452 ( .A1(n_407), .A2(n_388), .A3(n_369), .B(n_380), .Y(n_452) );
OAI31xp33_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_390), .A3(n_339), .B(n_286), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_417), .B(n_384), .C(n_380), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_399), .B(n_384), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_432), .Y(n_457) );
AOI31xp33_ASAP7_75t_L g458 ( .A1(n_427), .A2(n_384), .A3(n_15), .B(n_24), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_417), .B(n_384), .C(n_380), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_431), .B(n_359), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_432), .B(n_338), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_430), .B(n_381), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_430), .B(n_381), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_422), .B(n_381), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_411), .B(n_225), .C(n_213), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_420), .B(n_338), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_420), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_398), .B(n_404), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
OAI31xp33_ASAP7_75t_L g474 ( .A1(n_419), .A2(n_266), .A3(n_248), .B(n_239), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_400), .A2(n_381), .B(n_338), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_404), .B(n_381), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_406), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_404), .B(n_23), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_406), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_428), .B(n_319), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_428), .B(n_187), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_401), .A2(n_319), .B1(n_309), .B2(n_176), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_404), .B(n_319), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_427), .B(n_187), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_444), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_438), .B(n_424), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_473), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_454), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g490 ( .A(n_454), .B(n_429), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_438), .B(n_416), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_437), .B(n_418), .C(n_426), .D(n_176), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
OR2x4_ASAP7_75t_L g494 ( .A(n_458), .B(n_406), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_436), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_473), .Y(n_496) );
NOR2xp33_ASAP7_75t_R g497 ( .A(n_454), .B(n_416), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_440), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_416), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_443), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_439), .B(n_416), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_435), .B(n_183), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_443), .B(n_183), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_464), .B(n_187), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_448), .B(n_485), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_464), .B(n_187), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_466), .B(n_187), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_441), .B(n_183), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_454), .B(n_183), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_468), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_441), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_468), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_466), .B(n_183), .Y(n_515) );
OAI31xp33_ASAP7_75t_L g516 ( .A1(n_437), .A2(n_220), .A3(n_200), .B(n_226), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_467), .B(n_26), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_445), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_460), .B(n_226), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_471), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_467), .B(n_27), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_462), .B(n_217), .C(n_215), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_477), .B(n_225), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_472), .B(n_30), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_462), .B(n_215), .C(n_217), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_463), .B(n_215), .C(n_217), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_445), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_451), .B(n_31), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_477), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_479), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_463), .B(n_32), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_456), .B(n_220), .Y(n_537) );
NOR3xp33_ASAP7_75t_SL g538 ( .A(n_446), .B(n_33), .C(n_45), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_478), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_453), .B(n_213), .C(n_200), .D(n_199), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
AOI31xp33_ASAP7_75t_L g542 ( .A1(n_476), .A2(n_442), .A3(n_483), .B(n_480), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_449), .B(n_47), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_542), .A2(n_453), .B(n_474), .Y(n_544) );
NOR2xp33_ASAP7_75t_SL g545 ( .A(n_489), .B(n_474), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_486), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_498), .B(n_457), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_520), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_524), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_521), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_488), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_512), .B(n_450), .Y(n_553) );
OAI322xp33_ASAP7_75t_L g554 ( .A1(n_507), .A2(n_457), .A3(n_450), .B1(n_455), .B2(n_459), .C1(n_480), .C2(n_481), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g555 ( .A1(n_489), .A2(n_469), .A3(n_455), .B1(n_459), .B2(n_481), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g556 ( .A(n_495), .B(n_484), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_518), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
AOI31xp33_ASAP7_75t_L g559 ( .A1(n_490), .A2(n_442), .A3(n_470), .B(n_484), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_512), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_539), .A2(n_475), .B1(n_461), .B2(n_215), .C(n_217), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_501), .B(n_502), .Y(n_563) );
OAI322xp33_ASAP7_75t_L g564 ( .A1(n_525), .A2(n_199), .A3(n_215), .B1(n_217), .B2(n_452), .C1(n_442), .C2(n_447), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_534), .A2(n_461), .B1(n_482), .B2(n_470), .C(n_232), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_494), .A2(n_442), .B1(n_470), .B2(n_461), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_506), .B(n_452), .Y(n_567) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_531), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_531), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_489), .B(n_442), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_541), .Y(n_572) );
NAND2xp33_ASAP7_75t_R g573 ( .A(n_497), .B(n_447), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_538), .A2(n_447), .B1(n_452), .B2(n_251), .C(n_461), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_535), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_512), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_506), .B(n_452), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_514), .B(n_452), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_508), .B(n_447), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_492), .A2(n_470), .B1(n_57), .B2(n_59), .Y(n_580) );
AOI22x1_ASAP7_75t_L g581 ( .A1(n_495), .A2(n_53), .B1(n_61), .B2(n_63), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_504), .A2(n_64), .B1(n_65), .B2(n_66), .C(n_68), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_494), .A2(n_69), .B1(n_72), .B2(n_73), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_514), .B(n_76), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_490), .A2(n_511), .B(n_530), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_531), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_491), .B(n_500), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g588 ( .A1(n_516), .A2(n_487), .B(n_491), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_513), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_493), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_508), .B(n_515), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_556), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_560), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_567), .B(n_515), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_544), .B(n_522), .C(n_517), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_567), .B(n_509), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_503), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_549), .B(n_493), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_550), .B(n_500), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_572), .B(n_503), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_571), .B(n_509), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_580), .A2(n_522), .B(n_517), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_577), .B(n_499), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_548), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_588), .B(n_527), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_551), .B(n_532), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_570), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_545), .A2(n_487), .B1(n_532), .B2(n_536), .Y(n_610) );
AOI321xp33_ASAP7_75t_L g611 ( .A1(n_555), .A2(n_536), .A3(n_543), .B1(n_505), .B2(n_526), .C(n_519), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_562), .B(n_543), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_589), .B(n_537), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_570), .B(n_497), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_559), .A2(n_523), .B(n_529), .Y(n_616) );
CKINVDCx16_ASAP7_75t_R g617 ( .A(n_566), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_577), .B(n_537), .Y(n_618) );
AOI221x1_ASAP7_75t_L g619 ( .A1(n_583), .A2(n_510), .B1(n_540), .B2(n_585), .C(n_576), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_587), .B(n_580), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_553), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_575), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_581), .A2(n_584), .B(n_578), .C(n_568), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_607), .B(n_554), .Y(n_624) );
NOR2xp67_ASAP7_75t_SL g625 ( .A(n_623), .B(n_584), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_607), .A2(n_578), .B(n_564), .C(n_574), .Y(n_626) );
NOR2xp33_ASAP7_75t_SL g627 ( .A(n_592), .B(n_553), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_604), .B(n_579), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_616), .A2(n_582), .B(n_561), .C(n_553), .Y(n_629) );
XNOR2xp5_ASAP7_75t_L g630 ( .A(n_592), .B(n_591), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_593), .A2(n_565), .B(n_569), .C(n_586), .Y(n_631) );
XNOR2x1_ASAP7_75t_L g632 ( .A(n_615), .B(n_591), .Y(n_632) );
OAI31xp33_ASAP7_75t_L g633 ( .A1(n_595), .A2(n_579), .A3(n_573), .B(n_590), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_598), .Y(n_634) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_615), .B(n_573), .Y(n_635) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_609), .B(n_557), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_599), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_605), .B(n_586), .Y(n_638) );
NAND3x1_ASAP7_75t_SL g639 ( .A(n_603), .B(n_557), .C(n_558), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_620), .A2(n_558), .B1(n_618), .B2(n_617), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_636), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_632), .B(n_597), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_624), .A2(n_610), .B1(n_618), .B2(n_601), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_640), .B(n_605), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_637), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_624), .A2(n_619), .B(n_611), .C(n_621), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_633), .A2(n_600), .B(n_596), .C(n_594), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_640), .A2(n_622), .B1(n_606), .B2(n_612), .C(n_594), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_637), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_625), .A2(n_614), .B(n_608), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g651 ( .A(n_627), .B(n_596), .C(n_602), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_629), .A2(n_613), .B(n_626), .C(n_631), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_635), .A2(n_629), .B(n_630), .Y(n_653) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_631), .B(n_639), .C(n_628), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_639), .A2(n_640), .B(n_633), .C(n_624), .Y(n_656) );
AOI211xp5_ASAP7_75t_SL g657 ( .A1(n_638), .A2(n_624), .B(n_623), .C(n_627), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_649), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_649), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_641), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_653), .A2(n_657), .B1(n_652), .B2(n_656), .C(n_646), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_647), .B1(n_650), .B2(n_654), .C(n_648), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_660), .B(n_651), .C(n_642), .D(n_643), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_658), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_664), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_663), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
AOI22xp5_ASAP7_75t_SL g668 ( .A1(n_667), .A2(n_666), .B1(n_660), .B2(n_659), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_662), .B1(n_645), .B2(n_655), .C(n_644), .Y(n_669) );
endmodule