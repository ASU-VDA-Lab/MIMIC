module fake_jpeg_19755_n_259 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_18),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_2),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_2),
.B(n_3),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_5),
.B(n_6),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_59),
.B1(n_23),
.B2(n_20),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_43),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_R g95 ( 
.A(n_49),
.B(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_67),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_62),
.B1(n_69),
.B2(n_38),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_28),
.B(n_21),
.C(n_45),
.Y(n_102)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_31),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_77),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_107),
.B1(n_24),
.B2(n_33),
.Y(n_120)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_48),
.B(n_56),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_93),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_26),
.B1(n_35),
.B2(n_34),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_30),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_26),
.B1(n_45),
.B2(n_38),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_21),
.B(n_35),
.C(n_34),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_24),
.B(n_7),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_28),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_15),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_10),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_123),
.B1(n_128),
.B2(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_32),
.B1(n_24),
.B2(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_32),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_74),
.B1(n_90),
.B2(n_88),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_6),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_104),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_71),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_80),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_85),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_143),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_91),
.B(n_84),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_122),
.B(n_126),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_92),
.B1(n_104),
.B2(n_96),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_124),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_99),
.B(n_84),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_157),
.B(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_104),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_112),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_159),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_112),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_165),
.C(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_118),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_70),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_126),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_83),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_125),
.B1(n_119),
.B2(n_128),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_119),
.B(n_113),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_184),
.B(n_185),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_144),
.B1(n_162),
.B2(n_116),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_165),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_160),
.C(n_158),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_154),
.C(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_143),
.B1(n_126),
.B2(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_182),
.B(n_188),
.C(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_122),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_141),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_153),
.C(n_141),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_126),
.B(n_135),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_202),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_152),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_176),
.C(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_142),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_144),
.B1(n_148),
.B2(n_151),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_212)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_136),
.B1(n_83),
.B2(n_137),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_137),
.B1(n_135),
.B2(n_140),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_180),
.B(n_177),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_183),
.CI(n_171),
.CON(n_207),
.SN(n_207)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_218),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_172),
.C(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_189),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_168),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_167),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_175),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_203),
.B1(n_202),
.B2(n_168),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_209),
.B1(n_208),
.B2(n_178),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_221),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_175),
.B(n_179),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_217),
.B(n_205),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_193),
.C(n_187),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_174),
.B(n_194),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_229),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_140),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_231),
.B1(n_210),
.B2(n_219),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_200),
.B1(n_169),
.B2(n_178),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_224),
.C(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_247),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_246),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_228),
.B(n_225),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_222),
.B(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_246),
.B(n_245),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_248),
.B(n_237),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_241),
.CI(n_238),
.CON(n_257),
.SN(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_254),
.C(n_256),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_257),
.Y(n_259)
);


endmodule