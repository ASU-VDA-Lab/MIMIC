module fake_netlist_6_4845_n_1085 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1085);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1085;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_468;
wire n_372;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_940;
wire n_770;
wire n_795;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_964;
wire n_802;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_116),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_29),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_24),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_56),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_105),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_35),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_153),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_60),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_109),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_17),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_157),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_158),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_150),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_111),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_115),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_142),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_49),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_84),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_93),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_57),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_123),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_110),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_79),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_28),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_118),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_92),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_154),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_8),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_2),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_67),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_178),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_34),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_204),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_260),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_195),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_196),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_196),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_202),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_195),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_197),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_202),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_203),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_246),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_203),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_223),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_267),
.B1(n_275),
.B2(n_268),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_212),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_286),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_263),
.B1(n_251),
.B2(n_224),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_283),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_212),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_229),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_263),
.B1(n_235),
.B2(n_258),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_205),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_289),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_206),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_267),
.A2(n_225),
.B1(n_254),
.B2(n_248),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_208),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_211),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_213),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_297),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_275),
.A2(n_231),
.B1(n_247),
.B2(n_245),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_287),
.B(n_214),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_262),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g367 ( 
.A1(n_266),
.A2(n_219),
.B(n_216),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_318),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_318),
.B(n_279),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_333),
.B(n_313),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_348),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_279),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

AND3x2_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_300),
.C(n_197),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_197),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_361),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_335),
.B(n_297),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_220),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_304),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_361),
.B(n_304),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

AND3x2_ASAP7_75t_L g408 ( 
.A(n_321),
.B(n_1),
.C(n_3),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_306),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_222),
.C(n_221),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_361),
.B(n_306),
.Y(n_415)
);

AND3x2_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_1),
.C(n_3),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_361),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_333),
.B(n_31),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

BUFx6f_ASAP7_75t_SL g421 ( 
.A(n_337),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_325),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_337),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_360),
.B(n_309),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_334),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

NOR2x1p5_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_309),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_311),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_362),
.B(n_311),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

BUFx6f_ASAP7_75t_SL g439 ( 
.A(n_357),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g443 ( 
.A1(n_357),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_443)
);

XOR2x2_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_344),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_367),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_419),
.B(n_398),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_429),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_374),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_371),
.B(n_364),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_402),
.B(n_314),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_314),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_429),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_429),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_R g465 ( 
.A(n_422),
.B(n_327),
.Y(n_465)
);

XNOR2x2_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_363),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_346),
.Y(n_467)
);

XNOR2x2_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_363),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_429),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_423),
.A2(n_345),
.B(n_338),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_346),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_379),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_414),
.B(n_339),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_382),
.B(n_341),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_405),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_391),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_379),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_400),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_432),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_378),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_378),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_380),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_388),
.B(n_366),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_417),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_356),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_422),
.B(n_233),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_341),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_349),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_385),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_385),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_237),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_412),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_349),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_419),
.B(n_358),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_401),
.B(n_359),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_386),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_445),
.A2(n_442),
.B(n_407),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_483),
.B(n_407),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_473),
.B(n_424),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_447),
.B(n_398),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_404),
.Y(n_530)
);

AO22x1_ASAP7_75t_L g531 ( 
.A1(n_525),
.A2(n_443),
.B1(n_239),
.B2(n_240),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_421),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_445),
.A2(n_407),
.B(n_373),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_481),
.B(n_431),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_413),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_421),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_473),
.B(n_389),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_413),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_481),
.B(n_433),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_469),
.B(n_390),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_459),
.B(n_421),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_448),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_487),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_500),
.A2(n_407),
.B(n_373),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_483),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_478),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_355),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_447),
.A2(n_443),
.B1(n_433),
.B2(n_440),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_500),
.A2(n_426),
.B1(n_440),
.B2(n_427),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_509),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_451),
.B(n_390),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_485),
.B(n_390),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_456),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_355),
.C(n_244),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_404),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_495),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_522),
.A2(n_439),
.B1(n_438),
.B2(n_427),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_452),
.B(n_404),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_504),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_467),
.B(n_474),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_453),
.B(n_404),
.Y(n_567)
);

O2A1O1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_523),
.A2(n_418),
.B(n_438),
.C(n_435),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_467),
.B(n_430),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_457),
.A2(n_460),
.B(n_461),
.C(n_458),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_477),
.A2(n_439),
.B1(n_430),
.B2(n_435),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_464),
.B(n_418),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_518),
.Y(n_574)
);

BUFx6f_ASAP7_75t_SL g575 ( 
.A(n_474),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_450),
.B(n_408),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_484),
.A2(n_418),
.B1(n_434),
.B2(n_441),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_511),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_499),
.B(n_409),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_SL g581 ( 
.A(n_483),
.B(n_390),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_466),
.A2(n_441),
.B1(n_434),
.B2(n_409),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_471),
.B(n_392),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_471),
.B(n_392),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

INVx8_ASAP7_75t_L g587 ( 
.A(n_480),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_472),
.B(n_488),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_379),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_537),
.B(n_490),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_SL g591 ( 
.A(n_529),
.B(n_465),
.C(n_505),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_548),
.B(n_492),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_547),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_587),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_SL g596 ( 
.A(n_576),
.B(n_465),
.C(n_468),
.Y(n_596)
);

AOI22x1_ASAP7_75t_L g597 ( 
.A1(n_526),
.A2(n_524),
.B1(n_515),
.B2(n_521),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_566),
.B(n_516),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_587),
.Y(n_599)
);

OR2x6_ASAP7_75t_SL g600 ( 
.A(n_544),
.B(n_444),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_561),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_528),
.B(n_512),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_587),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_534),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_586),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_547),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_SL g608 ( 
.A(n_572),
.B(n_455),
.C(n_502),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_556),
.B(n_454),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_540),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_530),
.B(n_493),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_571),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_557),
.B(n_517),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_579),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_SL g619 ( 
.A(n_572),
.B(n_520),
.C(n_416),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_570),
.A2(n_497),
.B(n_494),
.C(n_501),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_574),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_541),
.B(n_496),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_532),
.B(n_514),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_535),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_550),
.A2(n_508),
.B1(n_507),
.B2(n_503),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_535),
.Y(n_633)
);

INVx3_ASAP7_75t_SL g634 ( 
.A(n_539),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_549),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_580),
.B(n_475),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_543),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_546),
.A2(n_482),
.B(n_411),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_581),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_538),
.B(n_352),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_565),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_569),
.B(n_482),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_589),
.Y(n_643)
);

BUFx4f_ASAP7_75t_L g644 ( 
.A(n_569),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_573),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_527),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_527),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_555),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_589),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_612),
.A2(n_553),
.B(n_533),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_613),
.A2(n_585),
.B(n_583),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_601),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_590),
.A2(n_542),
.B(n_568),
.Y(n_655)
);

NAND2x1_ASAP7_75t_L g656 ( 
.A(n_611),
.B(n_551),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_630),
.Y(n_657)
);

O2A1O1Ixp5_ASAP7_75t_L g658 ( 
.A1(n_624),
.A2(n_531),
.B(n_554),
.C(n_563),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_560),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_607),
.Y(n_660)
);

OAI22x1_ASAP7_75t_L g661 ( 
.A1(n_637),
.A2(n_634),
.B1(n_627),
.B2(n_625),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_638),
.A2(n_567),
.B(n_558),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_597),
.A2(n_567),
.B(n_577),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_645),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_636),
.A2(n_411),
.B(n_392),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_623),
.B(n_582),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_646),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_624),
.A2(n_369),
.B(n_372),
.C(n_370),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_651),
.B(n_369),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_602),
.B(n_352),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_592),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_620),
.A2(n_372),
.B(n_387),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_616),
.A2(n_651),
.B(n_643),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_607),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_643),
.B(n_352),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_632),
.A2(n_387),
.B(n_392),
.Y(n_678)
);

NOR2x1_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_594),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_644),
.B(n_392),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_635),
.B(n_352),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_644),
.A2(n_631),
.B(n_617),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_632),
.A2(n_387),
.B(n_411),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_637),
.B(n_575),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_591),
.B(n_387),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_609),
.B(n_411),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_614),
.B(n_411),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_631),
.A2(n_437),
.B(n_33),
.Y(n_688)
);

AOI21x1_ASAP7_75t_SL g689 ( 
.A1(n_640),
.A2(n_437),
.B(n_4),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_437),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_642),
.A2(n_437),
.B(n_36),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_631),
.A2(n_437),
.B(n_37),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_631),
.A2(n_39),
.B(n_32),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_595),
.B(n_5),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_618),
.B(n_6),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_599),
.B(n_40),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_592),
.A2(n_194),
.B(n_42),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_650),
.B(n_7),
.Y(n_699)
);

BUFx2_ASAP7_75t_R g700 ( 
.A(n_600),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_615),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_611),
.A2(n_43),
.B(n_41),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_596),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_703)
);

AO21x1_ASAP7_75t_L g704 ( 
.A1(n_639),
.A2(n_9),
.B(n_10),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_596),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_615),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_617),
.A2(n_45),
.B(n_44),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_591),
.B(n_11),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_652),
.A2(n_639),
.B(n_647),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_659),
.Y(n_711)
);

AOI221x1_ASAP7_75t_L g712 ( 
.A1(n_705),
.A2(n_605),
.B1(n_593),
.B2(n_608),
.C(n_598),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_653),
.A2(n_649),
.B(n_647),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_654),
.Y(n_714)
);

OA21x2_ASAP7_75t_L g715 ( 
.A1(n_667),
.A2(n_619),
.B(n_626),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_663),
.A2(n_641),
.B(n_628),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_655),
.A2(n_649),
.B(n_647),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_668),
.A2(n_608),
.B1(n_650),
.B2(n_634),
.Y(n_718)
);

NAND2x1_ASAP7_75t_L g719 ( 
.A(n_662),
.B(n_647),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_675),
.A2(n_649),
.B(n_606),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_696),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_666),
.A2(n_649),
.B(n_606),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_665),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_657),
.Y(n_724)
);

AO31x2_ASAP7_75t_L g725 ( 
.A1(n_670),
.A2(n_661),
.A3(n_704),
.B(n_677),
.Y(n_725)
);

OAI22x1_ASAP7_75t_L g726 ( 
.A1(n_703),
.A2(n_603),
.B1(n_610),
.B2(n_646),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_700),
.B(n_621),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_684),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_682),
.A2(n_606),
.B(n_598),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_691),
.A2(n_683),
.B(n_678),
.Y(n_730)
);

BUFx12f_ASAP7_75t_L g731 ( 
.A(n_669),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_672),
.B(n_593),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_679),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_678),
.A2(n_607),
.B(n_594),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_676),
.Y(n_735)
);

AO32x2_ASAP7_75t_L g736 ( 
.A1(n_689),
.A2(n_619),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_701),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_683),
.A2(n_607),
.B(n_47),
.Y(n_738)
);

AO31x2_ASAP7_75t_L g739 ( 
.A1(n_688),
.A2(n_122),
.A3(n_191),
.B(n_190),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_692),
.A2(n_120),
.A3(n_189),
.B(n_188),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_709),
.B(n_12),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_658),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_703),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_656),
.A2(n_18),
.B(n_19),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_664),
.A2(n_125),
.B(n_187),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_660),
.B(n_46),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_698),
.A2(n_126),
.B(n_185),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_702),
.A2(n_708),
.B(n_674),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_671),
.A2(n_124),
.A3(n_184),
.B(n_183),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_680),
.A2(n_193),
.B(n_119),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_676),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_693),
.A2(n_182),
.B(n_113),
.Y(n_752)
);

AO31x2_ASAP7_75t_L g753 ( 
.A1(n_686),
.A2(n_112),
.A3(n_180),
.B(n_177),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_694),
.B(n_20),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_681),
.Y(n_755)
);

CKINVDCx11_ASAP7_75t_R g756 ( 
.A(n_676),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_687),
.A2(n_108),
.A3(n_176),
.B(n_175),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_685),
.A2(n_699),
.B(n_695),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_659),
.B(n_21),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_690),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_104),
.B(n_174),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_707),
.A2(n_100),
.B(n_173),
.Y(n_763)
);

AO21x1_ASAP7_75t_L g764 ( 
.A1(n_662),
.A2(n_673),
.B(n_690),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_660),
.A2(n_22),
.B(n_23),
.Y(n_765)
);

NOR2x1_ASAP7_75t_R g766 ( 
.A(n_697),
.B(n_181),
.Y(n_766)
);

OA21x2_ASAP7_75t_L g767 ( 
.A1(n_667),
.A2(n_121),
.B(n_171),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_665),
.B(n_48),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_657),
.B(n_50),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_663),
.A2(n_129),
.B(n_170),
.Y(n_770)
);

AO31x2_ASAP7_75t_L g771 ( 
.A1(n_667),
.A2(n_99),
.A3(n_169),
.B(n_167),
.Y(n_771)
);

AOI21xp33_ASAP7_75t_L g772 ( 
.A1(n_668),
.A2(n_24),
.B(n_25),
.Y(n_772)
);

OA21x2_ASAP7_75t_L g773 ( 
.A1(n_667),
.A2(n_98),
.B(n_165),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_665),
.B(n_51),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_705),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_714),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_743),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_755),
.B(n_30),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_731),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_723),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_721),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_726),
.A2(n_30),
.B1(n_53),
.B2(n_54),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_712),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_711),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_737),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_716),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_62),
.Y(n_787)
);

BUFx4f_ASAP7_75t_SL g788 ( 
.A(n_759),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_764),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_756),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_754),
.A2(n_744),
.B1(n_772),
.B2(n_765),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_736),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_751),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_758),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_733),
.B(n_66),
.Y(n_796)
);

BUFx4_ASAP7_75t_SL g797 ( 
.A(n_727),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_751),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_715),
.B(n_68),
.Y(n_799)
);

AOI21xp33_ASAP7_75t_L g800 ( 
.A1(n_775),
.A2(n_69),
.B(n_70),
.Y(n_800)
);

BUFx8_ASAP7_75t_L g801 ( 
.A(n_741),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_724),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_735),
.Y(n_803)
);

INVx6_ASAP7_75t_L g804 ( 
.A(n_719),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_715),
.Y(n_805)
);

BUFx12f_ASAP7_75t_L g806 ( 
.A(n_746),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_768),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_760),
.B(n_72),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_749),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_725),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_73),
.Y(n_811)
);

INVx6_ASAP7_75t_L g812 ( 
.A(n_766),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_732),
.B(n_74),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_725),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_753),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_SL g816 ( 
.A1(n_730),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_749),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_728),
.Y(n_818)
);

CKINVDCx11_ASAP7_75t_R g819 ( 
.A(n_761),
.Y(n_819)
);

BUFx8_ASAP7_75t_SL g820 ( 
.A(n_774),
.Y(n_820)
);

INVx6_ASAP7_75t_L g821 ( 
.A(n_722),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_738),
.A2(n_172),
.B1(n_81),
.B2(n_82),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_762),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_729),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_769),
.A2(n_164),
.B1(n_87),
.B2(n_88),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_734),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_739),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_757),
.Y(n_828)
);

INVx6_ASAP7_75t_L g829 ( 
.A(n_720),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_752),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_784),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_818),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_784),
.B(n_771),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_821),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_785),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_826),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_821),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_781),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_821),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_809),
.A2(n_748),
.B(n_745),
.Y(n_840)
);

AO21x2_ASAP7_75t_L g841 ( 
.A1(n_815),
.A2(n_742),
.B(n_710),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_789),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_776),
.B(n_810),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_805),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_828),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_814),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_817),
.B(n_717),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_786),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_827),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_827),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_799),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_793),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_829),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_804),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_799),
.B(n_773),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_829),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_822),
.A2(n_770),
.B(n_747),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_R g858 ( 
.A(n_796),
.B(n_773),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_829),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_SL g860 ( 
.A1(n_824),
.A2(n_767),
.B1(n_763),
.B2(n_750),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_778),
.B(n_713),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_823),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_823),
.B(n_740),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_778),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_803),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_823),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_780),
.B(n_767),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_804),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_811),
.B(n_740),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_804),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_777),
.A2(n_739),
.B1(n_95),
.B2(n_96),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_803),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_868),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_844),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_836),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_831),
.B(n_792),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_840),
.A2(n_783),
.B(n_800),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_842),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_844),
.Y(n_879)
);

AO21x2_ASAP7_75t_L g880 ( 
.A1(n_840),
.A2(n_783),
.B(n_800),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_853),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_853),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_864),
.B(n_792),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_835),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_844),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_871),
.A2(n_819),
.B1(n_777),
.B2(n_782),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_835),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_847),
.B(n_806),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_842),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_845),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_845),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_861),
.B(n_782),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_867),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_852),
.B(n_794),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_834),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_843),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_843),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_852),
.B(n_787),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_857),
.A2(n_822),
.B(n_830),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_846),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_893),
.B(n_833),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_878),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_893),
.B(n_850),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_890),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_890),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_896),
.B(n_850),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_891),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_896),
.B(n_849),
.Y(n_908)
);

INVx3_ASAP7_75t_SL g909 ( 
.A(n_876),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_875),
.B(n_838),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_833),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_891),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_878),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_881),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_881),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_900),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_897),
.B(n_849),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_900),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_889),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_884),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_876),
.B(n_848),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_902),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_909),
.B(n_873),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_909),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_919),
.B(n_915),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_904),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_905),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_921),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_910),
.B(n_883),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_921),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_907),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_901),
.B(n_883),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_915),
.B(n_873),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_913),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_914),
.B(n_888),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_924),
.B(n_908),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_924),
.B(n_908),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_926),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_932),
.B(n_911),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_924),
.B(n_912),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_927),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_929),
.B(n_903),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_932),
.B(n_791),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_923),
.B(n_917),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_922),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_931),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_925),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_933),
.B(n_916),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_948),
.Y(n_950)
);

AND2x4_ASAP7_75t_SL g951 ( 
.A(n_946),
.B(n_925),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_937),
.B(n_933),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_939),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_942),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_948),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_940),
.B(n_936),
.Y(n_956)
);

AO221x2_ASAP7_75t_L g957 ( 
.A1(n_950),
.A2(n_954),
.B1(n_953),
.B2(n_947),
.C(n_955),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_956),
.A2(n_941),
.B1(n_937),
.B2(n_938),
.Y(n_958)
);

OAI22xp33_ASAP7_75t_L g959 ( 
.A1(n_950),
.A2(n_892),
.B1(n_935),
.B2(n_940),
.Y(n_959)
);

INVxp67_ASAP7_75t_SL g960 ( 
.A(n_951),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_SL g961 ( 
.A(n_951),
.B(n_944),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_952),
.B(n_941),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_957),
.B(n_962),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_961),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_958),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_959),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_957),
.B(n_952),
.Y(n_968)
);

AOI221xp5_ASAP7_75t_L g969 ( 
.A1(n_959),
.A2(n_941),
.B1(n_938),
.B2(n_886),
.C(n_949),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_960),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_961),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_961),
.A2(n_936),
.B1(n_892),
.B2(n_949),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_968),
.A2(n_963),
.B(n_970),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_945),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_SL g975 ( 
.A1(n_964),
.A2(n_936),
.B(n_832),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_967),
.Y(n_976)
);

OAI32xp33_ASAP7_75t_L g977 ( 
.A1(n_971),
.A2(n_966),
.A3(n_969),
.B1(n_972),
.B2(n_923),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_963),
.A2(n_949),
.B(n_899),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_965),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_965),
.B(n_945),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_SL g981 ( 
.A1(n_978),
.A2(n_943),
.B(n_930),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_979),
.B(n_928),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_976),
.B(n_779),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_L g984 ( 
.A1(n_977),
.A2(n_816),
.B(n_825),
.C(n_795),
.Y(n_984)
);

NAND3x2_ASAP7_75t_L g985 ( 
.A(n_973),
.B(n_975),
.C(n_980),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_974),
.A2(n_930),
.B1(n_928),
.B2(n_812),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_802),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_934),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_984),
.A2(n_899),
.B(n_934),
.C(n_825),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_985),
.A2(n_801),
.B(n_867),
.Y(n_990)
);

AOI221xp5_ASAP7_75t_L g991 ( 
.A1(n_986),
.A2(n_795),
.B1(n_880),
.B2(n_877),
.C(n_816),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_797),
.Y(n_992)
);

AOI211xp5_ASAP7_75t_L g993 ( 
.A1(n_982),
.A2(n_797),
.B(n_796),
.C(n_808),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_987),
.B(n_801),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_988),
.A2(n_812),
.B1(n_901),
.B2(n_889),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_994),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_995),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_992),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

BUFx8_ASAP7_75t_L g1000 ( 
.A(n_993),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_989),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_991),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_994),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_994),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_994),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_981),
.Y(n_1007)
);

AOI211x1_ASAP7_75t_SL g1008 ( 
.A1(n_997),
.A2(n_872),
.B(n_870),
.C(n_868),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1001),
.A2(n_812),
.B1(n_788),
.B2(n_854),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_996),
.B(n_788),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_SL g1011 ( 
.A(n_999),
.B(n_830),
.C(n_813),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_1000),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_787),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1004),
.B(n_920),
.Y(n_1014)
);

NAND5xp2_ASAP7_75t_L g1015 ( 
.A(n_1005),
.B(n_820),
.C(n_860),
.D(n_807),
.E(n_859),
.Y(n_1015)
);

NOR3x1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.B(n_854),
.C(n_911),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_SL g1017 ( 
.A1(n_1002),
.A2(n_790),
.B1(n_798),
.B2(n_888),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_1012),
.B(n_1000),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1007),
.B(n_807),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1009),
.A2(n_1017),
.B1(n_1010),
.B2(n_1011),
.C(n_1014),
.Y(n_1020)
);

NAND4xp25_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_839),
.C(n_837),
.D(n_834),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1013),
.A2(n_790),
.B1(n_880),
.B2(n_877),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1008),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

AO21x1_ASAP7_75t_L g1025 ( 
.A1(n_1007),
.A2(n_872),
.B(n_858),
.Y(n_1025)
);

NOR4xp25_ASAP7_75t_L g1026 ( 
.A(n_1024),
.B(n_918),
.C(n_794),
.D(n_870),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_1019),
.Y(n_1027)
);

NAND5xp2_ASAP7_75t_L g1028 ( 
.A(n_1020),
.B(n_859),
.C(n_856),
.D(n_898),
.E(n_855),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_1018),
.B(n_798),
.Y(n_1029)
);

NAND5xp2_ASAP7_75t_L g1030 ( 
.A(n_1023),
.B(n_856),
.C(n_898),
.D(n_855),
.E(n_862),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_1022),
.B(n_881),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1025),
.B(n_903),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_1021),
.B(n_882),
.Y(n_1033)
);

OR5x1_ASAP7_75t_L g1034 ( 
.A(n_1021),
.B(n_790),
.C(n_798),
.D(n_865),
.E(n_803),
.Y(n_1034)
);

XNOR2xp5_ASAP7_75t_L g1035 ( 
.A(n_1029),
.B(n_91),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1027),
.B(n_868),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1033),
.B(n_906),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_862),
.C(n_882),
.Y(n_1038)
);

NOR4xp25_ASAP7_75t_L g1039 ( 
.A(n_1032),
.B(n_894),
.C(n_917),
.D(n_906),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1026),
.B(n_882),
.Y(n_1040)
);

AOI221x1_ASAP7_75t_L g1041 ( 
.A1(n_1030),
.A2(n_846),
.B1(n_866),
.B2(n_851),
.C(n_863),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1028),
.B(n_894),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1034),
.A2(n_899),
.B(n_895),
.C(n_834),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_1035),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_1036),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1040),
.A2(n_888),
.B1(n_895),
.B2(n_851),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_1037),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1038),
.B(n_837),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1041),
.B(n_837),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_1043),
.B(n_869),
.C(n_839),
.Y(n_1051)
);

XOR2x1_ASAP7_75t_L g1052 ( 
.A(n_1036),
.B(n_97),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1036),
.B(n_895),
.Y(n_1053)
);

NAND4xp75_ASAP7_75t_L g1054 ( 
.A(n_1040),
.B(n_130),
.C(n_132),
.D(n_133),
.Y(n_1054)
);

AND3x4_ASAP7_75t_L g1055 ( 
.A(n_1036),
.B(n_839),
.C(n_863),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_1036),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1047),
.A2(n_888),
.B1(n_869),
.B2(n_866),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1048),
.B(n_888),
.Y(n_1058)
);

OA21x2_ASAP7_75t_L g1059 ( 
.A1(n_1045),
.A2(n_887),
.B(n_884),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1056),
.A2(n_880),
.B(n_877),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1055),
.A2(n_887),
.B1(n_838),
.B2(n_863),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_1054),
.B(n_880),
.Y(n_1062)
);

NAND4xp75_ASAP7_75t_L g1063 ( 
.A(n_1049),
.B(n_1050),
.C(n_1052),
.D(n_1056),
.Y(n_1063)
);

XNOR2xp5_ASAP7_75t_L g1064 ( 
.A(n_1044),
.B(n_134),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_1064),
.A2(n_1051),
.B1(n_1046),
.B2(n_863),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1057),
.A2(n_1065),
.B1(n_1063),
.B2(n_1062),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_1059),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1060),
.A2(n_877),
.B1(n_841),
.B2(n_847),
.Y(n_1071)
);

AO22x2_ASAP7_75t_L g1072 ( 
.A1(n_1066),
.A2(n_885),
.B1(n_879),
.B2(n_874),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1068),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_841),
.B1(n_847),
.B2(n_879),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_1069),
.C(n_1067),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1076),
.A2(n_1072),
.B1(n_1071),
.B2(n_1074),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_841),
.B1(n_847),
.B2(n_879),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_847),
.B1(n_885),
.B2(n_874),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1079),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1078),
.A2(n_139),
.B(n_140),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_1080),
.A2(n_141),
.B(n_143),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1081),
.A2(n_144),
.B(n_146),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1082),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_1084)
);

AOI211xp5_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_1083),
.B(n_151),
.C(n_152),
.Y(n_1085)
);


endmodule