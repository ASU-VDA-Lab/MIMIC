module fake_ariane_2278_n_2100 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2100);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2100;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_212;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g194 ( 
.A(n_34),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_4),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_41),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_22),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_118),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_63),
.Y(n_215)
);

HB1xp67_ASAP7_75t_SL g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_16),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_126),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_134),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_28),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_177),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_51),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_117),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_161),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_175),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_167),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_52),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_47),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_27),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_187),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_21),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_83),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_23),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_43),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_21),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_35),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_162),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_76),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_77),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_97),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_15),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_119),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_38),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_45),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_80),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_105),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_183),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_112),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_67),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_106),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_81),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_75),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_168),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_160),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_26),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_58),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_107),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_19),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_58),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_140),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_3),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_75),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_80),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_136),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_98),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_7),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_69),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_130),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_36),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_110),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_50),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_9),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_141),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_48),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_147),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_57),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_138),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_111),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_26),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_31),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_62),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_76),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_45),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_71),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_178),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_82),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_54),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_96),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_60),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_189),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_122),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_165),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_18),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_5),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_52),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_20),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_174),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_1),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_70),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_95),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_154),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_94),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_63),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_169),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_40),
.Y(n_350)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_47),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_2),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_103),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_89),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_30),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_171),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_25),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_78),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_39),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_91),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_73),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_73),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_120),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_54),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_142),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_102),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_14),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_101),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_124),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_90),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_129),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_1),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_115),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_51),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_82),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_145),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_48),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_42),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_191),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_9),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_61),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_49),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_60),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_88),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_34),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_132),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_195),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_335),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_205),
.B(n_196),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_248),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_196),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_198),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_198),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_274),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_200),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_200),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_202),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_202),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_203),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_203),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_329),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_229),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_205),
.B(n_0),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_229),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_275),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_295),
.B(n_0),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_335),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_275),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_288),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_268),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_R g417 ( 
.A(n_243),
.B(n_84),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_344),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_268),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_263),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_276),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_276),
.B(n_5),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_294),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_294),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_327),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_345),
.B(n_8),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_327),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_263),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_353),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_270),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_270),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_343),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_290),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_288),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_206),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_238),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_333),
.B(n_8),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_206),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_238),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_210),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_305),
.B(n_10),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_211),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_238),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_290),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_215),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_253),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_355),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_219),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_355),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_253),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_222),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_253),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_224),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_262),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_226),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_359),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_206),
.B(n_11),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_234),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_262),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_236),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_262),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_267),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_267),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_264),
.B(n_11),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_267),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_305),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_244),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_307),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_307),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_240),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_359),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_246),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_249),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_204),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_307),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_313),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_313),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_394),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_421),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_431),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_398),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_407),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_449),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g497 ( 
.A1(n_404),
.A2(n_259),
.B(n_213),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_451),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_390),
.B(n_243),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_245),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_390),
.B(n_269),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_399),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_399),
.B(n_247),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_392),
.B(n_269),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_454),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_457),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_392),
.B(n_269),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_247),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_395),
.B(n_278),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_395),
.B(n_278),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_417),
.B(n_207),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_396),
.B(n_278),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_455),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_459),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_459),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_461),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_478),
.B(n_396),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_471),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_473),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_473),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_465),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_467),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_397),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_470),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_477),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_477),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_472),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_479),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_397),
.B(n_326),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_484),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_400),
.B(n_326),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_400),
.B(n_326),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_401),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_480),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_481),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_485),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_401),
.B(n_348),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_402),
.B(n_207),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_402),
.B(n_348),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_391),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_403),
.B(n_348),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_R g567 ( 
.A(n_437),
.B(n_441),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_413),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_501),
.B(n_228),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_499),
.B(n_213),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_501),
.B(n_228),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_497),
.A2(n_405),
.B(n_403),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_517),
.B(n_444),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_523),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_517),
.B(n_429),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_491),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_440),
.Y(n_579)
);

BUFx6f_ASAP7_75t_SL g580 ( 
.A(n_502),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_540),
.B(n_482),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_447),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_540),
.B(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_415),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_540),
.B(n_409),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_491),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_499),
.B(n_405),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_513),
.B(n_503),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_513),
.B(n_460),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_540),
.B(n_412),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_540),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_540),
.B(n_446),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_496),
.B(n_476),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_524),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_503),
.B(n_406),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_523),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_508),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_213),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_525),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_508),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_514),
.B(n_476),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_524),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_543),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_557),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_494),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_534),
.B(n_450),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_498),
.B(n_423),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_316),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_543),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_490),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_533),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_533),
.Y(n_626)
);

INVx4_ASAP7_75t_SL g627 ( 
.A(n_543),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_490),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_509),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_543),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_503),
.B(n_406),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_509),
.A2(n_340),
.B1(n_469),
.B2(n_255),
.Y(n_634)
);

INVx6_ASAP7_75t_L g635 ( 
.A(n_502),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_504),
.B(n_408),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_543),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_510),
.B(n_408),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_316),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_514),
.B(n_410),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_506),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_534),
.B(n_464),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_514),
.B(n_410),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_506),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_530),
.A2(n_340),
.B1(n_256),
.B2(n_261),
.Y(n_651)
);

INVx3_ASAP7_75t_R g652 ( 
.A(n_541),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_515),
.B(n_416),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_515),
.B(n_416),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_497),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g658 ( 
.A(n_541),
.B(n_313),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_507),
.Y(n_659)
);

NOR2x1p5_ASAP7_75t_L g660 ( 
.A(n_538),
.B(n_240),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_511),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_504),
.B(n_420),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_515),
.B(n_420),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_511),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_519),
.B(n_422),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_519),
.B(n_422),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_511),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_516),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_538),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_539),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_518),
.Y(n_672)
);

INVx6_ASAP7_75t_L g673 ( 
.A(n_502),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_519),
.B(n_551),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_525),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_526),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_424),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_526),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_526),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_531),
.B(n_424),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_551),
.B(n_425),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_526),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_505),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_529),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_551),
.B(n_425),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_497),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_529),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_529),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_539),
.B(n_426),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_492),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_494),
.Y(n_691)
);

INVx4_ASAP7_75t_SL g692 ( 
.A(n_502),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_497),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_497),
.B(n_426),
.Y(n_694)
);

BUFx10_ASAP7_75t_L g695 ( 
.A(n_545),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_518),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_495),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_554),
.B(n_428),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_567),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_545),
.B(n_428),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_495),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_497),
.B(n_432),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_520),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_541),
.B(n_351),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_529),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_537),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_432),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_521),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_439),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_505),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_521),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_549),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_522),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_549),
.B(n_433),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_537),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_537),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_552),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_537),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_554),
.B(n_433),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_625),
.B(n_550),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_658),
.A2(n_512),
.B1(n_556),
.B2(n_505),
.Y(n_724)
);

O2A1O1Ixp5_ASAP7_75t_L g725 ( 
.A1(n_596),
.A2(n_577),
.B(n_590),
.C(n_585),
.Y(n_725)
);

OA22x2_ASAP7_75t_L g726 ( 
.A1(n_634),
.A2(n_553),
.B1(n_560),
.B2(n_550),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_587),
.A2(n_264),
.B1(n_368),
.B2(n_279),
.C(n_280),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_625),
.B(n_553),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_626),
.B(n_560),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_658),
.B(n_567),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_575),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_626),
.B(n_505),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_641),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_714),
.B(n_522),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_579),
.B(n_505),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_689),
.B(n_505),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_700),
.B(n_512),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_716),
.B(n_512),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_581),
.A2(n_556),
.B1(n_563),
.B2(n_512),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_636),
.B(n_512),
.Y(n_741)
);

AOI221xp5_ASAP7_75t_L g742 ( 
.A1(n_574),
.A2(n_271),
.B1(n_273),
.B2(n_258),
.C(n_257),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_577),
.A2(n_556),
.B1(n_563),
.B2(n_512),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_570),
.B(n_556),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_593),
.A2(n_528),
.B(n_527),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_641),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_688),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_711),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_688),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_SL g750 ( 
.A(n_714),
.B(n_419),
.C(n_418),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_720),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_619),
.B(n_565),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_663),
.B(n_556),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_677),
.B(n_556),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_614),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_711),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_704),
.A2(n_442),
.B1(n_443),
.B2(n_436),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_720),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_572),
.B(n_563),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_563),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_571),
.A2(n_683),
.B1(n_620),
.B2(n_680),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_643),
.B(n_653),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_692),
.B(n_563),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_L g765 ( 
.A1(n_596),
.A2(n_563),
.B(n_528),
.C(n_532),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_694),
.A2(n_532),
.B(n_527),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_643),
.B(n_561),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_653),
.B(n_561),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_655),
.B(n_561),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_655),
.B(n_566),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_576),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_698),
.B(n_566),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_719),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_651),
.A2(n_250),
.B1(n_254),
.B2(n_257),
.C(n_258),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_692),
.B(n_245),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_692),
.B(n_548),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_698),
.B(n_566),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_648),
.B(n_535),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_648),
.B(n_535),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_692),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_712),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_720),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_594),
.B(n_536),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_710),
.B(n_565),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_648),
.B(n_536),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_576),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_598),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_592),
.A2(n_442),
.B(n_443),
.C(n_436),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_571),
.A2(n_289),
.B1(n_544),
.B2(n_542),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_666),
.B(n_542),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_666),
.B(n_544),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_598),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_620),
.B(n_548),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_605),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_710),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_646),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_666),
.B(n_546),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_683),
.B(n_316),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_712),
.B(n_546),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_712),
.B(n_548),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_605),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_646),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_691),
.B(n_569),
.C(n_225),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_718),
.B(n_555),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

NOR2x2_ASAP7_75t_L g808 ( 
.A(n_704),
.B(n_434),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_683),
.B(n_316),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_571),
.A2(n_289),
.B1(n_558),
.B2(n_547),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_600),
.B(n_547),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_681),
.B(n_708),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_718),
.B(n_555),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_690),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_578),
.B(n_569),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_681),
.B(n_558),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_608),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_608),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_571),
.A2(n_559),
.B1(n_568),
.B2(n_564),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_580),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_718),
.B(n_555),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_681),
.B(n_559),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_706),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_708),
.B(n_564),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_597),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_656),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_674),
.B(n_568),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_708),
.B(n_555),
.Y(n_828)
);

NOR2x1_ASAP7_75t_L g829 ( 
.A(n_654),
.B(n_487),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_624),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_580),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_706),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_674),
.B(n_208),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_722),
.B(n_500),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_722),
.A2(n_225),
.B(n_235),
.C(n_208),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_622),
.B(n_259),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_582),
.A2(n_235),
.B1(n_250),
.B2(n_254),
.C(n_271),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_618),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_606),
.A2(n_500),
.B(n_284),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_615),
.A2(n_231),
.B1(n_194),
.B2(n_351),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_722),
.B(n_500),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_571),
.A2(n_216),
.B1(n_199),
.B2(n_209),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_635),
.B(n_216),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_578),
.B(n_492),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_628),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_571),
.A2(n_303),
.B1(n_291),
.B2(n_283),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_635),
.B(n_260),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_654),
.B(n_486),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_683),
.B(n_386),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_635),
.B(n_265),
.Y(n_850)
);

NOR2x1p5_ASAP7_75t_L g851 ( 
.A(n_670),
.B(n_281),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_638),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_615),
.A2(n_231),
.B1(n_194),
.B2(n_386),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_718),
.B(n_259),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_718),
.B(n_284),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_697),
.B(n_493),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_615),
.B(n_500),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_704),
.B(n_273),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_664),
.B(n_500),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_659),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_667),
.B(n_279),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_589),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_707),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_662),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_635),
.B(n_287),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_SL g866 ( 
.A(n_697),
.B(n_493),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_L g867 ( 
.A(n_622),
.B(n_293),
.C(n_292),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_704),
.B(n_280),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_583),
.B(n_284),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_583),
.B(n_286),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_683),
.A2(n_266),
.B1(n_389),
.B2(n_282),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_685),
.B(n_285),
.Y(n_872)
);

AND3x1_ASAP7_75t_L g873 ( 
.A(n_652),
.B(n_297),
.C(n_285),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_669),
.B(n_297),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_672),
.B(n_310),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_311),
.C(n_310),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_583),
.B(n_286),
.Y(n_877)
);

AO22x1_ASAP7_75t_L g878 ( 
.A1(n_699),
.A2(n_339),
.B1(n_296),
.B2(n_388),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_311),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_670),
.B(n_435),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_614),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_703),
.B(n_318),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_705),
.A2(n_338),
.B(n_373),
.C(n_318),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_660),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_709),
.B(n_328),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_629),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_713),
.B(n_328),
.Y(n_887)
);

INVx6_ASAP7_75t_L g888 ( 
.A(n_629),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_583),
.B(n_286),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_715),
.B(n_331),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_583),
.B(n_298),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_683),
.B(n_331),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_707),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_591),
.B(n_298),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_823),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_814),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_807),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_763),
.Y(n_898)
);

OR2x6_ASAP7_75t_L g899 ( 
.A(n_781),
.B(n_600),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_762),
.B(n_629),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_807),
.B(n_671),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_757),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_807),
.B(n_671),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_751),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_888),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_784),
.B(n_673),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_880),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_618),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_807),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_612),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_826),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_826),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_772),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_787),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_733),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_788),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_784),
.B(n_673),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_793),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_823),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_723),
.B(n_701),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_826),
.B(n_656),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_826),
.B(n_671),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_795),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_755),
.B(n_673),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_771),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_728),
.B(n_621),
.C(n_301),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_892),
.A2(n_580),
.B1(n_673),
.B2(n_612),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_803),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_827),
.B(n_695),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_782),
.B(n_695),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_817),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_736),
.B(n_612),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_782),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_729),
.B(n_695),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_832),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_737),
.B(n_612),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_758),
.B(n_591),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_843),
.A2(n_612),
.B1(n_640),
.B2(n_584),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_820),
.B(n_831),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_832),
.Y(n_941)
);

NOR3xp33_ASAP7_75t_SL g942 ( 
.A(n_750),
.B(n_302),
.C(n_300),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_818),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_748),
.B(n_652),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_848),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_746),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_830),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_811),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_845),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_888),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_888),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_796),
.B(n_690),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_831),
.B(n_612),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_SL g954 ( 
.A(n_835),
.B(n_306),
.C(n_304),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_852),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_797),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_860),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_815),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_SL g959 ( 
.A(n_886),
.B(n_599),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_771),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_864),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_SL g962 ( 
.A(n_835),
.B(n_314),
.C(n_308),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_771),
.Y(n_963)
);

AND3x1_ASAP7_75t_L g964 ( 
.A(n_866),
.B(n_368),
.C(n_338),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_863),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_771),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_798),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_834),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_785),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_841),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_828),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_812),
.B(n_609),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_838),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_825),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_827),
.B(n_610),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_827),
.B(n_892),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_804),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_863),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_893),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_767),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_768),
.B(n_631),
.Y(n_981)
);

NOR2x1_ASAP7_75t_R g982 ( 
.A(n_730),
.B(n_603),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_774),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_769),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_770),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_773),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_797),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_SL g988 ( 
.A1(n_726),
.A2(n_453),
.B1(n_456),
.B2(n_438),
.Y(n_988)
);

BUFx2_ASAP7_75t_SL g989 ( 
.A(n_734),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_892),
.A2(n_602),
.B1(n_588),
.B2(n_458),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_844),
.Y(n_991)
);

AND2x6_ASAP7_75t_SL g992 ( 
.A(n_858),
.B(n_373),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_883),
.B(n_323),
.C(n_322),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_778),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_843),
.B(n_610),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_856),
.B(n_694),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_838),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_801),
.A2(n_596),
.B1(n_609),
.B2(n_686),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_735),
.B(n_613),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_858),
.A2(n_483),
.B1(n_468),
.B2(n_686),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_779),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_873),
.Y(n_1002)
);

AO22x1_ASAP7_75t_L g1003 ( 
.A1(n_805),
.A2(n_358),
.B1(n_324),
.B2(n_365),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_819),
.B(n_591),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_811),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_780),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_753),
.B(n_640),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_833),
.B(n_609),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_868),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_862),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_858),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_730),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_786),
.B(n_613),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_791),
.B(n_644),
.Y(n_1015)
);

AO22x1_ASAP7_75t_L g1016 ( 
.A1(n_876),
.A2(n_325),
.B1(n_337),
.B2(n_342),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_792),
.B(n_644),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_833),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_738),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_L g1020 ( 
.A(n_836),
.Y(n_1020)
);

BUFx4f_ASAP7_75t_SL g1021 ( 
.A(n_884),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_738),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_747),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_747),
.Y(n_1024)
);

BUFx5_ASAP7_75t_L g1025 ( 
.A(n_836),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_764),
.B(n_656),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_799),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_766),
.B(n_591),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_749),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_742),
.A2(n_686),
.B1(n_656),
.B2(n_693),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_833),
.B(n_675),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_749),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_878),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_847),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_752),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_752),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_759),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_816),
.B(n_675),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_822),
.B(n_676),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_824),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_800),
.B(n_573),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_759),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_783),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_783),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_765),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_857),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_808),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_806),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_739),
.A2(n_721),
.B(n_717),
.C(n_678),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_732),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_874),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_724),
.B(n_678),
.Y(n_1053)
);

NOR2x1_ASAP7_75t_R g1054 ( 
.A(n_739),
.B(n_330),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_741),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_754),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_790),
.B(n_693),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_847),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_764),
.B(n_627),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_SL g1060 ( 
.A(n_883),
.B(n_350),
.C(n_346),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_810),
.B(n_591),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_829),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_809),
.B(n_573),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_849),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_861),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_850),
.B(n_633),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_801),
.B(n_601),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_726),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_875),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_879),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_777),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_882),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_761),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_744),
.B(n_679),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_851),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_837),
.B(n_679),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_777),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_744),
.B(n_682),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_885),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_727),
.B(n_356),
.C(n_352),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_SL g1081 ( 
.A(n_775),
.B(n_362),
.C(n_360),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_806),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_813),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_887),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_760),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_890),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_760),
.B(n_743),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1028),
.A2(n_870),
.B(n_869),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_907),
.A2(n_881),
.B(n_756),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1028),
.A2(n_725),
.B(n_745),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_SL g1091 ( 
.A1(n_918),
.A2(n_789),
.B1(n_850),
.B2(n_865),
.C(n_872),
.Y(n_1091)
);

OAI22x1_ASAP7_75t_L g1092 ( 
.A1(n_1002),
.A2(n_842),
.B1(n_794),
.B2(n_865),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1065),
.B(n_840),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_898),
.B(n_853),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1001),
.B(n_1006),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_L g1096 ( 
.A(n_987),
.B(n_794),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_999),
.A2(n_821),
.B(n_813),
.Y(n_1097)
);

OA21x2_ASAP7_75t_L g1098 ( 
.A1(n_1067),
.A2(n_839),
.B(n_789),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_897),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_947),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1027),
.B(n_740),
.Y(n_1101)
);

AO31x2_ASAP7_75t_L g1102 ( 
.A1(n_995),
.A2(n_721),
.A3(n_682),
.B(n_684),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1045),
.A2(n_821),
.B(n_854),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1040),
.B(n_776),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_980),
.B(n_776),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_895),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_969),
.B(n_194),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_984),
.B(n_684),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_1067),
.A2(n_855),
.B(n_854),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_933),
.A2(n_802),
.B(n_702),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1048),
.A2(n_687),
.A3(n_717),
.B(n_595),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1045),
.A2(n_855),
.B(n_870),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_937),
.A2(n_702),
.B(n_694),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1061),
.A2(n_889),
.B(n_877),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1048),
.A2(n_894),
.B(n_889),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_921),
.A2(n_871),
.B1(n_846),
.B2(n_867),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_1083),
.A2(n_687),
.A3(n_623),
.B(n_617),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_985),
.B(n_702),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1083),
.A2(n_604),
.A3(n_586),
.B(n_595),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1074),
.A2(n_891),
.B(n_877),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1061),
.A2(n_894),
.B(n_891),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_976),
.B(n_627),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1078),
.A2(n_604),
.B(n_586),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_959),
.A2(n_693),
.B1(n_489),
.B2(n_488),
.C(n_379),
.Y(n_1124)
);

NAND2xp33_ASAP7_75t_L g1125 ( 
.A(n_922),
.B(n_601),
.Y(n_1125)
);

OAI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_935),
.A2(n_1080),
.B(n_1081),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_925),
.A2(n_616),
.B(n_607),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1002),
.B(n_194),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_998),
.A2(n_970),
.B(n_968),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_976),
.B(n_627),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_981),
.A2(n_616),
.B(n_607),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1010),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_986),
.B(n_633),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_1087),
.A2(n_299),
.B(n_298),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_994),
.B(n_633),
.Y(n_1135)
);

BUFx2_ASAP7_75t_SL g1136 ( 
.A(n_950),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_1087),
.A2(n_317),
.B(n_299),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_949),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1058),
.B(n_693),
.Y(n_1139)
);

NAND2x1_ASAP7_75t_L g1140 ( 
.A(n_922),
.B(n_909),
.Y(n_1140)
);

BUFx2_ASAP7_75t_R g1141 ( 
.A(n_906),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_906),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1050),
.A2(n_623),
.B(n_617),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1052),
.B(n_693),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_895),
.Y(n_1145)
);

OAI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_958),
.A2(n_376),
.B(n_363),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1014),
.A2(n_632),
.B(n_630),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_SL g1148 ( 
.A1(n_900),
.A2(n_632),
.B(n_630),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_897),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_920),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1004),
.A2(n_642),
.B(n_645),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1020),
.B(n_601),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1069),
.B(n_645),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1004),
.A2(n_642),
.B(n_647),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_922),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_958),
.A2(n_944),
.B(n_1049),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_902),
.A2(n_649),
.B(n_647),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_976),
.B(n_627),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_902),
.A2(n_650),
.B(n_649),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1070),
.B(n_650),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1072),
.B(n_657),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1020),
.A2(n_379),
.B1(n_375),
.B2(n_380),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_668),
.B(n_665),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1020),
.A2(n_375),
.B1(n_384),
.B2(n_383),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1063),
.A2(n_668),
.B(n_665),
.Y(n_1165)
);

AO22x1_ASAP7_75t_L g1166 ( 
.A1(n_1009),
.A2(n_382),
.B1(n_489),
.B2(n_488),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1015),
.A2(n_1038),
.B(n_1017),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1033),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_904),
.A2(n_661),
.B(n_657),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_975),
.A2(n_601),
.B(n_637),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1079),
.A2(n_317),
.B(n_299),
.C(n_370),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_945),
.B(n_231),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_SL g1173 ( 
.A1(n_1005),
.A2(n_1037),
.B(n_966),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_920),
.A2(n_661),
.A3(n_370),
.B(n_317),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1021),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_952),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_940),
.B(n_601),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1033),
.Y(n_1178)
);

AOI31xp67_ASAP7_75t_L g1179 ( 
.A1(n_900),
.A2(n_370),
.A3(n_637),
.B(n_197),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_948),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1084),
.A2(n_386),
.B(n_637),
.C(n_197),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_904),
.A2(n_637),
.B(n_197),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1039),
.A2(n_637),
.B(n_387),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_971),
.A2(n_381),
.B(n_272),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_948),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_897),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1005),
.A2(n_12),
.B(n_13),
.Y(n_1187)
);

OAI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_946),
.A2(n_386),
.B(n_378),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1086),
.B(n_12),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1073),
.A2(n_386),
.B(n_197),
.C(n_374),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1073),
.A2(n_386),
.B(n_197),
.C(n_372),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_903),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1055),
.A2(n_197),
.B(n_369),
.C(n_367),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1037),
.A2(n_13),
.B(n_15),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_936),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1055),
.A2(n_377),
.B(n_366),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_955),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_975),
.B(n_17),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1008),
.A2(n_364),
.B1(n_361),
.B2(n_357),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_950),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1031),
.B(n_17),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1055),
.A2(n_354),
.B(n_349),
.C(n_347),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1008),
.A2(n_341),
.B1(n_336),
.B2(n_334),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_936),
.A2(n_231),
.A3(n_19),
.B(n_20),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_908),
.B(n_18),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_923),
.A2(n_108),
.B(n_192),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1031),
.B(n_1018),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_951),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1056),
.A2(n_332),
.B(n_320),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1053),
.B(n_22),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_952),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_923),
.A2(n_965),
.B(n_941),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_941),
.A2(n_100),
.B(n_186),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_965),
.A2(n_99),
.B(n_179),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1056),
.A2(n_319),
.B(n_315),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1053),
.B(n_23),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_959),
.A2(n_85),
.B(n_176),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_978),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1011),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1008),
.A2(n_312),
.B1(n_309),
.B2(n_277),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_979),
.A2(n_93),
.B(n_116),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1056),
.A2(n_1064),
.B(n_931),
.Y(n_1222)
);

CKINVDCx8_ASAP7_75t_R g1223 ( 
.A(n_992),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_979),
.A2(n_24),
.A3(n_29),
.B(n_30),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_951),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1064),
.B(n_252),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_991),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1064),
.A2(n_251),
.B(n_242),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1085),
.B(n_24),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1085),
.B(n_31),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1013),
.A2(n_32),
.A3(n_33),
.B(n_36),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_930),
.B(n_957),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1076),
.A2(n_241),
.B(n_239),
.C(n_237),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1064),
.A2(n_233),
.B(n_232),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1064),
.A2(n_230),
.B1(n_227),
.B2(n_223),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_948),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1013),
.A2(n_163),
.B(n_128),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_938),
.A2(n_173),
.B(n_131),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1007),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_930),
.B(n_33),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_940),
.B(n_156),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1051),
.A2(n_221),
.B(n_220),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_938),
.A2(n_218),
.B(n_217),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_983),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_961),
.B(n_37),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1012),
.B(n_37),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_974),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_896),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1019),
.A2(n_149),
.B(n_137),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1192),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1129),
.A2(n_939),
.B(n_931),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1095),
.B(n_967),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1167),
.A2(n_972),
.B(n_1051),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1126),
.A2(n_954),
.B(n_962),
.C(n_927),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1125),
.A2(n_912),
.B(n_910),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1134),
.A2(n_1026),
.B(n_1029),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1090),
.A2(n_1019),
.B(n_1024),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1090),
.A2(n_1044),
.B(n_1024),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1227),
.B(n_977),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1100),
.Y(n_1260)
);

NAND2x1_ASAP7_75t_L g1261 ( 
.A(n_1173),
.B(n_922),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1151),
.A2(n_1043),
.B(n_1042),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1241),
.B(n_1210),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1151),
.A2(n_1043),
.B(n_1042),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1154),
.A2(n_1044),
.B(n_1029),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_1155),
.B(n_897),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1137),
.A2(n_1026),
.B(n_901),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1239),
.B(n_916),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1088),
.A2(n_1026),
.B(n_905),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1186),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1154),
.A2(n_1051),
.B(n_997),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1111),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1200),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1184),
.A2(n_972),
.B(n_1030),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1182),
.A2(n_973),
.B(n_997),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1216),
.B(n_996),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1239),
.B(n_1232),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1138),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1106),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1116),
.A2(n_990),
.B(n_993),
.C(n_1060),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1181),
.A2(n_1066),
.B(n_932),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1241),
.B(n_996),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1207),
.B(n_1012),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1157),
.A2(n_973),
.B(n_997),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_973),
.B(n_914),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1159),
.A2(n_924),
.B(n_915),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1181),
.A2(n_919),
.B(n_943),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1155),
.B(n_897),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1229),
.A2(n_1046),
.B(n_972),
.C(n_989),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1197),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1247),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1229),
.A2(n_1046),
.B(n_1068),
.C(n_929),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1159),
.A2(n_917),
.B(n_934),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1175),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1169),
.A2(n_934),
.B(n_928),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1132),
.A2(n_1000),
.B1(n_964),
.B2(n_934),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_922),
.B(n_1025),
.Y(n_1298)
);

AND2x2_ASAP7_75t_SL g1299 ( 
.A(n_1125),
.B(n_1241),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1155),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1200),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1233),
.A2(n_1196),
.B(n_1089),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1155),
.B(n_910),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1219),
.B(n_1244),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1111),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_1122),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1180),
.B(n_940),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1114),
.A2(n_1025),
.B(n_910),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1091),
.A2(n_1062),
.B(n_1059),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1145),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_L g1311 ( 
.A(n_1156),
.B(n_1016),
.C(n_1054),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1246),
.A2(n_896),
.B1(n_1009),
.B2(n_1075),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1114),
.A2(n_1025),
.B(n_910),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1162),
.A2(n_988),
.B1(n_1025),
.B2(n_1057),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1111),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1092),
.A2(n_1082),
.B1(n_1037),
.B2(n_1022),
.C(n_1032),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1177),
.B(n_1034),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1121),
.A2(n_1025),
.B(n_910),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1233),
.A2(n_956),
.B(n_953),
.C(n_911),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1111),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1121),
.A2(n_1025),
.B(n_912),
.Y(n_1321)
);

AOI21xp33_ASAP7_75t_L g1322 ( 
.A1(n_1094),
.A2(n_982),
.B(n_1077),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1112),
.A2(n_1059),
.B(n_942),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1112),
.A2(n_1025),
.B(n_912),
.Y(n_1324)
);

OAI21xp33_ASAP7_75t_L g1325 ( 
.A1(n_1146),
.A2(n_956),
.B(n_1036),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1150),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1150),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1103),
.A2(n_912),
.B(n_913),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1219),
.B(n_1003),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1212),
.A2(n_912),
.B(n_913),
.Y(n_1330)
);

CKINVDCx6p67_ASAP7_75t_R g1331 ( 
.A(n_1208),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1195),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1248),
.B(n_987),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1141),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1195),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1144),
.A2(n_1222),
.B(n_1097),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1243),
.A2(n_1026),
.B(n_1059),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1221),
.A2(n_913),
.B(n_1057),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1122),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1101),
.B(n_1036),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1122),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1218),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1093),
.A2(n_1047),
.B1(n_1057),
.B2(n_911),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1245),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1221),
.A2(n_913),
.B(n_1057),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1117),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1176),
.A2(n_911),
.B1(n_953),
.B2(n_1034),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1142),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1117),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1208),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1164),
.A2(n_1057),
.B1(n_1034),
.B2(n_953),
.Y(n_1351)
);

INVx8_ASAP7_75t_L g1352 ( 
.A(n_1130),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1237),
.A2(n_913),
.B(n_1057),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1117),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1237),
.A2(n_1082),
.B(n_1035),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1171),
.A2(n_909),
.B(n_212),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1117),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1171),
.A2(n_966),
.A3(n_1082),
.B(n_1022),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1124),
.A2(n_1035),
.B(n_909),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1163),
.A2(n_1082),
.B(n_1035),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1186),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1223),
.A2(n_899),
.B1(n_1035),
.B2(n_966),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1119),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1189),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1119),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1140),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1180),
.B(n_960),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1119),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1119),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1176),
.A2(n_1077),
.B1(n_1071),
.B2(n_899),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1249),
.A2(n_1032),
.B(n_1023),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1238),
.A2(n_1032),
.B(n_1023),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1128),
.B(n_1022),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1115),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1242),
.A2(n_960),
.B(n_899),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1130),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1098),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1238),
.A2(n_1032),
.B(n_1023),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1213),
.A2(n_1032),
.B(n_1023),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1142),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1102),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1202),
.A2(n_960),
.B(n_214),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1214),
.A2(n_1023),
.B(n_1022),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1185),
.B(n_960),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1102),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1211),
.A2(n_1077),
.B1(n_1071),
.B2(n_963),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1185),
.B(n_1077),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1102),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1190),
.A2(n_1077),
.A3(n_1071),
.B(n_963),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1211),
.A2(n_1071),
.B1(n_963),
.B2(n_926),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1107),
.B(n_1071),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1230),
.A2(n_1105),
.B(n_1104),
.C(n_1193),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1168),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1225),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1099),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1170),
.A2(n_926),
.B(n_133),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1153),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1131),
.A2(n_926),
.B(n_201),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1172),
.B(n_39),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1205),
.A2(n_1168),
.B1(n_1178),
.B2(n_1199),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1163),
.A2(n_123),
.B(n_41),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1193),
.A2(n_40),
.B(n_42),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1098),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1099),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1225),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_SL g1406 ( 
.A(n_1178),
.B(n_1130),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1120),
.A2(n_43),
.B(n_44),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1158),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1102),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1099),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1206),
.A2(n_44),
.B(n_49),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1177),
.B(n_81),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1198),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1123),
.A2(n_53),
.B(n_56),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1160),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1147),
.A2(n_57),
.B(n_59),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1348),
.Y(n_1417)
);

CKINVDCx16_ASAP7_75t_R g1418 ( 
.A(n_1406),
.Y(n_1418)
);

CKINVDCx8_ASAP7_75t_R g1419 ( 
.A(n_1348),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1295),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1352),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1260),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1371),
.A2(n_1127),
.B(n_1143),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1252),
.B(n_1250),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1278),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1352),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1263),
.B(n_1096),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1311),
.A2(n_1240),
.B1(n_1166),
.B2(n_1220),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1291),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1295),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1292),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1310),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1314),
.A2(n_1201),
.B1(n_1188),
.B2(n_1108),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1297),
.A2(n_1203),
.B1(n_1236),
.B2(n_1152),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1295),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1381),
.A2(n_1165),
.B(n_1190),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1280),
.A2(n_1236),
.B1(n_1152),
.B2(n_1136),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1334),
.Y(n_1439)
);

INVx5_ASAP7_75t_SL g1440 ( 
.A(n_1331),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1299),
.A2(n_1139),
.B1(n_1133),
.B2(n_1135),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1393),
.A2(n_1177),
.B1(n_1158),
.B2(n_1235),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_SL g1443 ( 
.A(n_1254),
.B(n_1217),
.C(n_1215),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1332),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1299),
.A2(n_1191),
.B1(n_1118),
.B2(n_1209),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1293),
.B(n_1191),
.C(n_1228),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1402),
.B(n_1234),
.C(n_1183),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1381),
.A2(n_1165),
.B(n_1226),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1364),
.A2(n_1161),
.B1(n_1194),
.B2(n_1187),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1277),
.B(n_1099),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1263),
.A2(n_1226),
.B1(n_1110),
.B2(n_1158),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1344),
.A2(n_1113),
.B1(n_1109),
.B2(n_1149),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1304),
.B(n_1149),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1279),
.Y(n_1454)
);

AO31x2_ASAP7_75t_L g1455 ( 
.A1(n_1316),
.A2(n_1179),
.A3(n_1174),
.B(n_1148),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1312),
.A2(n_1109),
.B1(n_1149),
.B2(n_1204),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1276),
.A2(n_1149),
.B1(n_1204),
.B2(n_1224),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1400),
.A2(n_1231),
.B1(n_1224),
.B2(n_1204),
.C(n_65),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1279),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1276),
.A2(n_1204),
.B1(n_1224),
.B2(n_1231),
.Y(n_1460)
);

INVx8_ASAP7_75t_L g1461 ( 
.A(n_1352),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1413),
.A2(n_1231),
.B1(n_1224),
.B2(n_1174),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1282),
.A2(n_1231),
.B1(n_1174),
.B2(n_62),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1412),
.B(n_59),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1284),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1301),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1282),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1274),
.A2(n_1340),
.B1(n_1343),
.B2(n_1351),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1302),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1255),
.A2(n_72),
.B(n_77),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1376),
.B(n_78),
.Y(n_1471)
);

NOR2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1393),
.B(n_79),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1350),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1342),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1350),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1283),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1399),
.A2(n_1392),
.B1(n_1329),
.B2(n_1322),
.C(n_1382),
.Y(n_1477)
);

CKINVDCx6p67_ASAP7_75t_R g1478 ( 
.A(n_1331),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1283),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1352),
.B(n_1300),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1268),
.A2(n_1284),
.B1(n_1290),
.B2(n_1333),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1251),
.A2(n_1253),
.B(n_1336),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1316),
.A2(n_1385),
.A3(n_1388),
.B(n_1409),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1259),
.B(n_1412),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1380),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1281),
.A2(n_1356),
.B1(n_1391),
.B2(n_1362),
.Y(n_1486)
);

AOI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1325),
.A2(n_1356),
.B(n_1281),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1373),
.B(n_1405),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1340),
.A2(n_1415),
.B1(n_1397),
.B2(n_1281),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1326),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1347),
.A2(n_1319),
.B(n_1307),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1376),
.B(n_1339),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1338),
.A2(n_1353),
.B(n_1345),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1273),
.B(n_1394),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1273),
.B(n_1394),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1270),
.B(n_1361),
.Y(n_1496)
);

NOR3xp33_ASAP7_75t_L g1497 ( 
.A(n_1317),
.B(n_1359),
.C(n_1407),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1306),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1326),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1309),
.A2(n_1385),
.B1(n_1388),
.B2(n_1409),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1376),
.B(n_1339),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1339),
.B(n_1341),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1341),
.A2(n_1307),
.B1(n_1386),
.B2(n_1390),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1387),
.A2(n_1306),
.B1(n_1408),
.B2(n_1341),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1376),
.B(n_1387),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1387),
.B(n_1367),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1327),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1309),
.A2(n_1361),
.B1(n_1270),
.B2(n_1306),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1327),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1335),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1287),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1408),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1272),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1309),
.A2(n_1401),
.B1(n_1315),
.B2(n_1320),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1257),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_R g1516 ( 
.A(n_1300),
.B(n_1408),
.Y(n_1516)
);

INVx4_ASAP7_75t_SL g1517 ( 
.A(n_1300),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1287),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1375),
.A2(n_1300),
.B1(n_1356),
.B2(n_1370),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1367),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1367),
.A2(n_1384),
.B1(n_1323),
.B2(n_1288),
.Y(n_1521)
);

NAND2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1300),
.B(n_1366),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1401),
.A2(n_1315),
.B1(n_1320),
.B2(n_1305),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1384),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1395),
.B(n_1404),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1404),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1261),
.A2(n_1298),
.B(n_1355),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1395),
.B(n_1410),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1323),
.B(n_1305),
.C(n_1272),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1401),
.A2(n_1288),
.B1(n_1349),
.B2(n_1357),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1410),
.B(n_1288),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1257),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1349),
.A2(n_1357),
.B1(n_1346),
.B2(n_1354),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1414),
.A2(n_1407),
.B(n_1416),
.C(n_1338),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1366),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1363),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1266),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1257),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1266),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1541)
);

INVx8_ASAP7_75t_L g1542 ( 
.A(n_1366),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1266),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1346),
.A2(n_1354),
.B1(n_1363),
.B2(n_1369),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_SL g1545 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1365),
.A2(n_1368),
.A3(n_1369),
.B(n_1374),
.Y(n_1546)
);

CKINVDCx6p67_ASAP7_75t_R g1547 ( 
.A(n_1289),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1398),
.Y(n_1548)
);

NAND2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1308),
.B(n_1313),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1414),
.B(n_1416),
.C(n_1411),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1298),
.A2(n_1353),
.B(n_1345),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1289),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1323),
.B(n_1303),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1360),
.A2(n_1411),
.B1(n_1365),
.B2(n_1368),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1358),
.B(n_1389),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1289),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1303),
.B(n_1269),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1377),
.B(n_1403),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1377),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1303),
.A2(n_1267),
.B1(n_1374),
.B2(n_1269),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1389),
.B(n_1358),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_SL g1562 ( 
.A(n_1337),
.B(n_1358),
.C(n_1389),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1389),
.B(n_1358),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1358),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1286),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1389),
.B(n_1286),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1258),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1308),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1256),
.A2(n_1294),
.B1(n_1296),
.B2(n_1285),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1313),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1294),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1318),
.B(n_1321),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1296),
.A2(n_1258),
.B1(n_1262),
.B2(n_1264),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1425),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1469),
.A2(n_1262),
.B1(n_1264),
.B2(n_1265),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1465),
.A2(n_1428),
.B1(n_1477),
.B2(n_1467),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1465),
.A2(n_1265),
.B1(n_1318),
.B2(n_1321),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_SL g1578 ( 
.A1(n_1467),
.A2(n_1396),
.B(n_1378),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1434),
.A2(n_1418),
.B1(n_1433),
.B2(n_1481),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1433),
.A2(n_1324),
.B1(n_1271),
.B2(n_1378),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1458),
.A2(n_1324),
.B1(n_1271),
.B2(n_1372),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1468),
.A2(n_1464),
.B1(n_1463),
.B2(n_1472),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1438),
.A2(n_1372),
.B1(n_1379),
.B2(n_1383),
.C(n_1328),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1485),
.A2(n_1285),
.B1(n_1275),
.B2(n_1328),
.Y(n_1584)
);

BUFx12f_ASAP7_75t_L g1585 ( 
.A(n_1439),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1482),
.A2(n_1330),
.B(n_1275),
.Y(n_1586)
);

OAI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1443),
.A2(n_1330),
.B(n_1449),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1468),
.A2(n_1463),
.B1(n_1484),
.B2(n_1446),
.Y(n_1588)
);

BUFx12f_ASAP7_75t_L g1589 ( 
.A(n_1439),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1424),
.B(n_1488),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_L g1591 ( 
.A(n_1470),
.B(n_1548),
.C(n_1456),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1450),
.B(n_1453),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1422),
.A2(n_1460),
.B1(n_1457),
.B2(n_1447),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1437),
.B(n_1429),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1440),
.A2(n_1478),
.B1(n_1449),
.B2(n_1451),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1466),
.B(n_1473),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1473),
.Y(n_1597)
);

AOI222xp33_ASAP7_75t_L g1598 ( 
.A1(n_1460),
.A2(n_1431),
.B1(n_1491),
.B2(n_1457),
.C1(n_1519),
.C2(n_1489),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1519),
.A2(n_1489),
.B1(n_1445),
.B2(n_1462),
.Y(n_1599)
);

AOI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1462),
.A2(n_1487),
.B1(n_1508),
.B2(n_1550),
.C(n_1500),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1427),
.A2(n_1504),
.B1(n_1441),
.B2(n_1503),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1421),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1440),
.A2(n_1451),
.B1(n_1502),
.B2(n_1442),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1432),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1475),
.B(n_1494),
.Y(n_1605)
);

AOI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1550),
.A2(n_1500),
.B1(n_1514),
.B2(n_1497),
.C(n_1530),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1444),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1474),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1440),
.A2(n_1502),
.B1(n_1435),
.B2(n_1430),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1475),
.B(n_1495),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1497),
.A2(n_1535),
.B(n_1452),
.Y(n_1611)
);

OAI21xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1520),
.A2(n_1536),
.B(n_1496),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1420),
.A2(n_1417),
.B1(n_1471),
.B2(n_1427),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1513),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1486),
.A2(n_1471),
.B1(n_1564),
.B2(n_1523),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1523),
.A2(n_1498),
.B1(n_1452),
.B2(n_1530),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1498),
.A2(n_1514),
.B1(n_1506),
.B2(n_1436),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1436),
.A2(n_1559),
.B1(n_1555),
.B2(n_1505),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1516),
.A2(n_1561),
.B1(n_1563),
.B2(n_1566),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1513),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1509),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1501),
.B(n_1524),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1535),
.A2(n_1551),
.B(n_1573),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1529),
.A2(n_1532),
.B1(n_1537),
.B2(n_1562),
.C(n_1565),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1527),
.A2(n_1522),
.B(n_1545),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1525),
.B(n_1528),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1461),
.A2(n_1512),
.B1(n_1448),
.B2(n_1421),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1524),
.B(n_1526),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1417),
.A2(n_1419),
.B1(n_1520),
.B2(n_1521),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1421),
.A2(n_1426),
.B1(n_1461),
.B2(n_1480),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1421),
.A2(n_1426),
.B1(n_1492),
.B2(n_1480),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1531),
.B(n_1492),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1461),
.A2(n_1448),
.B1(n_1426),
.B2(n_1507),
.Y(n_1634)
);

AO31x2_ASAP7_75t_L g1635 ( 
.A1(n_1569),
.A2(n_1557),
.A3(n_1533),
.B(n_1515),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1426),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1480),
.A2(n_1536),
.B1(n_1547),
.B2(n_1552),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1552),
.A2(n_1538),
.B1(n_1543),
.B2(n_1540),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1476),
.A2(n_1516),
.B1(n_1454),
.B2(n_1459),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1557),
.B(n_1554),
.C(n_1553),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1553),
.A2(n_1573),
.B1(n_1549),
.B2(n_1568),
.C(n_1571),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1454),
.A2(n_1459),
.B1(n_1479),
.B2(n_1510),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1541),
.B(n_1542),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1490),
.A2(n_1499),
.B1(n_1510),
.B2(n_1558),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1556),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1490),
.A2(n_1534),
.B1(n_1541),
.B2(n_1539),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1483),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1546),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1517),
.A2(n_1560),
.B1(n_1568),
.B2(n_1572),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1423),
.A2(n_1549),
.B(n_1567),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1534),
.A2(n_1533),
.B1(n_1539),
.B2(n_1515),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1570),
.A2(n_1493),
.B1(n_1567),
.B2(n_1518),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_SL g1654 ( 
.A(n_1570),
.B(n_1517),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1511),
.A2(n_1544),
.B1(n_1570),
.B2(n_1493),
.C(n_1560),
.Y(n_1655)
);

AOI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1544),
.A2(n_1493),
.B(n_1570),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1483),
.A2(n_1311),
.B1(n_1428),
.B2(n_866),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1546),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1660)
);

AOI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1455),
.A2(n_1402),
.B(n_1477),
.Y(n_1661)
);

OAI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1455),
.A2(n_1467),
.B(n_1469),
.C(n_1126),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1437),
.B(n_1484),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1665)
);

OAI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1467),
.A2(n_1469),
.B(n_1126),
.C(n_1428),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1465),
.A2(n_1469),
.B(n_1311),
.C(n_412),
.Y(n_1668)
);

OA21x2_ASAP7_75t_L g1669 ( 
.A1(n_1535),
.A2(n_1316),
.B(n_1487),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1424),
.B(n_1484),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1428),
.A2(n_1280),
.B1(n_1126),
.B2(n_1311),
.C(n_1477),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1466),
.B(n_1473),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1676)
);

OAI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1467),
.A2(n_1469),
.B(n_1126),
.C(n_1428),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1482),
.A2(n_1125),
.B(n_1299),
.Y(n_1678)
);

OA21x2_ASAP7_75t_L g1679 ( 
.A1(n_1535),
.A2(n_1316),
.B(n_1487),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1481),
.B(n_1156),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1465),
.A2(n_412),
.B1(n_964),
.B2(n_742),
.C(n_1162),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_L g1682 ( 
.A1(n_1477),
.A2(n_1402),
.B(n_1469),
.Y(n_1682)
);

AO31x2_ASAP7_75t_L g1683 ( 
.A1(n_1535),
.A2(n_1316),
.A3(n_1569),
.B(n_1385),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1428),
.A2(n_1311),
.B1(n_866),
.B2(n_921),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1428),
.A2(n_1418),
.B1(n_1469),
.B2(n_866),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1469),
.A2(n_658),
.B1(n_1314),
.B2(n_1000),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1466),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1482),
.A2(n_1125),
.B(n_1299),
.Y(n_1691)
);

AOI222xp33_ASAP7_75t_L g1692 ( 
.A1(n_1465),
.A2(n_658),
.B1(n_1000),
.B2(n_409),
.C1(n_742),
.C2(n_446),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1437),
.B(n_1484),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1428),
.A2(n_1467),
.B1(n_1299),
.B2(n_1469),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1424),
.B(n_1484),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1437),
.B(n_1484),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1428),
.A2(n_1418),
.B1(n_1469),
.B2(n_866),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1424),
.Y(n_1698)
);

INVx8_ASAP7_75t_L g1699 ( 
.A(n_1461),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1428),
.A2(n_1311),
.B1(n_866),
.B2(n_921),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1428),
.A2(n_1280),
.B1(n_1126),
.B2(n_1311),
.C(n_1477),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1424),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1484),
.B(n_1424),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1604),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1659),
.B(n_1624),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1692),
.A2(n_1686),
.B1(n_1671),
.B2(n_1675),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1624),
.B(n_1683),
.Y(n_1707)
);

INVx4_ASAP7_75t_R g1708 ( 
.A(n_1690),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1612),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1607),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1624),
.B(n_1683),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1660),
.B(n_1614),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1621),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1590),
.B(n_1698),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1683),
.B(n_1611),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1608),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1648),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1683),
.B(n_1635),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1635),
.B(n_1669),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1702),
.B(n_1680),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1635),
.B(n_1669),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1651),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1622),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1574),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1635),
.B(n_1669),
.Y(n_1726)
);

CKINVDCx20_ASAP7_75t_R g1727 ( 
.A(n_1589),
.Y(n_1727)
);

NOR2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1591),
.B(n_1690),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1673),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1627),
.B(n_1640),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1650),
.B(n_1654),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1663),
.A2(n_1686),
.B1(n_1689),
.B2(n_1687),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1679),
.B(n_1653),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1592),
.B(n_1594),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1625),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1679),
.B(n_1664),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1584),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1576),
.A2(n_1682),
.B1(n_1697),
.B2(n_1688),
.C(n_1681),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1679),
.B(n_1693),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1576),
.A2(n_1701),
.B1(n_1579),
.B2(n_1694),
.C(n_1677),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1696),
.B(n_1606),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1674),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1642),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1658),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1593),
.B(n_1597),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1593),
.B(n_1620),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1596),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1652),
.B(n_1655),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1629),
.B(n_1580),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1580),
.B(n_1652),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1605),
.B(n_1610),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1619),
.B(n_1599),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1649),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1644),
.B(n_1626),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1623),
.B(n_1600),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1577),
.B(n_1586),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1657),
.B(n_1598),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1577),
.B(n_1599),
.Y(n_1759)
);

BUFx5_ASAP7_75t_L g1760 ( 
.A(n_1578),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1588),
.B(n_1601),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1619),
.B(n_1618),
.Y(n_1762)
);

OAI211xp5_ASAP7_75t_L g1763 ( 
.A1(n_1668),
.A2(n_1666),
.B(n_1700),
.C(n_1685),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1583),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1761),
.A2(n_1603),
.B1(n_1595),
.B2(n_1678),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1713),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1763),
.A2(n_1582),
.B1(n_1588),
.B2(n_1675),
.C(n_1676),
.Y(n_1767)
);

NAND4xp25_ASAP7_75t_L g1768 ( 
.A(n_1729),
.B(n_1582),
.C(n_1662),
.D(n_1670),
.Y(n_1768)
);

OAI221xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1741),
.A2(n_1676),
.B1(n_1671),
.B2(n_1684),
.C(n_1663),
.Y(n_1769)
);

AO21x2_ASAP7_75t_L g1770 ( 
.A1(n_1720),
.A2(n_1661),
.B(n_1656),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1729),
.A2(n_1687),
.B1(n_1665),
.B2(n_1667),
.C(n_1670),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1763),
.A2(n_1667),
.B1(n_1665),
.B2(n_1689),
.C(n_1684),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1587),
.C(n_1691),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1633),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1709),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1609),
.C(n_1630),
.Y(n_1776)
);

NAND4xp25_ASAP7_75t_L g1777 ( 
.A(n_1739),
.B(n_1706),
.C(n_1761),
.D(n_1732),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1706),
.A2(n_1616),
.B1(n_1613),
.B2(n_1617),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1713),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1732),
.A2(n_1616),
.B1(n_1617),
.B2(n_1618),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1754),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1709),
.B(n_1646),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1712),
.B(n_1581),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1712),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1737),
.B(n_1647),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1724),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1724),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1743),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1764),
.A2(n_1581),
.B(n_1628),
.C(n_1647),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1644),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1758),
.A2(n_1634),
.B1(n_1639),
.B2(n_1641),
.C(n_1636),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1747),
.A2(n_1631),
.B1(n_1632),
.B2(n_1646),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1740),
.B(n_1615),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1740),
.B(n_1575),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1764),
.A2(n_1637),
.B(n_1575),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1723),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1728),
.A2(n_1638),
.B(n_1602),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1721),
.B(n_1742),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1734),
.B(n_1645),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1704),
.Y(n_1803)
);

OAI211xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1721),
.A2(n_1645),
.B(n_1643),
.C(n_1699),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1705),
.B(n_1602),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1744),
.A2(n_1646),
.B1(n_1643),
.B2(n_1602),
.C(n_1699),
.Y(n_1806)
);

INVx3_ASAP7_75t_SL g1807 ( 
.A(n_1727),
.Y(n_1807)
);

NAND2xp33_ASAP7_75t_R g1808 ( 
.A(n_1718),
.B(n_1699),
.Y(n_1808)
);

OAI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1738),
.A2(n_1602),
.B(n_1646),
.C(n_1715),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1742),
.B(n_1734),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1704),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1731),
.B(n_1715),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1705),
.B(n_1750),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1710),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1753),
.A2(n_1747),
.B1(n_1759),
.B2(n_1736),
.Y(n_1815)
);

OAI33xp33_ASAP7_75t_L g1816 ( 
.A1(n_1736),
.A2(n_1730),
.A3(n_1753),
.B1(n_1744),
.B2(n_1714),
.B3(n_1734),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1715),
.B(n_1738),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1705),
.B(n_1750),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1730),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1817),
.B(n_1756),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1813),
.B(n_1760),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1813),
.B(n_1760),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1818),
.B(n_1760),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1812),
.B(n_1755),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1775),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1786),
.B(n_1775),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1807),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1776),
.A2(n_1773),
.B(n_1767),
.C(n_1785),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1756),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1807),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1782),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1775),
.B(n_1756),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1818),
.B(n_1760),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1796),
.B(n_1730),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1766),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1782),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1797),
.B(n_1760),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1760),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1780),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1785),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1810),
.B(n_1742),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1774),
.B(n_1760),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1774),
.B(n_1760),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1784),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1799),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1809),
.B(n_1760),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1801),
.B(n_1710),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1778),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1788),
.B(n_1716),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1795),
.B(n_1760),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1783),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1787),
.B(n_1746),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1784),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1788),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1789),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1795),
.B(n_1760),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1805),
.B(n_1787),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1807),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1805),
.B(n_1707),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1789),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1792),
.B(n_1707),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1803),
.B(n_1725),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1803),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1792),
.B(n_1707),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1802),
.B(n_1746),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1802),
.B(n_1717),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1812),
.B(n_1755),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1812),
.B(n_1711),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1864),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1864),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1819),
.B(n_1811),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1864),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1840),
.B(n_1815),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1837),
.B(n_1790),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1847),
.A2(n_1800),
.B(n_1816),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_SL g1877 ( 
.A(n_1827),
.B(n_1768),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1831),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1837),
.B(n_1790),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1828),
.A2(n_1815),
.B1(n_1777),
.B2(n_1768),
.C(n_1779),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1836),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1819),
.B(n_1811),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1819),
.B(n_1814),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1814),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1849),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1841),
.B(n_1798),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1837),
.B(n_1812),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1838),
.B(n_1812),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1859),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1836),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1845),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1845),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1829),
.A2(n_1773),
.B1(n_1781),
.B2(n_1779),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1838),
.B(n_1752),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1850),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1849),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1838),
.B(n_1821),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1820),
.B(n_1867),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1821),
.B(n_1752),
.Y(n_1900)
);

INVx2_ASAP7_75t_SL g1901 ( 
.A(n_1859),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1841),
.B(n_1759),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1820),
.B(n_1735),
.Y(n_1903)
);

OAI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1828),
.A2(n_1777),
.B(n_1711),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1848),
.B(n_1829),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1821),
.B(n_1752),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1867),
.B(n_1735),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1822),
.B(n_1748),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1867),
.B(n_1735),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1848),
.B(n_1759),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1832),
.B(n_1765),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1854),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1887),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1888),
.B(n_1824),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1832),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1877),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1878),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_SL g1918 ( 
.A(n_1911),
.B(n_1808),
.C(n_1847),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1907),
.B(n_1834),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1874),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1895),
.B(n_1822),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1878),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1907),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1879),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_SL g1925 ( 
.A(n_1875),
.B(n_1825),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1890),
.B(n_1827),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1895),
.B(n_1822),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1879),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1881),
.B(n_1771),
.C(n_1769),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1882),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1909),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1882),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1891),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1886),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1891),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_SL g1936 ( 
.A(n_1876),
.B(n_1830),
.C(n_1852),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1892),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1823),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1886),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1892),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1893),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1893),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1910),
.B(n_1835),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1901),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1909),
.B(n_1834),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1912),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1901),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1897),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1885),
.Y(n_1949)
);

AND4x1_ASAP7_75t_L g1950 ( 
.A(n_1888),
.B(n_1800),
.C(n_1869),
.D(n_1823),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1897),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1899),
.B(n_1834),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1900),
.B(n_1823),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1906),
.B(n_1833),
.Y(n_1954)
);

NOR3xp33_ASAP7_75t_L g1955 ( 
.A(n_1905),
.B(n_1830),
.C(n_1772),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1912),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1902),
.B(n_1835),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1920),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_SL g1959 ( 
.A(n_1950),
.B(n_1899),
.C(n_1898),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1916),
.A2(n_1929),
.B(n_1936),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1917),
.Y(n_1961)
);

AOI322xp5_ASAP7_75t_L g1962 ( 
.A1(n_1913),
.A2(n_1869),
.A3(n_1762),
.B1(n_1751),
.B2(n_1833),
.C1(n_1898),
.C2(n_1889),
.Y(n_1962)
);

OAI211xp5_ASAP7_75t_L g1963 ( 
.A1(n_1915),
.A2(n_1859),
.B(n_1852),
.C(n_1825),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1917),
.Y(n_1964)
);

OAI32xp33_ASAP7_75t_L g1965 ( 
.A1(n_1955),
.A2(n_1929),
.A3(n_1923),
.B1(n_1952),
.B2(n_1931),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1949),
.B(n_1903),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1926),
.B(n_1903),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1918),
.A2(n_1751),
.B1(n_1791),
.B2(n_1728),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1914),
.A2(n_1859),
.B1(n_1889),
.B2(n_1833),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1944),
.A2(n_1866),
.B(n_1853),
.C(n_1826),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1919),
.A2(n_1853),
.B1(n_1753),
.B2(n_1749),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1919),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1922),
.Y(n_1973)
);

O2A1O1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1947),
.A2(n_1866),
.B(n_1853),
.C(n_1826),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1947),
.B(n_1896),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1945),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1922),
.A2(n_1866),
.B(n_1869),
.C(n_1856),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1934),
.A2(n_1762),
.B1(n_1751),
.B2(n_1749),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1950),
.B(n_1872),
.Y(n_1979)
);

OAI211xp5_ASAP7_75t_L g1980 ( 
.A1(n_1925),
.A2(n_1825),
.B(n_1880),
.C(n_1875),
.Y(n_1980)
);

NAND2xp33_ASAP7_75t_SL g1981 ( 
.A(n_1952),
.B(n_1880),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1943),
.A2(n_1856),
.B(n_1872),
.Y(n_1982)
);

AOI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1924),
.A2(n_1770),
.B(n_1794),
.Y(n_1983)
);

OAI21x1_ASAP7_75t_SL g1984 ( 
.A1(n_1945),
.A2(n_1846),
.B(n_1883),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1924),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1928),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1928),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1914),
.B(n_1906),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1914),
.B(n_1908),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1957),
.B(n_1883),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1930),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1914),
.B(n_1884),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1921),
.B(n_1908),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1930),
.B(n_1858),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1968),
.A2(n_1762),
.B1(n_1733),
.B2(n_1770),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1958),
.B(n_1921),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1972),
.B(n_1927),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1972),
.B(n_1927),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1960),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1961),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1959),
.A2(n_1733),
.B1(n_1770),
.B2(n_1749),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1964),
.Y(n_2002)
);

OAI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1979),
.A2(n_1954),
.B1(n_1953),
.B2(n_1938),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1973),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1976),
.B(n_1938),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1963),
.A2(n_1953),
.B(n_1954),
.Y(n_2006)
);

NAND2x1_ASAP7_75t_L g2007 ( 
.A(n_1984),
.B(n_1932),
.Y(n_2007)
);

OAI21xp33_ASAP7_75t_L g2008 ( 
.A1(n_1965),
.A2(n_1956),
.B(n_1941),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1987),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1979),
.A2(n_1733),
.B1(n_1804),
.B2(n_1719),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1992),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1981),
.B(n_1956),
.C(n_1941),
.Y(n_2012)
);

NOR3xp33_ASAP7_75t_L g2013 ( 
.A(n_1965),
.B(n_1935),
.C(n_1942),
.Y(n_2013)
);

AOI32xp33_ASAP7_75t_L g2014 ( 
.A1(n_1981),
.A2(n_1711),
.A3(n_1757),
.B1(n_1843),
.B2(n_1844),
.Y(n_2014)
);

OAI21xp33_ASAP7_75t_SL g2015 ( 
.A1(n_1962),
.A2(n_1940),
.B(n_1937),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1985),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1976),
.B(n_1884),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1989),
.B(n_1843),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1986),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1991),
.Y(n_2020)
);

AOI21xp33_ASAP7_75t_L g2021 ( 
.A1(n_1971),
.A2(n_1951),
.B(n_1939),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1997),
.B(n_1998),
.Y(n_2022)
);

NAND3xp33_ASAP7_75t_SL g2023 ( 
.A(n_1999),
.B(n_1977),
.C(n_1980),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1996),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2019),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1999),
.B(n_1967),
.Y(n_2026)
);

OAI21xp33_ASAP7_75t_SL g2027 ( 
.A1(n_2014),
.A2(n_1988),
.B(n_1989),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2001),
.A2(n_1988),
.B1(n_1969),
.B2(n_1966),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_2016),
.B(n_2013),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2000),
.Y(n_2030)
);

XNOR2xp5_ASAP7_75t_L g2031 ( 
.A(n_2003),
.B(n_2005),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_2016),
.B(n_1975),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2002),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2004),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_L g2035 ( 
.A(n_2012),
.B(n_1974),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2015),
.A2(n_1983),
.B(n_1970),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_2013),
.A2(n_1982),
.B(n_1978),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2009),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2011),
.B(n_1993),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2020),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2017),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_2039),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2039),
.B(n_1993),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2032),
.B(n_2008),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2032),
.B(n_2006),
.Y(n_2045)
);

NAND2x1_ASAP7_75t_L g2046 ( 
.A(n_2035),
.B(n_1984),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_2041),
.B(n_2018),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2024),
.B(n_1990),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2029),
.Y(n_2049)
);

NOR2x1_ASAP7_75t_L g2050 ( 
.A(n_2023),
.B(n_2007),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_2036),
.A2(n_1995),
.B1(n_2010),
.B2(n_2021),
.Y(n_2051)
);

AOI211xp5_ASAP7_75t_L g2052 ( 
.A1(n_2023),
.A2(n_1990),
.B(n_1994),
.C(n_1935),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2025),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_2043),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_2050),
.A2(n_2037),
.B(n_2026),
.Y(n_2055)
);

O2A1O1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_2044),
.A2(n_2028),
.B(n_2038),
.C(n_2034),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2051),
.A2(n_2031),
.B1(n_2027),
.B2(n_2022),
.Y(n_2057)
);

AOI221xp5_ASAP7_75t_L g2058 ( 
.A1(n_2049),
.A2(n_2033),
.B1(n_2030),
.B2(n_2040),
.C(n_1948),
.Y(n_2058)
);

OAI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2046),
.A2(n_1946),
.B(n_1937),
.Y(n_2059)
);

AOI321xp33_ASAP7_75t_L g2060 ( 
.A1(n_2052),
.A2(n_1948),
.A3(n_1951),
.B1(n_1934),
.B2(n_1939),
.C(n_1793),
.Y(n_2060)
);

NAND4xp75_ASAP7_75t_L g2061 ( 
.A(n_2045),
.B(n_1948),
.C(n_1932),
.D(n_1946),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_2042),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_2048),
.A2(n_1942),
.B1(n_1940),
.B2(n_1933),
.C(n_1719),
.Y(n_2063)
);

OAI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2053),
.A2(n_1933),
.B(n_1839),
.C(n_1842),
.Y(n_2064)
);

O2A1O1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_2047),
.A2(n_1873),
.B(n_1871),
.C(n_1870),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2054),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2057),
.A2(n_2047),
.B1(n_1873),
.B2(n_1871),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_2062),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2055),
.B(n_1870),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_R g2070 ( 
.A(n_2056),
.B(n_1839),
.Y(n_2070)
);

OAI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_2061),
.A2(n_1844),
.B(n_1843),
.Y(n_2071)
);

NAND2xp33_ASAP7_75t_R g2072 ( 
.A(n_2059),
.B(n_2060),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2068),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_2072),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_SL g2075 ( 
.A(n_2070),
.B(n_2064),
.Y(n_2075)
);

OAI222xp33_ASAP7_75t_L g2076 ( 
.A1(n_2067),
.A2(n_2065),
.B1(n_2058),
.B2(n_2063),
.C1(n_1806),
.C2(n_1844),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_2066),
.B(n_1714),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2069),
.B(n_1858),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2071),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2078),
.Y(n_2080)
);

OR4x1_ASAP7_75t_L g2081 ( 
.A(n_2073),
.B(n_1846),
.C(n_1861),
.D(n_1854),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2074),
.A2(n_1719),
.B1(n_1726),
.B2(n_1722),
.Y(n_2082)
);

NAND4xp25_ASAP7_75t_SL g2083 ( 
.A(n_2079),
.B(n_2075),
.C(n_2076),
.D(n_2077),
.Y(n_2083)
);

NOR3xp33_ASAP7_75t_SL g2084 ( 
.A(n_2076),
.B(n_1850),
.C(n_1863),
.Y(n_2084)
);

INVxp67_ASAP7_75t_SL g2085 ( 
.A(n_2073),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2083),
.A2(n_1726),
.B1(n_1722),
.B2(n_1720),
.Y(n_2086)
);

AOI221xp5_ASAP7_75t_L g2087 ( 
.A1(n_2084),
.A2(n_1858),
.B1(n_1757),
.B2(n_1860),
.C(n_1726),
.Y(n_2087)
);

OR3x2_ASAP7_75t_L g2088 ( 
.A(n_2080),
.B(n_1708),
.C(n_1855),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2085),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_2089),
.A2(n_2088),
.B1(n_2087),
.B2(n_2086),
.Y(n_2090)
);

OA21x2_ASAP7_75t_L g2091 ( 
.A1(n_2090),
.A2(n_2082),
.B(n_2081),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2091),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2091),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2092),
.B(n_1849),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_2093),
.A2(n_1863),
.B(n_1860),
.Y(n_2095)
);

OAI222xp33_ASAP7_75t_L g2096 ( 
.A1(n_2094),
.A2(n_1860),
.B1(n_1865),
.B2(n_1862),
.C1(n_1851),
.C2(n_1857),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_R g2097 ( 
.A(n_2095),
.B(n_1842),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_SL g2098 ( 
.A1(n_2097),
.A2(n_1865),
.B1(n_1862),
.B2(n_1868),
.Y(n_2098)
);

AOI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_2098),
.A2(n_2096),
.B1(n_1855),
.B2(n_1861),
.C(n_1865),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_1851),
.B(n_1857),
.C(n_1862),
.Y(n_2100)
);


endmodule