module fake_jpeg_18367_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_21),
.B1(n_16),
.B2(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_10),
.B1(n_16),
.B2(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_2),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_27),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_17),
.B(n_19),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_31),
.B(n_20),
.C(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_21),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_36),
.B(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_25),
.C(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_14),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_36),
.B1(n_38),
.B2(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_34),
.C(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_42),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_45),
.B1(n_12),
.B2(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_12),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_9),
.Y(n_53)
);


endmodule