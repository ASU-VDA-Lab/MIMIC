module real_jpeg_3613_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx4f_ASAP7_75t_L g123 ( 
.A(n_0),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_155),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_155),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_1),
.A2(n_74),
.B1(n_75),
.B2(n_155),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_2),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_133),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_2),
.A2(n_74),
.B1(n_75),
.B2(n_133),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_64),
.B1(n_74),
.B2(n_75),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_6),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_95),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_74),
.B1(n_75),
.B2(n_95),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_7),
.A2(n_26),
.B1(n_74),
.B2(n_75),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_41),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_53),
.C(n_55),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_8),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_52),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_8),
.B(n_71),
.C(n_74),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_222),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_8),
.B(n_123),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_8),
.B(n_77),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_222),
.Y(n_287)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_20),
.B(n_345),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_12),
.B(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_13),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_87),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_87),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_13),
.A2(n_74),
.B1(n_75),
.B2(n_87),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_15),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_16),
.A2(n_27),
.B1(n_29),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_16),
.A2(n_54),
.B1(n_55),
.B2(n_187),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_16),
.A2(n_74),
.B1(n_75),
.B2(n_187),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_17),
.A2(n_40),
.B1(n_74),
.B2(n_75),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_23),
.B(n_344),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_24),
.B(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_30),
.B1(n_41),
.B2(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_27),
.A2(n_85),
.B(n_222),
.C(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_27),
.B(n_222),
.Y(n_223)
);

AOI32xp33_ASAP7_75t_L g234 ( 
.A1(n_27),
.A2(n_33),
.A3(n_35),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_30),
.A2(n_41),
.B1(n_154),
.B2(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_31),
.A2(n_63),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_31),
.A2(n_85),
.B1(n_86),
.B2(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_31),
.A2(n_94),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_31),
.B(n_132),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_31),
.A2(n_130),
.B(n_308),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_33),
.B1(n_53),
.B2(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_32),
.B(n_212),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_32),
.B(n_36),
.Y(n_236)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_340),
.B(n_342),
.Y(n_45)
);

AOI21x1_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_100),
.B(n_339),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_88),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_48),
.B(n_88),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_67),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_59),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_51),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_52),
.B(n_184),
.Y(n_288)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_55),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_55),
.B(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_61),
.B(n_65),
.C(n_67),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.C(n_84),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_80),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_93),
.C(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_77),
.B(n_78),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_69),
.A2(n_77),
.B1(n_128),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_69),
.A2(n_77),
.B1(n_149),
.B2(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_69),
.A2(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_69),
.B(n_208),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_79),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_109),
.B1(n_110),
.B2(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_73),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_73),
.A2(n_229),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_73),
.A2(n_109),
.B1(n_205),
.B2(n_255),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_74),
.B(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_77),
.B(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_83),
.B1(n_99),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_81),
.A2(n_83),
.B1(n_107),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_81),
.A2(n_83),
.B1(n_195),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_81),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_81),
.A2(n_226),
.B(n_288),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_83),
.A2(n_151),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_83),
.A2(n_183),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_153),
.B(n_156),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.C(n_96),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_89),
.A2(n_93),
.B1(n_113),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_163),
.B(n_336),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_158),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_134),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_103),
.B(n_134),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_106),
.B(n_108),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_111),
.C(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_109),
.A2(n_207),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B(n_129),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_117),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_126),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_119),
.B1(n_129),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_123),
.B(n_124),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_120),
.A2(n_123),
.B1(n_146),
.B2(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_120),
.A2(n_222),
.B(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_121),
.A2(n_122),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_121),
.A2(n_122),
.B1(n_202),
.B2(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_121),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_121),
.A2(n_122),
.B1(n_247),
.B2(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_201),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_122),
.B(n_216),
.Y(n_249)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_123),
.A2(n_215),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_150),
.C(n_152),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_143),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_144),
.A2(n_147),
.B1(n_148),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_144),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_152),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_157),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_158),
.A2(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_159),
.B(n_162),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_188),
.B(n_335),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_165),
.B(n_168),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_169),
.B(n_172),
.Y(n_333)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_174),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.C(n_185),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_175),
.A2(n_176),
.B1(n_323),
.B2(n_325),
.Y(n_322)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_177),
.B(n_179),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_178),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_185),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_186),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_330),
.B(n_334),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_299),
.B(n_327),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_241),
.B(n_298),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_217),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_217),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_203),
.C(n_209),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_193),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_197),
.C(n_200),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_203),
.B(n_209),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_231),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_218),
.B(n_232),
.C(n_240),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_230),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_219),
.B(n_225),
.C(n_227),
.Y(n_312)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_233),
.B(n_238),
.Y(n_303)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_293),
.B(n_297),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_282),
.B(n_292),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_264),
.B(n_281),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_258),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_258),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_250),
.B1(n_256),
.B2(n_257),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_253),
.C(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_275),
.B(n_280),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B(n_274),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_278),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.C(n_290),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_314),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_313),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_311),
.C(n_312),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.C(n_309),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_309),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_326),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_326),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_320),
.C(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_341),
.Y(n_344)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule