module fake_jpeg_31713_n_212 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_20),
.B(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_3),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_51),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_55),
.B(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_71),
.B1(n_75),
.B2(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_47),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_42),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_69),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_49),
.B1(n_48),
.B2(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_28),
.B1(n_16),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_28),
.B1(n_16),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_31),
.B1(n_25),
.B2(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_35),
.A2(n_31),
.B1(n_30),
.B2(n_7),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_31),
.B1(n_30),
.B2(n_7),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_39),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_37),
.B(n_5),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_107),
.Y(n_131)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_9),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_113),
.Y(n_115)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_10),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_138),
.Y(n_148)
);

NAND2x1_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_68),
.Y(n_118)
);

NOR2x1_ASAP7_75t_R g147 ( 
.A(n_118),
.B(n_68),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_52),
.B1(n_79),
.B2(n_82),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_137),
.B1(n_112),
.B2(n_134),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_59),
.B(n_63),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_128),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_59),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_135),
.C(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_70),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_67),
.C(n_58),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_86),
.B(n_80),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_134),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_80),
.B1(n_84),
.B2(n_82),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_64),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_54),
.B1(n_65),
.B2(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_92),
.B(n_54),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_125),
.C(n_115),
.Y(n_159)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_147),
.B1(n_118),
.B2(n_115),
.C(n_117),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_152),
.B1(n_156),
.B2(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_105),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_155),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_93),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_153),
.C(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_65),
.B1(n_109),
.B2(n_111),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_61),
.C(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_89),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_89),
.B1(n_72),
.B2(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_120),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_167),
.B1(n_151),
.B2(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_125),
.B1(n_118),
.B2(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_129),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.C(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_183),
.B1(n_184),
.B2(n_167),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_153),
.C(n_146),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.C(n_174),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_139),
.C(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_191),
.C(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_189),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_164),
.B1(n_166),
.B2(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_190),
.B1(n_192),
.B2(n_187),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_163),
.B(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_172),
.C(n_136),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_198),
.B(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_181),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_141),
.B(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_192),
.B1(n_172),
.B2(n_168),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_173),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_201),
.Y(n_204)
);

OAI21x1_ASAP7_75t_SL g202 ( 
.A1(n_195),
.A2(n_91),
.B(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_120),
.B1(n_102),
.B2(n_77),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_193),
.B(n_198),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_200),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_205),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_209),
.A2(n_204),
.B(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_207),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_208),
.Y(n_212)
);


endmodule