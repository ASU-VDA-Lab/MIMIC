module fake_netlist_1_9034_n_1287 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1287);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1287;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1130;
wire n_584;
wire n_1042;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVxp33_ASAP7_75t_L g298 ( .A(n_80), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_91), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_112), .B(n_286), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_91), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_105), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_238), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_17), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_63), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_62), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_11), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_174), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_248), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_167), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_231), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_138), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_55), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_276), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_186), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_166), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_78), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_148), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_58), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_125), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_214), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_77), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_75), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_66), .Y(n_327) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_57), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_281), .Y(n_329) );
INVxp33_ASAP7_75t_L g330 ( .A(n_199), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_106), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_16), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_171), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_55), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_68), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_113), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_69), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_10), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_4), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_81), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_40), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_257), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_42), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_70), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_285), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_235), .Y(n_347) );
CKINVDCx14_ASAP7_75t_R g348 ( .A(n_256), .Y(n_348) );
INVxp33_ASAP7_75t_L g349 ( .A(n_206), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_119), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_61), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_96), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_211), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_2), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_85), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_196), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_180), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_76), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_66), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_131), .Y(n_360) );
INVxp33_ASAP7_75t_SL g361 ( .A(n_46), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_289), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_170), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_215), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_234), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_3), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_160), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_213), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_27), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_219), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_51), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_156), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_73), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_152), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_128), .Y(n_375) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_263), .B(n_252), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_54), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_43), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_150), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_114), .Y(n_380) );
CKINVDCx14_ASAP7_75t_R g381 ( .A(n_129), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_258), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_197), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_179), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_168), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_87), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_230), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_90), .B(n_54), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_7), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_24), .Y(n_390) );
CKINVDCx14_ASAP7_75t_R g391 ( .A(n_279), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_108), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_217), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_278), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_96), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_42), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_188), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_134), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_21), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_117), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_120), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_222), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_153), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_264), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_247), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_76), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_124), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_47), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_216), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_49), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_6), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_246), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_20), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_239), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_274), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_205), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_0), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_251), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_270), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_269), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_275), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_39), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_204), .Y(n_423) );
INVxp33_ASAP7_75t_L g424 ( .A(n_162), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_74), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_163), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_127), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_59), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_207), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_294), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_135), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_19), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_79), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_242), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_53), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g436 ( .A(n_68), .B(n_99), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_64), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_0), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_93), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_305), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_310), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_369), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_316), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_316), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_317), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_310), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_321), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_321), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_342), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_347), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_347), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_385), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_385), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_423), .B(n_1), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_298), .B(n_1), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_412), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_412), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_335), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_317), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_344), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_415), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_357), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_348), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_318), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_308), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_357), .Y(n_466) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_318), .A2(n_103), .B(n_102), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_415), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_323), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_420), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_357), .Y(n_471) );
AND2x6_ASAP7_75t_L g472 ( .A(n_398), .B(n_104), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_323), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_334), .B(n_2), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_324), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_447), .B(n_330), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_472), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_467), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_460), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_474), .B(n_447), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_448), .B(n_349), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_472), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_460), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_448), .B(n_424), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_474), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_472), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_462), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_474), .B(n_334), .Y(n_489) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_467), .B(n_300), .Y(n_490) );
AO22x1_ASAP7_75t_L g491 ( .A1(n_472), .A2(n_315), .B1(n_361), .B2(n_331), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_449), .B(n_381), .Y(n_492) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_443), .A2(n_331), .B(n_324), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_467), .B(n_300), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_462), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_443), .B(n_423), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_467), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_449), .B(n_377), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_467), .B(n_336), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_444), .B(n_377), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_445), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_466), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_466), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_445), .B(n_343), .C(n_336), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_471), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_459), .B(n_343), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_471), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_471), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_463), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_464), .Y(n_516) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_472), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_464), .B(n_346), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_469), .B(n_407), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_469), .B(n_346), .Y(n_520) );
NAND2xp33_ASAP7_75t_L g521 ( .A(n_472), .B(n_357), .Y(n_521) );
AND2x6_ASAP7_75t_L g522 ( .A(n_473), .B(n_407), .Y(n_522) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_482), .B(n_420), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_488), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_480), .B(n_463), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_480), .B(n_455), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_480), .B(n_455), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_492), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_512), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
AND3x1_ASAP7_75t_SL g532 ( .A(n_515), .B(n_306), .C(n_301), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_492), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_480), .A2(n_442), .B1(n_454), .B2(n_361), .Y(n_535) );
INVx6_ASAP7_75t_L g536 ( .A(n_489), .Y(n_536) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_477), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_480), .B(n_473), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_485), .A2(n_486), .B1(n_498), .B2(n_489), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_476), .B(n_442), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_498), .B(n_475), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_475), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_476), .B(n_302), .Y(n_545) );
BUFx4f_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_488), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_498), .B(n_319), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_322), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_515), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_512), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_516), .A2(n_431), .B(n_394), .Y(n_552) );
BUFx8_ASAP7_75t_L g553 ( .A(n_522), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
INVx5_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_481), .B(n_302), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_488), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_516), .B(n_333), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_481), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_484), .B(n_441), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_484), .B(n_333), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_489), .B(n_319), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_477), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_516), .B(n_356), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_505), .B(n_356), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_520), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_477), .Y(n_570) );
CKINVDCx11_ASAP7_75t_R g571 ( .A(n_489), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_486), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_491), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_495), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_495), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_505), .B(n_402), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_495), .Y(n_577) );
INVx4_ASAP7_75t_L g578 ( .A(n_482), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_486), .Y(n_579) );
INVx5_ASAP7_75t_L g580 ( .A(n_519), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_501), .Y(n_581) );
AOI21x1_ASAP7_75t_L g582 ( .A1(n_491), .A2(n_431), .B(n_394), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
NOR3xp33_ASAP7_75t_SL g584 ( .A(n_509), .B(n_450), .C(n_446), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_519), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_489), .B(n_325), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_486), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_501), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_501), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_501), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_512), .Y(n_593) );
NOR3xp33_ASAP7_75t_SL g594 ( .A(n_509), .B(n_452), .C(n_451), .Y(n_594) );
NOR3xp33_ASAP7_75t_SL g595 ( .A(n_518), .B(n_456), .C(n_453), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_505), .B(n_325), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_503), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_520), .B(n_457), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_504), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_491), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_505), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_493), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_505), .B(n_327), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_506), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_506), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_511), .A2(n_378), .B(n_388), .C(n_332), .Y(n_608) );
AO22x1_ASAP7_75t_L g609 ( .A1(n_519), .A2(n_472), .B1(n_315), .B2(n_320), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_569), .Y(n_610) );
BUFx10_ASAP7_75t_L g611 ( .A(n_550), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_571), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_536), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_593), .A2(n_461), .B1(n_470), .B2(n_468), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_526), .B(n_511), .Y(n_616) );
OR2x6_ASAP7_75t_SL g617 ( .A(n_550), .B(n_465), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_598), .B(n_496), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_526), .B(n_496), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_529), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_553), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_598), .B(n_322), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_526), .B(n_519), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_603), .A2(n_490), .B(n_521), .Y(n_624) );
INVx4_ASAP7_75t_L g625 ( .A(n_571), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_536), .Y(n_626) );
BUFx8_ASAP7_75t_SL g627 ( .A(n_573), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_564), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_559), .A2(n_458), .B1(n_440), .B2(n_519), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_549), .Y(n_630) );
INVx5_ASAP7_75t_L g631 ( .A(n_554), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_553), .Y(n_632) );
INVx5_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_544), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_544), .B(n_299), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_523), .A2(n_308), .B1(n_437), .B2(n_328), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_559), .B(n_518), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_546), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_531), .A2(n_490), .B(n_521), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_595), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_527), .B(n_482), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_553), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_548), .A2(n_352), .B1(n_354), .B2(n_326), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_527), .B(n_482), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_536), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_548), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_548), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_527), .B(n_519), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_583), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_533), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_539), .A2(n_522), .B1(n_493), .B2(n_490), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_543), .B(n_522), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_531), .A2(n_490), .B(n_478), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_543), .B(n_487), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_532), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_542), .A2(n_493), .B(n_487), .Y(n_658) );
INVx4_ASAP7_75t_L g659 ( .A(n_555), .Y(n_659) );
BUFx3_ASAP7_75t_L g660 ( .A(n_546), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_560), .B(n_326), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_551), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_539), .A2(n_522), .B1(n_493), .B2(n_472), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_543), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_539), .B(n_522), .Y(n_665) );
BUFx12f_ASAP7_75t_L g666 ( .A(n_562), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_SL g667 ( .A1(n_592), .A2(n_600), .B(n_599), .C(n_567), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_535), .A2(n_522), .B1(n_354), .B2(n_493), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_562), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_599), .Y(n_670) );
INVx5_ASAP7_75t_L g671 ( .A(n_585), .Y(n_671) );
NOR2xp67_ASAP7_75t_R g672 ( .A(n_555), .B(n_487), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_584), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_602), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_540), .B(n_522), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_562), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_586), .B(n_411), .Y(n_677) );
BUFx12f_ASAP7_75t_L g678 ( .A(n_586), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_525), .A2(n_601), .B1(n_573), .B2(n_586), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_601), .A2(n_332), .B1(n_337), .B2(n_327), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_596), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_585), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_546), .A2(n_494), .B1(n_391), .B2(n_500), .Y(n_683) );
CKINVDCx8_ASAP7_75t_R g684 ( .A(n_596), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_596), .B(n_436), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_605), .B(n_522), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_605), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_605), .A2(n_494), .B1(n_500), .B2(n_497), .Y(n_688) );
AND2x6_ASAP7_75t_L g689 ( .A(n_599), .B(n_517), .Y(n_689) );
INVx4_ASAP7_75t_L g690 ( .A(n_555), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_538), .A2(n_497), .B(n_478), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_538), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_604), .B(n_307), .Y(n_693) );
BUFx3_ASAP7_75t_L g694 ( .A(n_604), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_558), .B(n_314), .Y(n_695) );
INVx3_ASAP7_75t_L g696 ( .A(n_578), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_524), .Y(n_697) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_530), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_541), .A2(n_497), .B(n_478), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_555), .B(n_517), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_524), .Y(n_701) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_600), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_568), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_534), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_580), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_545), .B(n_522), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_541), .A2(n_497), .B(n_478), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_566), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_534), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_609), .B(n_337), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_576), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_547), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_556), .B(n_338), .Y(n_713) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_530), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_561), .Y(n_715) );
CKINVDCx11_ASAP7_75t_R g716 ( .A(n_594), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_606), .B(n_338), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_572), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_572), .Y(n_719) );
CKINVDCx11_ASAP7_75t_R g720 ( .A(n_578), .Y(n_720) );
OAI21xp33_ASAP7_75t_L g721 ( .A1(n_607), .A2(n_494), .B(n_500), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_547), .B(n_339), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_579), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_580), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_579), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_608), .B(n_522), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_587), .Y(n_727) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_587), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_552), .A2(n_497), .B(n_478), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_609), .B(n_339), .Y(n_730) );
INVx1_ASAP7_75t_SL g731 ( .A(n_557), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_610), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_624), .A2(n_582), .B(n_565), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_618), .B(n_557), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_702), .A2(n_494), .B1(n_578), .B2(n_500), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_612), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_702), .A2(n_341), .B1(n_345), .B2(n_340), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_634), .B(n_565), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_630), .B(n_574), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_612), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_620), .A2(n_575), .B1(n_577), .B2(n_574), .Y(n_741) );
INVx4_ASAP7_75t_L g742 ( .A(n_720), .Y(n_742) );
AO31x2_ASAP7_75t_L g743 ( .A1(n_654), .A2(n_393), .A3(n_303), .B(n_304), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_SL g744 ( .A1(n_658), .A2(n_683), .B(n_731), .C(n_701), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_620), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_637), .A2(n_344), .B1(n_355), .B2(n_351), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_684), .A2(n_622), .B1(n_646), .B2(n_710), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_650), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_637), .A2(n_344), .B1(n_359), .B2(n_358), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_657), .A2(n_341), .B1(n_345), .B2(n_340), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_730), .A2(n_344), .B1(n_373), .B2(n_366), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_697), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_697), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_651), .B(n_371), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_619), .B(n_581), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_636), .A2(n_580), .B1(n_589), .B2(n_588), .Y(n_756) );
INVx3_ASAP7_75t_L g757 ( .A(n_662), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_661), .B(n_497), .C(n_478), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_717), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_652), .A2(n_588), .B1(n_590), .B2(n_589), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_636), .A2(n_580), .B1(n_597), .B2(n_590), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_652), .A2(n_597), .B1(n_582), .B2(n_497), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_710), .A2(n_371), .B1(n_432), .B2(n_406), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_704), .Y(n_764) );
OR2x6_ASAP7_75t_L g765 ( .A(n_666), .B(n_399), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_722), .Y(n_766) );
INVx4_ASAP7_75t_L g767 ( .A(n_720), .Y(n_767) );
AO21x2_ASAP7_75t_L g768 ( .A1(n_667), .A2(n_376), .B(n_311), .Y(n_768) );
INVx4_ASAP7_75t_L g769 ( .A(n_678), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_614), .B(n_406), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_704), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_676), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_657), .A2(n_435), .B1(n_438), .B2(n_432), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_643), .B(n_386), .Y(n_774) );
INVx4_ASAP7_75t_L g775 ( .A(n_625), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_617), .Y(n_776) );
CKINVDCx14_ASAP7_75t_R g777 ( .A(n_611), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_710), .A2(n_438), .B1(n_439), .B2(n_435), .Y(n_778) );
BUFx2_ASAP7_75t_L g779 ( .A(n_625), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_674), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_647), .A2(n_497), .B1(n_478), .B2(n_418), .Y(n_781) );
INVx4_ASAP7_75t_L g782 ( .A(n_642), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_694), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_642), .B(n_580), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_635), .Y(n_785) );
NAND3x1_ASAP7_75t_L g786 ( .A(n_629), .B(n_439), .C(n_390), .Y(n_786) );
INVx6_ASAP7_75t_L g787 ( .A(n_611), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_715), .B(n_530), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_677), .A2(n_389), .B1(n_396), .B2(n_395), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_643), .A2(n_408), .B1(n_413), .B2(n_410), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_687), .A2(n_478), .B1(n_418), .B2(n_409), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_635), .A2(n_417), .B1(n_428), .B2(n_422), .Y(n_792) );
NAND2x1_ASAP7_75t_L g793 ( .A(n_662), .B(n_591), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_703), .B(n_399), .Y(n_794) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_631), .B(n_530), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_668), .B(n_425), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_624), .A2(n_483), .B(n_479), .Y(n_797) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_694), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_640), .Y(n_799) );
AOI21xp5_ASAP7_75t_SL g800 ( .A1(n_688), .A2(n_517), .B(n_530), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_711), .B(n_425), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_682), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_685), .B(n_433), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_685), .A2(n_344), .B1(n_433), .B2(n_398), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_716), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_669), .A2(n_409), .B1(n_563), .B2(n_537), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_726), .A2(n_313), .B1(n_350), .B2(n_309), .Y(n_807) );
BUFx10_ASAP7_75t_L g808 ( .A(n_693), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_680), .A2(n_364), .B1(n_367), .B2(n_329), .C(n_312), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_681), .A2(n_563), .B1(n_570), .B2(n_537), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_621), .A2(n_401), .B1(n_404), .B2(n_379), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_664), .A2(n_360), .B1(n_362), .B2(n_353), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_680), .A2(n_363), .B1(n_368), .B2(n_365), .Y(n_813) );
OR2x6_ASAP7_75t_L g814 ( .A(n_632), .B(n_517), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_695), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_708), .B(n_537), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_709), .Y(n_817) );
AO21x2_ASAP7_75t_L g818 ( .A1(n_667), .A2(n_374), .B(n_372), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_654), .A2(n_483), .B(n_479), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_681), .A2(n_537), .B1(n_570), .B2(n_563), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_616), .A2(n_682), .B1(n_686), .B2(n_728), .Y(n_821) );
AND2x4_ASAP7_75t_L g822 ( .A(n_641), .B(n_537), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_679), .B(n_563), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_695), .A2(n_382), .B1(n_383), .B2(n_375), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_709), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g826 ( .A1(n_713), .A2(n_380), .B(n_384), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_673), .A2(n_392), .B1(n_397), .B2(n_387), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_692), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_693), .A2(n_400), .B1(n_405), .B2(n_403), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_712), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_613), .B(n_563), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_626), .B(n_570), .Y(n_832) );
AND2x4_ASAP7_75t_L g833 ( .A(n_641), .B(n_570), .Y(n_833) );
INVx4_ASAP7_75t_L g834 ( .A(n_631), .Y(n_834) );
INVx6_ASAP7_75t_L g835 ( .A(n_631), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_645), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_716), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_712), .A2(n_414), .B1(n_419), .B2(n_416), .Y(n_838) );
INVx4_ASAP7_75t_L g839 ( .A(n_631), .Y(n_839) );
AOI21xp5_ASAP7_75t_SL g840 ( .A1(n_721), .A2(n_517), .B(n_591), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_719), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_644), .B(n_4), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_675), .A2(n_591), .B1(n_517), .B2(n_421), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_718), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_623), .A2(n_591), .B1(n_517), .B2(n_426), .Y(n_845) );
INVx1_ASAP7_75t_SL g846 ( .A(n_656), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_663), .A2(n_591), .B1(n_427), .B2(n_430), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_648), .B(n_725), .Y(n_848) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_706), .A2(n_429), .B1(n_393), .B2(n_502), .C(n_499), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_627), .Y(n_850) );
NAND2x1_ASAP7_75t_L g851 ( .A(n_659), .B(n_502), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_727), .A2(n_370), .B1(n_434), .B2(n_357), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_723), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_627), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_633), .A2(n_434), .B1(n_370), .B2(n_7), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_653), .B(n_5), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_663), .A2(n_665), .B1(n_671), .B2(n_633), .Y(n_857) );
OAI21x1_ASAP7_75t_L g858 ( .A1(n_691), .A2(n_707), .B(n_699), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_633), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_628), .Y(n_860) );
BUFx10_ASAP7_75t_L g861 ( .A(n_705), .Y(n_861) );
INVx3_ASAP7_75t_L g862 ( .A(n_696), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_696), .A2(n_434), .B1(n_370), .B2(n_502), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_649), .B(n_5), .Y(n_864) );
OAI21x1_ASAP7_75t_L g865 ( .A1(n_858), .A2(n_699), .B(n_691), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_732), .Y(n_866) );
AOI21xp33_ASAP7_75t_L g867 ( .A1(n_747), .A2(n_705), .B(n_628), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_752), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_753), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_733), .A2(n_707), .B(n_729), .Y(n_870) );
OAI221xp5_ASAP7_75t_L g871 ( .A1(n_789), .A2(n_639), .B1(n_649), .B2(n_655), .C(n_615), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_785), .Y(n_872) );
INVx4_ASAP7_75t_L g873 ( .A(n_834), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_759), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g875 ( .A(n_747), .B(n_724), .C(n_700), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_804), .B(n_434), .C(n_370), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_748), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_734), .Y(n_878) );
OAI22xp33_ASAP7_75t_SL g879 ( .A1(n_776), .A2(n_671), .B1(n_633), .B2(n_670), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_765), .Y(n_880) );
AOI221x1_ASAP7_75t_SL g881 ( .A1(n_737), .A2(n_6), .B1(n_8), .B2(n_9), .C(n_10), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_763), .A2(n_670), .B1(n_671), .B2(n_698), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_770), .B(n_8), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_742), .A2(n_671), .B1(n_689), .B2(n_638), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_764), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_771), .Y(n_886) );
BUFx2_ASAP7_75t_L g887 ( .A(n_859), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_763), .A2(n_778), .B1(n_766), .B2(n_789), .Y(n_888) );
NAND2x1_ASAP7_75t_L g889 ( .A(n_834), .B(n_659), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_815), .B(n_660), .Y(n_890) );
OAI21x1_ASAP7_75t_L g891 ( .A1(n_762), .A2(n_689), .B(n_507), .Y(n_891) );
AOI211xp5_ASAP7_75t_L g892 ( .A1(n_778), .A2(n_434), .B(n_370), .C(n_499), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_750), .B(n_773), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_803), .A2(n_698), .B1(n_714), .B2(n_638), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_802), .Y(n_895) );
AOI21x1_ASAP7_75t_L g896 ( .A1(n_857), .A2(n_507), .B(n_503), .Y(n_896) );
AOI211xp5_ASAP7_75t_L g897 ( .A1(n_737), .A2(n_503), .B(n_508), .C(n_507), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_826), .A2(n_698), .B1(n_714), .B2(n_638), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_817), .Y(n_899) );
BUFx2_ASAP7_75t_L g900 ( .A(n_765), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_750), .B(n_773), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_744), .A2(n_714), .B(n_698), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_786), .A2(n_690), .B1(n_689), .B2(n_714), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_765), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_792), .A2(n_502), .B1(n_514), .B2(n_510), .C(n_508), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_802), .B(n_690), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_780), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_828), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_755), .B(n_844), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_825), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_767), .A2(n_672), .B1(n_12), .B2(n_9), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_801), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_829), .A2(n_502), .B1(n_507), .B2(n_503), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_745), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_790), .B(n_11), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_754), .B(n_12), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_813), .B(n_13), .Y(n_917) );
AOI33xp33_ASAP7_75t_L g918 ( .A1(n_827), .A2(n_514), .A3(n_510), .B1(n_508), .B2(n_16), .B3(n_17), .Y(n_918) );
NOR2x1_ASAP7_75t_L g919 ( .A(n_767), .B(n_513), .Y(n_919) );
BUFx4f_ASAP7_75t_SL g920 ( .A(n_740), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_846), .B(n_13), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_772), .Y(n_922) );
OAI21x1_ASAP7_75t_L g923 ( .A1(n_840), .A2(n_510), .B(n_508), .Y(n_923) );
OAI22xp33_ASAP7_75t_SL g924 ( .A1(n_787), .A2(n_14), .B1(n_15), .B2(n_18), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_768), .A2(n_514), .B(n_510), .Y(n_925) );
AOI322xp5_ASAP7_75t_L g926 ( .A1(n_774), .A2(n_824), .A3(n_813), .B1(n_827), .B2(n_777), .C1(n_854), .C2(n_749), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_842), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_808), .B(n_14), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_841), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_804), .A2(n_514), .B1(n_513), .B2(n_19), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_787), .A2(n_15), .B1(n_18), .B2(n_20), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_794), .A2(n_513), .B1(n_22), .B2(n_23), .C(n_24), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_746), .A2(n_513), .B1(n_22), .B2(n_23), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_808), .B(n_21), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_783), .Y(n_935) );
OAI211xp5_ASAP7_75t_L g936 ( .A1(n_811), .A2(n_513), .B(n_26), .C(n_27), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_746), .A2(n_25), .B1(n_26), .B2(n_28), .Y(n_937) );
BUFx6f_ASAP7_75t_L g938 ( .A(n_839), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_749), .A2(n_796), .B1(n_751), .B2(n_838), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_829), .A2(n_25), .B1(n_28), .B2(n_29), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_751), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_807), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_853), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_838), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_944) );
OR2x6_ASAP7_75t_L g945 ( .A(n_839), .B(n_33), .Y(n_945) );
AO21x2_ASAP7_75t_L g946 ( .A1(n_768), .A2(n_109), .B(n_107), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_855), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_775), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_782), .B(n_37), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_855), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_830), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_848), .B(n_38), .Y(n_952) );
INVx3_ASAP7_75t_L g953 ( .A(n_835), .Y(n_953) );
CKINVDCx6p67_ASAP7_75t_R g954 ( .A(n_736), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_811), .A2(n_41), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_955) );
BUFx2_ASAP7_75t_L g956 ( .A(n_769), .Y(n_956) );
INVx2_ASAP7_75t_SL g957 ( .A(n_835), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_824), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_809), .B(n_779), .Y(n_959) );
NAND3xp33_ASAP7_75t_SL g960 ( .A(n_805), .B(n_48), .C(n_50), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g961 ( .A1(n_775), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_860), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_797), .A2(n_111), .B(n_110), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_856), .A2(n_56), .B1(n_58), .B2(n_59), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_738), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_821), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_966) );
CKINVDCx9p33_ASAP7_75t_R g967 ( .A(n_850), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_800), .A2(n_116), .B(n_115), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_741), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_969) );
AO21x2_ASAP7_75t_L g970 ( .A1(n_818), .A2(n_121), .B(n_118), .Y(n_970) );
AOI322xp5_ASAP7_75t_L g971 ( .A1(n_837), .A2(n_65), .A3(n_67), .B1(n_69), .B2(n_70), .C1(n_71), .C2(n_72), .Y(n_971) );
AOI21xp33_ASAP7_75t_L g972 ( .A1(n_849), .A2(n_67), .B(n_71), .Y(n_972) );
BUFx6f_ASAP7_75t_L g973 ( .A(n_835), .Y(n_973) );
OAI211xp5_ASAP7_75t_SL g974 ( .A1(n_812), .A2(n_72), .B(n_73), .C(n_74), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_769), .B(n_78), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_739), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_783), .B(n_82), .Y(n_977) );
AOI211xp5_ASAP7_75t_L g978 ( .A1(n_799), .A2(n_83), .B(n_84), .C(n_85), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_743), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_L g980 ( .A1(n_823), .A2(n_83), .B(n_84), .C(n_86), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_798), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_981) );
OR2x2_ASAP7_75t_SL g982 ( .A(n_798), .B(n_88), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g983 ( .A1(n_756), .A2(n_89), .B1(n_92), .B2(n_93), .C(n_94), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_757), .B(n_89), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_893), .A2(n_761), .B1(n_864), .B2(n_788), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_873), .B(n_757), .Y(n_986) );
BUFx3_ASAP7_75t_L g987 ( .A(n_938), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_901), .B(n_836), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_888), .A2(n_788), .B1(n_818), .B2(n_847), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_926), .B(n_743), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_888), .A2(n_758), .B1(n_862), .B2(n_816), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_917), .A2(n_862), .B1(n_816), .B2(n_760), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_974), .A2(n_822), .B1(n_833), .B2(n_735), .Y(n_993) );
INVxp67_ASAP7_75t_L g994 ( .A(n_877), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_909), .B(n_861), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_874), .Y(n_996) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_881), .A2(n_863), .B1(n_852), .B2(n_845), .C(n_843), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_952), .A2(n_833), .B1(n_822), .B2(n_852), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_883), .B(n_743), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_866), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1001 ( .A(n_873), .B(n_743), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_952), .A2(n_861), .B1(n_863), .B2(n_781), .Y(n_1002) );
CKINVDCx11_ASAP7_75t_R g1003 ( .A(n_954), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_895), .B(n_791), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_959), .A2(n_814), .B1(n_819), .B2(n_795), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_939), .A2(n_814), .B1(n_832), .B2(n_831), .Y(n_1006) );
OA21x2_ASAP7_75t_L g1007 ( .A1(n_870), .A2(n_820), .B(n_810), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_865), .Y(n_1008) );
AOI21xp33_ASAP7_75t_L g1009 ( .A1(n_879), .A2(n_793), .B(n_814), .Y(n_1009) );
AOI21xp33_ASAP7_75t_L g1010 ( .A1(n_871), .A2(n_806), .B(n_851), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_909), .B(n_784), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_878), .B(n_92), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_927), .B(n_94), .Y(n_1013) );
BUFx2_ASAP7_75t_SL g1014 ( .A(n_949), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_938), .Y(n_1015) );
NOR2x1_ASAP7_75t_L g1016 ( .A(n_945), .B(n_95), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_939), .A2(n_95), .B1(n_97), .B2(n_98), .Y(n_1017) );
AOI211xp5_ASAP7_75t_L g1018 ( .A1(n_960), .A2(n_948), .B(n_924), .C(n_978), .Y(n_1018) );
NOR2xp33_ASAP7_75t_R g1019 ( .A(n_920), .B(n_97), .Y(n_1019) );
AOI222xp33_ASAP7_75t_L g1020 ( .A1(n_900), .A2(n_98), .B1(n_99), .B2(n_100), .C1(n_101), .C2(n_122), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_904), .B(n_100), .Y(n_1021) );
AOI211xp5_ASAP7_75t_L g1022 ( .A1(n_955), .A2(n_101), .B(n_123), .C(n_126), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_912), .A2(n_130), .B1(n_132), .B2(n_133), .C(n_136), .Y(n_1023) );
OAI211xp5_ASAP7_75t_L g1024 ( .A1(n_971), .A2(n_137), .B(n_139), .C(n_140), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_967), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_907), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_887), .B(n_297), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_977), .B(n_141), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_908), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_914), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_945), .A2(n_142), .B1(n_143), .B2(n_144), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_935), .B(n_145), .Y(n_1032) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_961), .A2(n_146), .B(n_147), .C(n_149), .Y(n_1033) );
BUFx3_ASAP7_75t_L g1034 ( .A(n_938), .Y(n_1034) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_938), .Y(n_1035) );
OAI31xp33_ASAP7_75t_L g1036 ( .A1(n_936), .A2(n_151), .A3(n_154), .B(n_155), .Y(n_1036) );
NOR2x1_ASAP7_75t_SL g1037 ( .A(n_945), .B(n_157), .Y(n_1037) );
OR2x6_ASAP7_75t_L g1038 ( .A(n_945), .B(n_158), .Y(n_1038) );
NOR2x1_ASAP7_75t_L g1039 ( .A(n_949), .B(n_159), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_892), .A2(n_161), .B1(n_164), .B2(n_165), .Y(n_1040) );
NOR4xp25_ASAP7_75t_SL g1041 ( .A(n_983), .B(n_169), .C(n_172), .D(n_173), .Y(n_1041) );
NOR2x1_ASAP7_75t_R g1042 ( .A(n_956), .B(n_175), .Y(n_1042) );
OR2x6_ASAP7_75t_L g1043 ( .A(n_873), .B(n_176), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_928), .B(n_177), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_954), .Y(n_1045) );
OAI211xp5_ASAP7_75t_L g1046 ( .A1(n_944), .A2(n_178), .B(n_181), .C(n_182), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_922), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_929), .B(n_183), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_947), .A2(n_184), .B1(n_185), .B2(n_187), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_880), .A2(n_189), .B1(n_190), .B2(n_191), .C(n_192), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_865), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_943), .B(n_193), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1053 ( .A1(n_972), .A2(n_194), .B(n_195), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_916), .B(n_198), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_872), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_947), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_950), .A2(n_203), .B1(n_208), .B2(n_209), .C(n_210), .Y(n_1057) );
INVx1_ASAP7_75t_SL g1058 ( .A(n_934), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_962), .Y(n_1059) );
AO21x2_ASAP7_75t_L g1060 ( .A1(n_925), .A2(n_212), .B(n_218), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_868), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_975), .B(n_220), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_868), .Y(n_1063) );
AOI221xp5_ASAP7_75t_SL g1064 ( .A1(n_982), .A2(n_221), .B1(n_224), .B2(n_225), .C(n_226), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_940), .A2(n_227), .B1(n_228), .B2(n_229), .C(n_232), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g1066 ( .A1(n_981), .A2(n_233), .B1(n_236), .B2(n_237), .C(n_241), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_962), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_869), .Y(n_1068) );
AO22x1_ASAP7_75t_L g1069 ( .A1(n_984), .A2(n_243), .B1(n_244), .B2(n_245), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_869), .Y(n_1070) );
AND2x4_ASAP7_75t_L g1071 ( .A(n_965), .B(n_249), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_915), .B(n_250), .Y(n_1072) );
NAND2xp5_ASAP7_75t_SL g1073 ( .A(n_918), .B(n_253), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1074 ( .A(n_980), .B(n_254), .C(n_255), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_944), .B(n_259), .Y(n_1075) );
AOI22xp5_ASAP7_75t_SL g1076 ( .A1(n_984), .A2(n_260), .B1(n_261), .B2(n_262), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_885), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_930), .A2(n_265), .B1(n_266), .B2(n_267), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_984), .Y(n_1079) );
NAND2xp33_ASAP7_75t_R g1080 ( .A(n_963), .B(n_268), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_1018), .A2(n_1017), .B1(n_1016), .B2(n_1064), .C(n_1013), .Y(n_1081) );
AO21x2_ASAP7_75t_L g1082 ( .A1(n_1008), .A2(n_925), .B(n_979), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1061), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_1001), .B(n_979), .Y(n_1084) );
INVxp67_ASAP7_75t_L g1085 ( .A(n_995), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_1038), .A2(n_966), .B1(n_930), .B2(n_882), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1059), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_1067), .Y(n_1088) );
AOI211xp5_ASAP7_75t_L g1089 ( .A1(n_1019), .A2(n_931), .B(n_911), .C(n_976), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1063), .B(n_899), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1063), .B(n_899), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1068), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1070), .B(n_886), .Y(n_1093) );
OAI22xp5_ASAP7_75t_SL g1094 ( .A1(n_1025), .A2(n_964), .B1(n_966), .B2(n_958), .Y(n_1094) );
OAI31xp33_ASAP7_75t_L g1095 ( .A1(n_1024), .A2(n_980), .A3(n_942), .B(n_969), .Y(n_1095) );
OAI31xp33_ASAP7_75t_L g1096 ( .A1(n_1013), .A2(n_958), .A3(n_876), .B(n_964), .Y(n_1096) );
INVx1_ASAP7_75t_SL g1097 ( .A(n_1003), .Y(n_1097) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_1035), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1070), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1077), .Y(n_1100) );
OAI33xp33_ASAP7_75t_L g1101 ( .A1(n_990), .A2(n_921), .A3(n_906), .B1(n_913), .B2(n_910), .B3(n_886), .Y(n_1101) );
INVx1_ASAP7_75t_SL g1102 ( .A(n_1003), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_996), .B(n_957), .Y(n_1103) );
NAND4xp25_ASAP7_75t_SL g1104 ( .A(n_1025), .B(n_937), .C(n_941), .D(n_933), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_999), .B(n_951), .Y(n_1105) );
AOI31xp67_ASAP7_75t_L g1106 ( .A1(n_1008), .A2(n_903), .A3(n_951), .B(n_910), .Y(n_1106) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_1035), .Y(n_1107) );
OAI21xp5_ASAP7_75t_SL g1108 ( .A1(n_1020), .A2(n_941), .B(n_937), .Y(n_1108) );
AOI31xp33_ASAP7_75t_L g1109 ( .A1(n_1042), .A2(n_919), .A3(n_933), .B(n_884), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1110 ( .A1(n_1017), .A2(n_932), .B1(n_890), .B2(n_875), .C(n_898), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1051), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1001), .B(n_946), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1030), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1001), .B(n_970), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1051), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1000), .B(n_973), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1026), .B(n_973), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1014), .B(n_973), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1029), .Y(n_1119) );
OAI31xp33_ASAP7_75t_L g1120 ( .A1(n_988), .A2(n_1072), .A3(n_1058), .B(n_1075), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1047), .B(n_973), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1055), .B(n_963), .Y(n_1122) );
OAI211xp5_ASAP7_75t_SL g1123 ( .A1(n_994), .A2(n_953), .B(n_894), .C(n_867), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_1038), .A2(n_894), .B1(n_963), .B2(n_968), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1079), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_992), .B(n_968), .Y(n_1126) );
INVx1_ASAP7_75t_SL g1127 ( .A(n_1045), .Y(n_1127) );
AOI21xp33_ASAP7_75t_SL g1128 ( .A1(n_1043), .A2(n_271), .B(n_272), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_992), .B(n_923), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_987), .B(n_923), .Y(n_1130) );
NOR2x1_ASAP7_75t_SL g1131 ( .A(n_1043), .B(n_896), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1007), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_987), .B(n_891), .Y(n_1133) );
OAI33xp33_ASAP7_75t_L g1134 ( .A1(n_1021), .A2(n_897), .A3(n_280), .B1(n_282), .B2(n_283), .B3(n_284), .Y(n_1134) );
AO31x2_ASAP7_75t_L g1135 ( .A1(n_1037), .A2(n_902), .A3(n_891), .B(n_889), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1015), .B(n_277), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1012), .B(n_905), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1015), .B(n_287), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1011), .B(n_288), .Y(n_1139) );
NAND4xp25_ASAP7_75t_L g1140 ( .A(n_991), .B(n_290), .C(n_291), .D(n_292), .Y(n_1140) );
HB1xp67_ASAP7_75t_SL g1141 ( .A(n_1027), .Y(n_1141) );
OAI33xp33_ASAP7_75t_L g1142 ( .A1(n_1073), .A2(n_293), .A3(n_296), .B1(n_1004), .B2(n_1078), .B3(n_1048), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_1043), .A2(n_991), .B1(n_998), .B2(n_1002), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1071), .Y(n_1144) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_1072), .A2(n_985), .B1(n_1005), .B2(n_1054), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_1034), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1062), .B(n_1044), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1071), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1084), .B(n_1071), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1113), .B(n_1005), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1119), .B(n_989), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1119), .B(n_989), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1087), .Y(n_1153) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_1088), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1105), .B(n_1034), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1116), .B(n_1006), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_1081), .A2(n_1073), .B1(n_1054), .B2(n_993), .C(n_998), .Y(n_1157) );
INVx5_ASAP7_75t_L g1158 ( .A(n_1136), .Y(n_1158) );
INVx1_ASAP7_75t_SL g1159 ( .A(n_1127), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1105), .B(n_1035), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1083), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1084), .B(n_1035), .Y(n_1162) );
NAND2x1_ASAP7_75t_L g1163 ( .A(n_1084), .B(n_1039), .Y(n_1163) );
NOR3xp33_ASAP7_75t_SL g1164 ( .A(n_1104), .B(n_1080), .C(n_1050), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1087), .B(n_1052), .Y(n_1165) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_1145), .A2(n_1080), .B1(n_1057), .B2(n_1074), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_1094), .B(n_1028), .Y(n_1167) );
NOR4xp25_ASAP7_75t_SL g1168 ( .A(n_1128), .B(n_1009), .C(n_1066), .D(n_997), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1103), .Y(n_1169) );
NAND2xp5_ASAP7_75t_SL g1170 ( .A(n_1120), .B(n_1076), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1117), .B(n_993), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1085), .B(n_986), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1125), .Y(n_1173) );
NAND4xp25_ASAP7_75t_L g1174 ( .A(n_1089), .B(n_1022), .C(n_1031), .D(n_1056), .Y(n_1174) );
AND2x2_ASAP7_75t_SL g1175 ( .A(n_1147), .B(n_986), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1121), .Y(n_1176) );
NAND4xp25_ASAP7_75t_L g1177 ( .A(n_1143), .B(n_1056), .C(n_1049), .D(n_1002), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1178 ( .A(n_1092), .B(n_986), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1092), .B(n_1032), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1100), .B(n_1069), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1100), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1129), .B(n_1060), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1129), .B(n_1049), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1146), .B(n_1010), .Y(n_1184) );
AND2x4_ASAP7_75t_L g1185 ( .A(n_1130), .B(n_1053), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1099), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1090), .B(n_1041), .Y(n_1187) );
NAND4xp25_ASAP7_75t_L g1188 ( .A(n_1108), .B(n_1036), .C(n_1065), .D(n_1023), .Y(n_1188) );
NOR3xp33_ASAP7_75t_SL g1189 ( .A(n_1140), .B(n_1046), .C(n_1033), .Y(n_1189) );
INVx2_ASAP7_75t_SL g1190 ( .A(n_1098), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1090), .B(n_1040), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_1097), .Y(n_1192) );
INVxp67_ASAP7_75t_L g1193 ( .A(n_1141), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1091), .B(n_1093), .Y(n_1194) );
INVx1_ASAP7_75t_SL g1195 ( .A(n_1102), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1091), .B(n_1093), .Y(n_1196) );
NOR3xp33_ASAP7_75t_L g1197 ( .A(n_1109), .B(n_1142), .C(n_1123), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1161), .Y(n_1198) );
AO22x1_ASAP7_75t_L g1199 ( .A1(n_1193), .A2(n_1086), .B1(n_1126), .B2(n_1112), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_1167), .A2(n_1101), .B1(n_1110), .B2(n_1134), .C(n_1096), .Y(n_1200) );
XOR2x2_ASAP7_75t_L g1201 ( .A(n_1195), .B(n_1118), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1154), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1169), .B(n_1122), .Y(n_1203) );
OAI321xp33_ASAP7_75t_L g1204 ( .A1(n_1170), .A2(n_1124), .A3(n_1112), .B1(n_1114), .B2(n_1118), .C(n_1130), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1153), .Y(n_1205) );
O2A1O1Ixp33_ASAP7_75t_L g1206 ( .A1(n_1197), .A2(n_1137), .B(n_1095), .C(n_1139), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g1207 ( .A1(n_1177), .A2(n_1148), .B1(n_1144), .B2(n_1114), .Y(n_1207) );
INVxp67_ASAP7_75t_L g1208 ( .A(n_1186), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1209 ( .A(n_1167), .B(n_1148), .Y(n_1209) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_1157), .A2(n_1144), .B1(n_1133), .B2(n_1138), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_1174), .A2(n_1133), .B1(n_1138), .B2(n_1098), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1194), .B(n_1111), .Y(n_1212) );
INVx1_ASAP7_75t_SL g1213 ( .A(n_1159), .Y(n_1213) );
NOR3xp33_ASAP7_75t_L g1214 ( .A(n_1188), .B(n_1107), .C(n_1132), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1196), .B(n_1115), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1173), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1181), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1176), .Y(n_1218) );
AOI21xp5_ASAP7_75t_L g1219 ( .A1(n_1166), .A2(n_1131), .B(n_1082), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1220 ( .A1(n_1158), .A2(n_1106), .B1(n_1135), .B2(n_1172), .Y(n_1220) );
OAI221xp5_ASAP7_75t_L g1221 ( .A1(n_1164), .A2(n_1106), .B1(n_1135), .B2(n_1150), .C(n_1192), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1186), .Y(n_1222) );
AOI221x1_ASAP7_75t_SL g1223 ( .A1(n_1151), .A2(n_1135), .B1(n_1152), .B2(n_1171), .C(n_1156), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1178), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1165), .Y(n_1225) );
AO22x1_ASAP7_75t_L g1226 ( .A1(n_1214), .A2(n_1158), .B1(n_1149), .B2(n_1185), .Y(n_1226) );
INVx1_ASAP7_75t_SL g1227 ( .A(n_1213), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_1212), .Y(n_1228) );
AOI21xp33_ASAP7_75t_L g1229 ( .A1(n_1206), .A2(n_1180), .B(n_1190), .Y(n_1229) );
XNOR2xp5_ASAP7_75t_L g1230 ( .A(n_1201), .B(n_1175), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1198), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1222), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1202), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1215), .B(n_1182), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1205), .Y(n_1235) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_1208), .B(n_1162), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1208), .Y(n_1237) );
A2O1A1Ixp33_ASAP7_75t_SL g1238 ( .A1(n_1221), .A2(n_1168), .B(n_1184), .C(n_1187), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1223), .B(n_1183), .Y(n_1239) );
NAND2xp5_ASAP7_75t_SL g1240 ( .A(n_1204), .B(n_1158), .Y(n_1240) );
XOR2x2_ASAP7_75t_L g1241 ( .A(n_1209), .B(n_1163), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1216), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1225), .B(n_1160), .Y(n_1243) );
INVx1_ASAP7_75t_SL g1244 ( .A(n_1224), .Y(n_1244) );
NAND2xp5_ASAP7_75t_SL g1245 ( .A(n_1214), .B(n_1190), .Y(n_1245) );
NOR2xp33_ASAP7_75t_R g1246 ( .A(n_1209), .B(n_1155), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1217), .Y(n_1247) );
XNOR2x1_ASAP7_75t_L g1248 ( .A(n_1199), .B(n_1179), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1218), .B(n_1182), .Y(n_1249) );
AOI31xp33_ASAP7_75t_L g1250 ( .A1(n_1230), .A2(n_1200), .A3(n_1211), .B(n_1207), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1239), .B(n_1203), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1237), .Y(n_1252) );
XNOR2x1_ASAP7_75t_L g1253 ( .A(n_1230), .B(n_1210), .Y(n_1253) );
AOI22xp5_ASAP7_75t_L g1254 ( .A1(n_1248), .A2(n_1241), .B1(n_1229), .B2(n_1245), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1231), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1232), .Y(n_1256) );
OAI31xp33_ASAP7_75t_SL g1257 ( .A1(n_1240), .A2(n_1227), .A3(n_1244), .B(n_1236), .Y(n_1257) );
INVx2_ASAP7_75t_L g1258 ( .A(n_1231), .Y(n_1258) );
NAND4xp75_ASAP7_75t_L g1259 ( .A(n_1238), .B(n_1219), .C(n_1189), .D(n_1191), .Y(n_1259) );
NOR2x1p5_ASAP7_75t_L g1260 ( .A(n_1249), .B(n_1185), .Y(n_1260) );
NAND3xp33_ASAP7_75t_L g1261 ( .A(n_1232), .B(n_1189), .C(n_1220), .Y(n_1261) );
XOR2x2_ASAP7_75t_L g1262 ( .A(n_1241), .B(n_1149), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1251), .B(n_1228), .Y(n_1263) );
BUFx8_ASAP7_75t_SL g1264 ( .A(n_1252), .Y(n_1264) );
NOR2xp33_ASAP7_75t_L g1265 ( .A(n_1253), .B(n_1243), .Y(n_1265) );
AOI21xp33_ASAP7_75t_L g1266 ( .A1(n_1250), .A2(n_1233), .B(n_1220), .Y(n_1266) );
INVx2_ASAP7_75t_SL g1267 ( .A(n_1260), .Y(n_1267) );
OAI211xp5_ASAP7_75t_L g1268 ( .A1(n_1257), .A2(n_1246), .B(n_1247), .C(n_1242), .Y(n_1268) );
NOR2x1_ASAP7_75t_SL g1269 ( .A(n_1261), .B(n_1243), .Y(n_1269) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_1254), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1262), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1256), .Y(n_1272) );
BUFx2_ASAP7_75t_L g1273 ( .A(n_1255), .Y(n_1273) );
AOI21xp33_ASAP7_75t_L g1274 ( .A1(n_1253), .A2(n_1235), .B(n_1236), .Y(n_1274) );
NOR3xp33_ASAP7_75t_L g1275 ( .A(n_1259), .B(n_1226), .C(n_1234), .Y(n_1275) );
NOR2xp67_ASAP7_75t_L g1276 ( .A(n_1258), .B(n_1254), .Y(n_1276) );
OAI21xp5_ASAP7_75t_L g1277 ( .A1(n_1270), .A2(n_1276), .B(n_1271), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1265), .B(n_1272), .Y(n_1278) );
OAI21xp5_ASAP7_75t_L g1279 ( .A1(n_1266), .A2(n_1268), .B(n_1274), .Y(n_1279) );
AND3x2_ASAP7_75t_L g1280 ( .A(n_1277), .B(n_1275), .C(n_1269), .Y(n_1280) );
XOR2xp5_ASAP7_75t_L g1281 ( .A(n_1279), .B(n_1263), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1281), .B(n_1278), .Y(n_1282) );
INVx1_ASAP7_75t_SL g1283 ( .A(n_1280), .Y(n_1283) );
BUFx2_ASAP7_75t_SL g1284 ( .A(n_1283), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1282), .Y(n_1285) );
OA22x2_ASAP7_75t_L g1286 ( .A1(n_1284), .A2(n_1267), .B1(n_1264), .B2(n_1273), .Y(n_1286) );
OR2x6_ASAP7_75t_L g1287 ( .A(n_1286), .B(n_1285), .Y(n_1287) );
endmodule