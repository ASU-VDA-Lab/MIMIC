module fake_jpeg_8035_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx6p67_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_6),
.B1(n_9),
.B2(n_8),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_18),
.B1(n_8),
.B2(n_7),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_23),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_14),
.C(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_22),
.B1(n_11),
.B2(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_25),
.C(n_26),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_27),
.B(n_26),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_37),
.B(n_33),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_32),
.B(n_25),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_34),
.C(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_29),
.A3(n_31),
.B1(n_35),
.B2(n_13),
.C1(n_12),
.C2(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_29),
.B1(n_35),
.B2(n_4),
.Y(n_43)
);


endmodule