module fake_aes_5557_n_576 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_576);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_576;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g81 ( .A(n_1), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_72), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_56), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_51), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_2), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_66), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_12), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_36), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_62), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_13), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_34), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_78), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_29), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_27), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_14), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_63), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_74), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_32), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_54), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_50), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_30), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_19), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_35), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_38), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_89), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_91), .B(n_0), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_94), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_90), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_91), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_101), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_111), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_111), .A2(n_0), .B(n_1), .Y(n_132) );
NOR2xp33_ASAP7_75t_SL g133 ( .A(n_82), .B(n_39), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_85), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_102), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_86), .B(n_3), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_86), .B(n_3), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_88), .B(n_4), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_135), .B(n_93), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_143), .Y(n_147) );
AND3x2_ASAP7_75t_L g148 ( .A(n_143), .B(n_88), .C(n_92), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_124), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_138), .B(n_120), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_129), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_138), .B(n_115), .Y(n_152) );
OR2x6_ASAP7_75t_L g153 ( .A(n_138), .B(n_92), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_138), .B(n_96), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_120), .B(n_96), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_135), .B(n_82), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_136), .B(n_116), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_120), .B(n_95), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_136), .B(n_137), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_138), .B(n_97), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_124), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_119), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_137), .B(n_95), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_156), .B(n_128), .Y(n_172) );
OR2x2_ASAP7_75t_SL g173 ( .A(n_149), .B(n_125), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_147), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_150), .B(n_132), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_147), .A2(n_125), .B1(n_84), .B2(n_132), .Y(n_177) );
AND3x1_ASAP7_75t_SL g178 ( .A(n_148), .B(n_108), .C(n_106), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_171), .B(n_134), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_167), .Y(n_180) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_155), .B(n_140), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_150), .B(n_128), .Y(n_183) );
BUFx8_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_153), .A2(n_141), .B1(n_140), .B2(n_131), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
AND2x6_ASAP7_75t_SL g188 ( .A(n_153), .B(n_141), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_155), .B(n_132), .Y(n_189) );
NOR3xp33_ASAP7_75t_SL g190 ( .A(n_158), .B(n_134), .C(n_122), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_153), .A2(n_122), .B1(n_133), .B2(n_131), .Y(n_191) );
INVxp67_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_168), .A2(n_127), .B(n_130), .C(n_121), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_146), .B(n_126), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_153), .A2(n_133), .B1(n_139), .B2(n_142), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_154), .B(n_139), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_154), .B(n_139), .Y(n_199) );
BUFx8_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_154), .B(n_126), .Y(n_201) );
BUFx2_ASAP7_75t_SL g202 ( .A(n_152), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_166), .B(n_126), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_175), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_180), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_207), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_192), .B(n_153), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_197), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g215 ( .A1(n_174), .A2(n_166), .B1(n_121), .B2(n_126), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_184), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_182), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_179), .A2(n_157), .B(n_170), .C(n_121), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_SL g220 ( .A1(n_179), .A2(n_139), .B(n_142), .C(n_121), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_181), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_185), .B(n_166), .Y(n_222) );
AOI221xp5_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_118), .B1(n_100), .B2(n_97), .C(n_112), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_172), .B(n_152), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_139), .B(n_142), .C(n_170), .Y(n_227) );
AOI33xp33_ASAP7_75t_L g228 ( .A1(n_193), .A2(n_112), .A3(n_113), .B1(n_130), .B2(n_127), .B3(n_123), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_205), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_188), .B(n_152), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_198), .A2(n_142), .B(n_121), .C(n_119), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_183), .B(n_152), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_184), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_198), .A2(n_132), .B1(n_142), .B2(n_130), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_199), .A2(n_132), .B1(n_130), .B2(n_119), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_160), .B(n_144), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_187), .B(n_99), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_199), .B(n_132), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_216), .B(n_187), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_217), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g247 ( .A1(n_223), .A2(n_113), .B1(n_190), .B2(n_119), .C(n_123), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_189), .B(n_176), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_176), .B(n_189), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
BUFx10_ASAP7_75t_L g253 ( .A(n_212), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_212), .B(n_200), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_238), .A2(n_195), .B(n_191), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_236), .A2(n_165), .B(n_161), .Y(n_256) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_160), .B(n_163), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_212), .A2(n_221), .B1(n_225), .B2(n_230), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_212), .B(n_218), .Y(n_259) );
AOI21xp33_ASAP7_75t_L g260 ( .A1(n_220), .A2(n_201), .B(n_205), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_210), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_216), .B(n_196), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_222), .A2(n_202), .B1(n_123), .B2(n_206), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_231), .A2(n_196), .B(n_206), .C(n_123), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_236), .A2(n_161), .B(n_165), .Y(n_265) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_161), .B(n_165), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_239), .A2(n_163), .B(n_145), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_233), .B(n_180), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_228), .B(n_151), .C(n_144), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_211), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_226), .A2(n_145), .B(n_87), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_210), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_244), .Y(n_273) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_268), .B(n_221), .Y(n_274) );
NAND5xp2_ASAP7_75t_SL g275 ( .A(n_247), .B(n_99), .C(n_114), .D(n_117), .E(n_173), .Y(n_275) );
AOI222xp33_ASAP7_75t_L g276 ( .A1(n_247), .A2(n_225), .B1(n_209), .B2(n_218), .C1(n_215), .C2(n_234), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_244), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_246), .B(n_213), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_268), .A2(n_233), .B1(n_242), .B2(n_214), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_268), .A2(n_233), .B1(n_200), .B2(n_213), .Y(n_280) );
BUFx12f_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_263), .A2(n_224), .B(n_232), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_249), .Y(n_283) );
AO221x2_ASAP7_75t_L g284 ( .A1(n_263), .A2(n_214), .B1(n_5), .B2(n_7), .C(n_8), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_244), .B(n_242), .Y(n_285) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_240), .B(n_242), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_250), .A2(n_226), .B(n_241), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_178), .B1(n_200), .B2(n_242), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_252), .A2(n_259), .B1(n_249), .B2(n_270), .Y(n_289) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_256), .A2(n_241), .B(n_229), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_259), .A2(n_237), .B1(n_178), .B2(n_229), .C(n_103), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_256), .A2(n_151), .B(n_210), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_252), .A2(n_235), .B1(n_210), .B2(n_117), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_255), .A2(n_114), .B(n_210), .C(n_109), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_255), .A2(n_151), .B(n_164), .C(n_7), .Y(n_295) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_256), .A2(n_151), .B(n_235), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_273), .B(n_252), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_270), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_274), .B(n_284), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_274), .B(n_251), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_284), .B(n_251), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_276), .A2(n_258), .B1(n_253), .B2(n_262), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_292), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_296), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_275), .A2(n_253), .B1(n_262), .B2(n_248), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_278), .B(n_248), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_281), .B(n_251), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_295), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_294), .B(n_265), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_296), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_298), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_305), .B(n_290), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_302), .B(n_290), .Y(n_324) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_319), .A2(n_294), .B(n_265), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_305), .B(n_265), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_302), .B(n_257), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_316), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_304), .B(n_257), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_304), .B(n_257), .Y(n_330) );
OAI33xp33_ASAP7_75t_L g331 ( .A1(n_306), .A2(n_293), .A3(n_275), .B1(n_269), .B2(n_10), .B3(n_11), .Y(n_331) );
INVx5_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_306), .B(n_257), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
INVx4_ASAP7_75t_L g336 ( .A(n_297), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_299), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_303), .A2(n_291), .B1(n_280), .B2(n_279), .C(n_288), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_311), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_299), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
AOI322xp5_ASAP7_75t_L g344 ( .A1(n_308), .A2(n_281), .A3(n_5), .B1(n_9), .B2(n_10), .C1(n_11), .C2(n_13), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_314), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_300), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
OA21x2_ASAP7_75t_L g350 ( .A1(n_310), .A2(n_287), .B(n_266), .Y(n_350) );
INVx5_ASAP7_75t_SL g351 ( .A(n_316), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_321), .B(n_323), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_346), .B(n_320), .Y(n_353) );
NOR2x1_ASAP7_75t_L g354 ( .A(n_333), .B(n_319), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_333), .B(n_313), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g356 ( .A(n_331), .B(n_307), .C(n_286), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_348), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_322), .B(n_320), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_348), .Y(n_360) );
BUFx2_ASAP7_75t_SL g361 ( .A(n_336), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_323), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_333), .B(n_301), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_322), .B(n_318), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_322), .B(n_318), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_336), .B(n_315), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_333), .B(n_301), .Y(n_369) );
NAND3xp33_ASAP7_75t_SL g370 ( .A(n_344), .B(n_312), .C(n_245), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_348), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_329), .B(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_329), .B(n_317), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_336), .B(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_342), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_346), .B(n_310), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_329), .B(n_315), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_342), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_307), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_336), .B(n_272), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_343), .Y(n_381) );
AND2x4_ASAP7_75t_SL g382 ( .A(n_336), .B(n_253), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_343), .B(n_255), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_326), .B(n_272), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_330), .B(n_271), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_4), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_332), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_330), .B(n_271), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_326), .B(n_272), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_324), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_326), .B(n_271), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_332), .B(n_14), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_347), .B(n_332), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_340), .A2(n_282), .B(n_250), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_345), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_356), .B(n_344), .C(n_340), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_379), .B(n_349), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_386), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_379), .B(n_349), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_358), .B(n_332), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_359), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_358), .B(n_334), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_372), .B(n_334), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_353), .B(n_328), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_382), .B(n_328), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_361), .B(n_364), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_362), .Y(n_410) );
NAND2x1_ASAP7_75t_SL g411 ( .A(n_354), .B(n_345), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_361), .B(n_332), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_372), .B(n_332), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_373), .B(n_332), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_363), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_387), .B(n_370), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_353), .B(n_341), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_366), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_387), .B(n_331), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_373), .B(n_332), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_382), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_354), .B(n_345), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_369), .B(n_341), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_395), .B(n_351), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_376), .B(n_324), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_366), .B(n_375), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_375), .B(n_324), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_378), .Y(n_430) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_394), .B(n_325), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_360), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_378), .B(n_327), .Y(n_433) );
INVxp33_ASAP7_75t_L g434 ( .A(n_388), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_381), .B(n_327), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_382), .B(n_351), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_392), .A2(n_327), .B(n_337), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_355), .A2(n_338), .B(n_337), .C(n_335), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_395), .B(n_351), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_384), .B(n_351), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_381), .B(n_325), .Y(n_441) );
NAND2x2_ASAP7_75t_L g442 ( .A(n_376), .B(n_351), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_377), .B(n_351), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_392), .B(n_325), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_352), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_365), .B(n_15), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g447 ( .A(n_357), .B(n_325), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_384), .B(n_350), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_365), .B(n_338), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_380), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_357), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_384), .B(n_350), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_408), .Y(n_453) );
NAND4xp25_ASAP7_75t_L g454 ( .A(n_398), .B(n_396), .C(n_367), .D(n_393), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_418), .A2(n_371), .B1(n_383), .B2(n_390), .C(n_397), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_445), .B(n_367), .Y(n_457) );
AOI22x1_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_380), .B1(n_371), .B2(n_368), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
NAND2xp33_ASAP7_75t_SL g460 ( .A(n_436), .B(n_368), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_421), .B(n_377), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_421), .B(n_390), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_407), .Y(n_463) );
A2O1A1O1Ixp25_ASAP7_75t_L g464 ( .A1(n_418), .A2(n_16), .B(n_17), .C(n_18), .D(n_19), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_405), .B(n_393), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_432), .B(n_397), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_446), .A2(n_397), .B1(n_390), .B2(n_245), .C(n_385), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_404), .B(n_385), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_410), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_442), .A2(n_397), .B1(n_390), .B2(n_368), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_446), .A2(n_391), .B1(n_384), .B2(n_389), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_413), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_400), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_425), .B(n_391), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_408), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_402), .B(n_391), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_436), .A2(n_380), .B(n_389), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_414), .B(n_368), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_409), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_399), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_432), .A2(n_380), .B(n_374), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g483 ( .A1(n_442), .A2(n_245), .B1(n_386), .B2(n_338), .C(n_335), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_401), .B(n_391), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_426), .B(n_374), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_449), .B(n_386), .Y(n_489) );
NOR4xp25_ASAP7_75t_L g490 ( .A(n_438), .B(n_337), .C(n_260), .D(n_269), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_406), .B(n_374), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_400), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_439), .A2(n_374), .B1(n_350), .B2(n_253), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_434), .A2(n_16), .B(n_17), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_450), .B(n_350), .Y(n_495) );
NOR2xp67_ASAP7_75t_SL g496 ( .A(n_443), .B(n_272), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_415), .A2(n_350), .B1(n_262), .B2(n_261), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_438), .A2(n_266), .B(n_261), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
XOR2xp5_ASAP7_75t_L g501 ( .A(n_454), .B(n_416), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_460), .A2(n_434), .B(n_411), .C(n_437), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_464), .A2(n_431), .B(n_424), .Y(n_503) );
AOI211x1_ASAP7_75t_SL g504 ( .A1(n_494), .A2(n_444), .B(n_441), .C(n_429), .Y(n_504) );
NAND2xp33_ASAP7_75t_L g505 ( .A(n_460), .B(n_422), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_476), .B(n_452), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_476), .A2(n_424), .B(n_440), .C(n_447), .Y(n_507) );
XNOR2x1_ASAP7_75t_L g508 ( .A(n_480), .B(n_419), .Y(n_508) );
AO221x1_ASAP7_75t_L g509 ( .A1(n_470), .A2(n_447), .B1(n_424), .B2(n_427), .C(n_448), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_461), .B(n_435), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_462), .A2(n_433), .B(n_260), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_453), .A2(n_261), .B1(n_262), .B2(n_235), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_469), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_462), .B(n_20), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_481), .Y(n_516) );
NOR2xp33_ASAP7_75t_SL g517 ( .A(n_458), .B(n_261), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_475), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_471), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_484), .Y(n_520) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_478), .B(n_20), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_472), .A2(n_235), .B1(n_151), .B2(n_164), .C(n_24), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
CKINVDCx14_ASAP7_75t_R g525 ( .A(n_487), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_455), .B(n_266), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_456), .A2(n_21), .B(n_22), .C(n_23), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_472), .A2(n_267), .B1(n_151), .B2(n_164), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_479), .B(n_26), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_467), .A2(n_267), .B1(n_164), .B2(n_33), .C1(n_37), .C2(n_40), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_503), .B(n_466), .C(n_488), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_516), .B(n_457), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_505), .A2(n_470), .B(n_482), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_500), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_516), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_517), .A2(n_483), .B(n_479), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_502), .A2(n_493), .B1(n_491), .B2(n_489), .C(n_486), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_517), .B(n_479), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_512), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_501), .A2(n_468), .B1(n_465), .B2(n_497), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_521), .A2(n_495), .B(n_477), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_509), .A2(n_490), .B1(n_498), .B2(n_492), .C(n_474), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g544 ( .A1(n_515), .A2(n_527), .B(n_531), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g545 ( .A1(n_513), .A2(n_496), .B(n_498), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_514), .Y(n_546) );
XOR2x2_ASAP7_75t_L g547 ( .A(n_508), .B(n_499), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_519), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_530), .A2(n_492), .B1(n_474), .B2(n_164), .C(n_44), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_523), .Y(n_550) );
OAI21xp33_ASAP7_75t_L g551 ( .A1(n_542), .A2(n_507), .B(n_511), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_541), .A2(n_506), .B1(n_510), .B2(n_524), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_534), .A2(n_525), .B(n_506), .C(n_529), .Y(n_553) );
NAND4xp25_ASAP7_75t_SL g554 ( .A(n_538), .B(n_520), .C(n_518), .D(n_522), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_532), .A2(n_528), .B1(n_526), .B2(n_504), .Y(n_555) );
AND3x2_ASAP7_75t_L g556 ( .A(n_533), .B(n_28), .C(n_31), .Y(n_556) );
OAI211xp5_ASAP7_75t_SL g557 ( .A1(n_544), .A2(n_41), .B(n_45), .C(n_46), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
OA22x2_ASAP7_75t_L g559 ( .A1(n_541), .A2(n_539), .B1(n_547), .B2(n_548), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_543), .A2(n_164), .B1(n_49), .B2(n_52), .C(n_53), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_554), .A2(n_550), .B1(n_546), .B2(n_540), .C(n_535), .Y(n_561) );
XOR2x1_ASAP7_75t_L g562 ( .A(n_558), .B(n_537), .Y(n_562) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_551), .A2(n_549), .B(n_545), .C(n_267), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_560), .B(n_48), .C(n_55), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g565 ( .A(n_552), .B(n_57), .Y(n_565) );
AND3x4_ASAP7_75t_L g566 ( .A(n_565), .B(n_559), .C(n_553), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_561), .A2(n_555), .B1(n_557), .B2(n_556), .Y(n_567) );
OA22x2_ASAP7_75t_L g568 ( .A1(n_563), .A2(n_58), .B1(n_59), .B2(n_61), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_568), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_566), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_570), .A2(n_567), .B1(n_562), .B2(n_564), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_569), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_572), .Y(n_573) );
AOI222xp33_ASAP7_75t_SL g574 ( .A1(n_573), .A2(n_571), .B1(n_65), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_574), .A2(n_64), .B1(n_70), .B2(n_71), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_575), .A2(n_73), .B1(n_76), .B2(n_77), .C(n_80), .Y(n_576) );
endmodule