module fake_jpeg_31732_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.C(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_51),
.Y(n_59)
);

NAND2x1_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_18),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_22),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_2),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_3),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_44),
.CI(n_52),
.CON(n_58),
.SN(n_58)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_68),
.B1(n_42),
.B2(n_43),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_30),
.B1(n_24),
.B2(n_33),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_38),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_82),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_8),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_62),
.C(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_40),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_67),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_90),
.B(n_61),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_88),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_67),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_66),
.B(n_68),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_83),
.B1(n_50),
.B2(n_72),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_90),
.B(n_84),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.C(n_94),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_96),
.CI(n_55),
.CON(n_102),
.SN(n_102)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_72),
.C(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_103),
.B1(n_102),
.B2(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_102),
.Y(n_106)
);


endmodule