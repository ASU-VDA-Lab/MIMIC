module fake_netlist_6_1254_n_1770 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1770);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1770;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_7),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_47),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_98),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_47),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_60),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_34),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_2),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_115),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_26),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_133),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_33),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_128),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_77),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_64),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_54),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_48),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_74),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_83),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_103),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_23),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_56),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_82),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_140),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_105),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_46),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_126),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_85),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_123),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_131),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_43),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_166),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_88),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_37),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_150),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_100),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_139),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_40),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_50),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_81),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_173),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_89),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_165),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_79),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_51),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_4),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_167),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_53),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_41),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_76),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_101),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_8),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_155),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_41),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_13),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_154),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_141),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_114),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_14),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_48),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_112),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_4),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_132),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_152),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_80),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_135),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_87),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_56),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_33),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_143),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_20),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_86),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_121),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_10),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_142),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_8),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_78),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_21),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_6),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_75),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_26),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_169),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_28),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_24),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_93),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_17),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_1),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_153),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_58),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_31),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_62),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_52),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_28),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_164),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_15),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_111),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_14),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_16),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_127),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_66),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_137),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_106),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_15),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_69),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_206),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_201),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_0),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_206),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_258),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_276),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_276),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_208),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_209),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_278),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_218),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_181),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_220),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_2),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_175),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_178),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_195),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_239),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_223),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_182),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_190),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_213),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_221),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_284),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_258),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_205),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_320),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_222),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_258),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_228),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_258),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_203),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_253),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_267),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_226),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_230),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_237),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_232),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_271),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_275),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_258),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_282),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_272),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_273),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_277),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_179),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_285),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_179),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_211),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_189),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_301),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_233),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_235),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_241),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_242),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_243),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_215),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_216),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_244),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_245),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_251),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_246),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_259),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_258),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_254),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_256),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_210),
.B(n_5),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_302),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_422),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_352),
.B(n_189),
.Y(n_437)
);

BUFx8_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_357),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_344),
.B(n_219),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_347),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_362),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_366),
.B(n_184),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

BUFx8_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_383),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_366),
.B(n_214),
.C(n_212),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

BUFx8_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_348),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_369),
.B(n_194),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_427),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_380),
.B(n_304),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_397),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_352),
.B(n_189),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_355),
.B(n_227),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_345),
.A2(n_310),
.B(n_305),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_343),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_177),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_356),
.B(n_184),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_177),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_370),
.B(n_231),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_343),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_346),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_359),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_364),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_425),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_378),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_372),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_407),
.B(n_231),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_381),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_384),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_370),
.B(n_231),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_346),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_374),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_385),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_349),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_391),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_349),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_421),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_361),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_394),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_370),
.B(n_247),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_412),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_350),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_413),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_393),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_467),
.B(n_414),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_415),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_474),
.A2(n_424),
.B1(n_429),
.B2(n_393),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_423),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_407),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_488),
.A2(n_396),
.B1(n_390),
.B2(n_387),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_443),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_371),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_475),
.B(n_483),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_463),
.B(n_176),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_458),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_398),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_442),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_457),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_454),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_475),
.B(n_371),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_426),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_465),
.B(n_176),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_445),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_477),
.B(n_426),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_501),
.B(n_388),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_503),
.B(n_430),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_371),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_452),
.B(n_176),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_492),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_459),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_431),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_445),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_446),
.A2(n_392),
.B1(n_420),
.B2(n_419),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_452),
.B(n_176),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_483),
.B(n_176),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_449),
.B(n_263),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_444),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_449),
.B(n_323),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_433),
.B(n_200),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_482),
.B(n_417),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_486),
.A2(n_494),
.B1(n_497),
.B2(n_495),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_489),
.B(n_200),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_449),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_461),
.B(n_200),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_449),
.B(n_336),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_502),
.B(n_236),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_505),
.A2(n_430),
.B1(n_234),
.B2(n_238),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_468),
.A2(n_403),
.B1(n_419),
.B2(n_411),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_451),
.B(n_489),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_489),
.B(n_200),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_432),
.B(n_392),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_468),
.B(n_200),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_466),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_466),
.B(n_202),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_432),
.B(n_395),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_470),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_433),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_451),
.B(n_250),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_451),
.B(n_250),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_473),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_473),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_451),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_436),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_476),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_480),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_480),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_464),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_435),
.B(n_395),
.Y(n_598)
);

BUFx4f_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_464),
.B(n_257),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

INVx4_ASAP7_75t_SL g602 ( 
.A(n_435),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_436),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_487),
.B(n_250),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_491),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_499),
.B(n_399),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_439),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_499),
.B(n_399),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_507),
.B(n_420),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_464),
.B(n_261),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_507),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_496),
.B(n_250),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_496),
.B(n_471),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_460),
.B(n_262),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_460),
.B(n_268),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_439),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_447),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_496),
.B(n_400),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_458),
.B(n_400),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_471),
.A2(n_409),
.B1(n_408),
.B2(n_403),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_447),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_447),
.B(n_250),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_471),
.B(n_401),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_450),
.A2(n_321),
.B1(n_291),
.B2(n_286),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_478),
.A2(n_409),
.B1(n_408),
.B2(n_406),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_450),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_450),
.B(n_283),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_453),
.B(n_287),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_453),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_434),
.B(n_315),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_453),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_456),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_500),
.B(n_186),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_479),
.B(n_411),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_479),
.A2(n_406),
.B1(n_274),
.B2(n_265),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_479),
.B(n_180),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_456),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_493),
.B(n_265),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_456),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_469),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_SL g646 ( 
.A(n_434),
.B(n_186),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_469),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_469),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_493),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_434),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_631),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_526),
.A2(n_274),
.B1(n_265),
.B2(n_258),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_631),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_586),
.Y(n_654)
);

O2A1O1Ixp5_ASAP7_75t_L g655 ( 
.A1(n_527),
.A2(n_335),
.B(n_337),
.C(n_338),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_526),
.B(n_326),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_535),
.B(n_329),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_606),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_493),
.Y(n_660)
);

CKINVDCx11_ASAP7_75t_R g661 ( 
.A(n_533),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_541),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_514),
.B(n_198),
.C(n_197),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_510),
.B(n_498),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_528),
.A2(n_199),
.B1(n_193),
.B2(n_187),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_519),
.B(n_180),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_560),
.B(n_438),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_513),
.B(n_498),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_568),
.B(n_522),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_498),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_543),
.B(n_506),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_586),
.A2(n_360),
.B(n_353),
.C(n_354),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_536),
.B(n_506),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_540),
.B(n_506),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_606),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_560),
.B(n_253),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_517),
.A2(n_295),
.B1(n_288),
.B2(n_289),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_549),
.B(n_290),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_511),
.B(n_183),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_546),
.B(n_292),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_579),
.B(n_183),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_518),
.B(n_521),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_556),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_621),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_599),
.B(n_438),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_525),
.B(n_293),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_621),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_599),
.A2(n_309),
.B1(n_294),
.B2(n_296),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_538),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_579),
.B(n_438),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_531),
.B(n_307),
.Y(n_691)
);

NAND4xp25_ASAP7_75t_SL g692 ( 
.A(n_551),
.B(n_353),
.C(n_350),
.D(n_354),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_636),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_313),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_636),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_554),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_559),
.B(n_314),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_316),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_530),
.A2(n_196),
.B1(n_185),
.B2(n_188),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_581),
.B(n_529),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_575),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_596),
.B(n_185),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_584),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_596),
.B(n_188),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_619),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_544),
.A2(n_191),
.B1(n_192),
.B2(n_279),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_589),
.B(n_265),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_572),
.B(n_187),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_544),
.A2(n_191),
.B1(n_192),
.B2(n_279),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_647),
.Y(n_710)
);

AND2x6_ASAP7_75t_SL g711 ( 
.A(n_542),
.B(n_358),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_613),
.B(n_196),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_590),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_592),
.B(n_265),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_647),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_594),
.B(n_274),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_649),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_595),
.B(n_274),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_613),
.B(n_438),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_601),
.B(n_274),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_612),
.B(n_324),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_555),
.B(n_448),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_614),
.B(n_331),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_557),
.B(n_333),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_583),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_542),
.B(n_339),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_542),
.B(n_552),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_569),
.B(n_641),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_641),
.B(n_448),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_532),
.A2(n_490),
.B1(n_484),
.B2(n_341),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_552),
.B(n_240),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_632),
.B(n_448),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_533),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_L g736 ( 
.A(n_563),
.B(n_57),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_548),
.B(n_297),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_597),
.B(n_448),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_583),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_597),
.B(n_455),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_515),
.B(n_455),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_527),
.A2(n_193),
.B1(n_199),
.B2(n_260),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_633),
.B(n_628),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_604),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_548),
.B(n_455),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_537),
.B(n_455),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_607),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_537),
.A2(n_611),
.B1(n_600),
.B2(n_617),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_610),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_545),
.B(n_358),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_622),
.B(n_248),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_537),
.B(n_249),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_578),
.A2(n_553),
.B1(n_622),
.B2(n_640),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_618),
.B(n_252),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_538),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_650),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_648),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_585),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_616),
.B(n_255),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_577),
.B(n_264),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_523),
.B(n_266),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_520),
.B(n_270),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_523),
.B(n_312),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_635),
.B(n_640),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_577),
.B(n_306),
.Y(n_767)
);

O2A1O1Ixp5_ASAP7_75t_L g768 ( 
.A1(n_578),
.A2(n_365),
.B(n_363),
.C(n_360),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_538),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_553),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_646),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_593),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_539),
.B(n_308),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_604),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_582),
.A2(n_327),
.B(n_325),
.C(n_260),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_539),
.B(n_303),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_564),
.B(n_318),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_564),
.B(n_299),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_567),
.B(n_322),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_538),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_567),
.B(n_319),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_593),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_598),
.B(n_281),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_598),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_627),
.B(n_90),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_553),
.A2(n_327),
.B1(n_325),
.B2(n_297),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_602),
.B(n_280),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_553),
.A2(n_645),
.B1(n_573),
.B2(n_562),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_509),
.B(n_70),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_624),
.B(n_11),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_561),
.B(n_73),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_573),
.A2(n_297),
.B1(n_84),
.B2(n_92),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_624),
.B(n_12),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_602),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_648),
.B(n_170),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_648),
.B(n_162),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_615),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_550),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_627),
.B(n_161),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_604),
.B(n_159),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_729),
.A2(n_574),
.B(n_634),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_684),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_728),
.B(n_629),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_762),
.B(n_629),
.C(n_605),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_654),
.B(n_512),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_654),
.B(n_512),
.Y(n_807)
);

AO22x1_ASAP7_75t_L g808 ( 
.A1(n_794),
.A2(n_558),
.B1(n_626),
.B2(n_562),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_700),
.B(n_580),
.Y(n_809)
);

AOI33xp33_ASAP7_75t_L g810 ( 
.A1(n_665),
.A2(n_642),
.A3(n_625),
.B1(n_630),
.B2(n_637),
.B3(n_620),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_667),
.B(n_605),
.C(n_615),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_701),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_660),
.A2(n_671),
.B(n_668),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_762),
.B(n_587),
.C(n_588),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_656),
.B(n_608),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_664),
.A2(n_550),
.B(n_591),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_676),
.B(n_644),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_755),
.A2(n_743),
.B(n_669),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_755),
.A2(n_588),
.B1(n_587),
.B2(n_576),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_673),
.A2(n_591),
.B(n_550),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_735),
.B(n_565),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_767),
.B(n_604),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_657),
.Y(n_823)
);

AO21x1_ASAP7_75t_L g824 ( 
.A1(n_732),
.A2(n_565),
.B(n_576),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_703),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_687),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_657),
.B(n_644),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_679),
.B(n_608),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_674),
.A2(n_591),
.B(n_550),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_743),
.A2(n_643),
.B(n_626),
.Y(n_830)
);

NAND2x1p5_ASAP7_75t_L g831 ( 
.A(n_795),
.B(n_603),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_713),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_693),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_780),
.A2(n_800),
.B(n_786),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_662),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_689),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_689),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_695),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_733),
.B(n_591),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_789),
.A2(n_608),
.B1(n_643),
.B2(n_603),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_710),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_670),
.A2(n_603),
.B(n_566),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_780),
.A2(n_566),
.B(n_524),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_768),
.A2(n_626),
.B(n_558),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_652),
.A2(n_603),
.B1(n_566),
.B2(n_524),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_732),
.A2(n_524),
.B(n_566),
.C(n_21),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_793),
.B(n_626),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_689),
.A2(n_524),
.B(n_626),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_689),
.A2(n_558),
.B(n_136),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_757),
.A2(n_558),
.B(n_124),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_652),
.A2(n_558),
.B(n_122),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_757),
.B(n_116),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_730),
.B(n_113),
.Y(n_854)
);

O2A1O1Ixp5_ASAP7_75t_L g855 ( 
.A1(n_658),
.A2(n_109),
.B(n_107),
.C(n_104),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_681),
.B(n_702),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_784),
.B(n_24),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_756),
.B(n_25),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_757),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_769),
.A2(n_799),
.B(n_682),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_737),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_769),
.B(n_799),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_SL g863 ( 
.A(n_685),
.B(n_29),
.Y(n_863)
);

AOI21xp33_ASAP7_75t_L g864 ( 
.A1(n_679),
.A2(n_29),
.B(n_30),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_770),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_801),
.A2(n_30),
.B(n_32),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_756),
.B(n_32),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_666),
.B(n_35),
.C(n_36),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_702),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_666),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_870)
);

AOI22x1_ASAP7_75t_L g871 ( 
.A1(n_715),
.A2(n_102),
.B1(n_97),
.B2(n_96),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_747),
.B(n_94),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_748),
.B(n_38),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_791),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_769),
.A2(n_45),
.B(n_52),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_769),
.A2(n_799),
.B(n_725),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_749),
.A2(n_766),
.B(n_761),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_799),
.A2(n_770),
.B(n_776),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_770),
.A2(n_782),
.B(n_773),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_651),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_763),
.A2(n_777),
.B(n_765),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_771),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_683),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_750),
.B(n_704),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_672),
.A2(n_653),
.B(n_781),
.C(n_663),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_696),
.B(n_678),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_778),
.A2(n_779),
.B(n_744),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_722),
.A2(n_704),
.B(n_712),
.C(n_727),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_744),
.A2(n_774),
.B(n_759),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_801),
.A2(n_663),
.B(n_723),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_759),
.A2(n_774),
.B(n_698),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_726),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_659),
.B(n_675),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

OAI22x1_ASAP7_75t_L g895 ( 
.A1(n_741),
.A2(n_751),
.B1(n_764),
.B2(n_745),
.Y(n_895)
);

OAI22x1_ASAP7_75t_L g896 ( 
.A1(n_690),
.A2(n_720),
.B1(n_758),
.B2(n_708),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_734),
.A2(n_680),
.B1(n_787),
.B2(n_736),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_787),
.A2(n_742),
.B1(n_798),
.B2(n_699),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_752),
.B(n_742),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_705),
.B(n_691),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_711),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_724),
.B(n_752),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_707),
.A2(n_717),
.B(n_721),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_775),
.A2(n_709),
.B(n_706),
.C(n_677),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_705),
.B(n_686),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_752),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_738),
.B(n_740),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_705),
.B(n_697),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_716),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_694),
.A2(n_797),
.B(n_796),
.Y(n_910)
);

O2A1O1Ixp5_ASAP7_75t_L g911 ( 
.A1(n_754),
.A2(n_655),
.B(n_719),
.C(n_714),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_665),
.B(n_723),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_746),
.B(n_688),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_731),
.B(n_740),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_718),
.A2(n_790),
.B(n_792),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

AOI21x1_ASAP7_75t_L g917 ( 
.A1(n_739),
.A2(n_760),
.B(n_772),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_783),
.A2(n_705),
.B(n_692),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_705),
.A2(n_729),
.B(n_645),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_701),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_729),
.A2(n_755),
.B(n_743),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_654),
.B(n_560),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_753),
.B(n_526),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_654),
.B(n_560),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_753),
.B(n_526),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_753),
.B(n_526),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_684),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_654),
.B(n_560),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_701),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_683),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_728),
.A2(n_526),
.B1(n_743),
.B2(n_669),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_753),
.B(n_526),
.Y(n_935)
);

AOI21x1_ASAP7_75t_L g936 ( 
.A1(n_660),
.A2(n_670),
.B(n_729),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_728),
.B(n_516),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_743),
.A2(n_526),
.B(n_732),
.C(n_762),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_676),
.B(n_516),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_940)
);

AO21x2_ASAP7_75t_L g941 ( 
.A1(n_789),
.A2(n_670),
.B(n_729),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_689),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_753),
.B(n_526),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_689),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_654),
.B(n_560),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_728),
.A2(n_526),
.B1(n_743),
.B2(n_669),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_700),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_753),
.B(n_526),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_654),
.B(n_560),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_743),
.A2(n_526),
.B(n_732),
.C(n_762),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_728),
.B(n_516),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_743),
.A2(n_526),
.B(n_732),
.C(n_762),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_728),
.B(n_516),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_684),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_743),
.A2(n_526),
.B(n_732),
.C(n_762),
.Y(n_960)
);

AO21x1_ASAP7_75t_L g961 ( 
.A1(n_656),
.A2(n_732),
.B(n_729),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_683),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_652),
.A2(n_656),
.B1(n_785),
.B2(n_755),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_729),
.A2(n_645),
.B(n_660),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_728),
.B(n_516),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_654),
.B(n_560),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_660),
.A2(n_670),
.B(n_729),
.Y(n_972)
);

BUFx8_ASAP7_75t_L g973 ( 
.A(n_771),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_689),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_834),
.A2(n_822),
.B(n_919),
.Y(n_975)
);

AO31x2_ASAP7_75t_L g976 ( 
.A1(n_961),
.A2(n_824),
.A3(n_960),
.B(n_938),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_905),
.B(n_900),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_925),
.B(n_928),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_935),
.B(n_943),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_836),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_948),
.A2(n_946),
.B1(n_934),
.B2(n_923),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_882),
.Y(n_982)
);

AO31x2_ASAP7_75t_L g983 ( 
.A1(n_890),
.A2(n_968),
.A3(n_819),
.B(n_846),
.Y(n_983)
);

INVx8_ASAP7_75t_L g984 ( 
.A(n_836),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_923),
.A2(n_818),
.B(n_877),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_812),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_818),
.A2(n_877),
.B(n_968),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_856),
.A2(n_912),
.B(n_888),
.C(n_857),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_924),
.B(n_926),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_931),
.B(n_945),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_836),
.Y(n_992)
);

OAI22xp33_ASAP7_75t_L g993 ( 
.A1(n_898),
.A2(n_869),
.B1(n_858),
.B2(n_867),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_887),
.A2(n_878),
.B(n_876),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_950),
.B(n_971),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_842),
.A2(n_913),
.B(n_936),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_908),
.A2(n_815),
.B(n_910),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_820),
.A2(n_829),
.B(n_915),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_920),
.A2(n_958),
.B(n_957),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_880),
.B(n_906),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_939),
.B(n_886),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_922),
.A2(n_949),
.B(n_962),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_816),
.A2(n_889),
.B(n_879),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_827),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_SL g1005 ( 
.A1(n_866),
.A2(n_852),
.B(n_885),
.Y(n_1005)
);

OAI22x1_ASAP7_75t_L g1006 ( 
.A1(n_899),
.A2(n_914),
.B1(n_952),
.B2(n_970),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_803),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_903),
.A2(n_860),
.B(n_881),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_927),
.A2(n_954),
.B(n_965),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_823),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_804),
.A2(n_897),
.B1(n_904),
.B2(n_940),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_959),
.A2(n_969),
.B(n_966),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_825),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_883),
.B(n_937),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_837),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_809),
.B(n_817),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_963),
.A2(n_964),
.B(n_805),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_955),
.A2(n_947),
.B(n_902),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_941),
.A2(n_884),
.B1(n_852),
.B2(n_828),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_911),
.A2(n_802),
.B(n_840),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_832),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_SL g1022 ( 
.A(n_864),
.B(n_865),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_802),
.A2(n_862),
.B(n_843),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_830),
.A2(n_972),
.B(n_814),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_SL g1025 ( 
.A1(n_941),
.A2(n_907),
.B(n_845),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_863),
.A2(n_932),
.B1(n_921),
.B2(n_841),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_837),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_SL g1028 ( 
.A1(n_907),
.A2(n_830),
.B(n_854),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_861),
.B(n_839),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_806),
.B(n_807),
.Y(n_1030)
);

NAND2x1_ASAP7_75t_L g1031 ( 
.A(n_851),
.B(n_944),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_SL g1032 ( 
.A1(n_875),
.A2(n_874),
.B(n_871),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_803),
.B(n_930),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_808),
.A2(n_872),
.B(n_893),
.Y(n_1034)
);

AO31x2_ASAP7_75t_L g1035 ( 
.A1(n_895),
.A2(n_870),
.A3(n_896),
.B(n_874),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_855),
.A2(n_810),
.B(n_844),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_848),
.A2(n_831),
.B(n_844),
.Y(n_1037)
);

AOI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_835),
.A2(n_826),
.B(n_833),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_930),
.B(n_956),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_865),
.A2(n_944),
.B(n_942),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_956),
.B(n_838),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_837),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_851),
.A2(n_859),
.A3(n_942),
.B(n_849),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_865),
.A2(n_974),
.B1(n_859),
.B2(n_909),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_811),
.A2(n_847),
.B(n_868),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_974),
.A2(n_909),
.B(n_853),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_831),
.A2(n_853),
.B(n_850),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_873),
.A2(n_909),
.B(n_847),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_974),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_933),
.B(n_821),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_909),
.A2(n_821),
.B(n_916),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_916),
.B(n_821),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_967),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_847),
.B(n_901),
.Y(n_1054)
);

AO21x1_ASAP7_75t_L g1055 ( 
.A1(n_847),
.A2(n_882),
.B(n_973),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_894),
.Y(n_1056)
);

AOI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_856),
.A2(n_928),
.B(n_925),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_939),
.B(n_924),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_836),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_834),
.A2(n_822),
.B(n_919),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_834),
.A2(n_822),
.B(n_919),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_880),
.B(n_906),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_938),
.A2(n_953),
.B(n_951),
.Y(n_1063)
);

INVx8_ASAP7_75t_L g1064 ( 
.A(n_836),
.Y(n_1064)
);

AO31x2_ASAP7_75t_L g1065 ( 
.A1(n_961),
.A2(n_824),
.A3(n_953),
.B(n_951),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_892),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_SL g1067 ( 
.A(n_895),
.B(n_733),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_925),
.A2(n_929),
.B(n_928),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_835),
.B(n_700),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_834),
.A2(n_822),
.B(n_919),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_SL g1071 ( 
.A(n_894),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_938),
.A2(n_953),
.B(n_951),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_892),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_928),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_866),
.A2(n_890),
.B(n_918),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_939),
.B(n_924),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_812),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1078)
);

INVx6_ASAP7_75t_SL g1079 ( 
.A(n_821),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_834),
.A2(n_822),
.B(n_919),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_938),
.A2(n_953),
.B(n_951),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_836),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_925),
.A2(n_928),
.B1(n_935),
.B2(n_929),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_925),
.B(n_928),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_961),
.A2(n_824),
.A3(n_953),
.B(n_951),
.Y(n_1087)
);

INVx5_ASAP7_75t_L g1088 ( 
.A(n_836),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_835),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_836),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_835),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_933),
.B(n_735),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_836),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_938),
.A2(n_953),
.B(n_951),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_835),
.B(n_700),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_939),
.B(n_924),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_925),
.B(n_928),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_938),
.A2(n_953),
.B1(n_960),
.B2(n_951),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_939),
.B(n_924),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_925),
.B(n_928),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_836),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_812),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_938),
.A2(n_953),
.B(n_960),
.C(n_951),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_939),
.B(n_924),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_938),
.B(n_953),
.C(n_951),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_883),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_856),
.A2(n_635),
.B1(n_571),
.B2(n_912),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_967),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_925),
.A2(n_928),
.B1(n_935),
.B2(n_929),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_938),
.A2(n_953),
.B(n_951),
.Y(n_1113)
);

NAND2x1_ASAP7_75t_L g1114 ( 
.A(n_851),
.B(n_859),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_917),
.A2(n_918),
.B(n_891),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_925),
.B(n_928),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_961),
.A2(n_824),
.A3(n_953),
.B(n_951),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_856),
.A2(n_928),
.B(n_925),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_988),
.A2(n_1118),
.B(n_1057),
.C(n_989),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1089),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1058),
.B(n_1076),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1110),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_982),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1092),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1010),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1108),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1004),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1097),
.B(n_1100),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1000),
.B(n_1062),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_990),
.B(n_995),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1013),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1071),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1062),
.B(n_1050),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_977),
.A2(n_997),
.B(n_1081),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_984),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1021),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1106),
.B(n_978),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1077),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1014),
.B(n_1052),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1063),
.A2(n_1095),
.B(n_1072),
.C(n_1113),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_984),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1104),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1007),
.B(n_1029),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_975),
.A2(n_1060),
.B(n_1061),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_984),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_1064),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1109),
.A2(n_981),
.B1(n_1107),
.B2(n_1006),
.Y(n_1148)
);

INVx4_ASAP7_75t_L g1149 ( 
.A(n_1059),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_979),
.B(n_1074),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1093),
.Y(n_1152)
);

OR2x6_ASAP7_75t_L g1153 ( 
.A(n_1064),
.B(n_1093),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1064),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1001),
.B(n_1086),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1079),
.Y(n_1156)
);

AOI221x1_ASAP7_75t_L g1157 ( 
.A1(n_1105),
.A2(n_1107),
.B1(n_1011),
.B2(n_987),
.C(n_1005),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_1055),
.A2(n_1075),
.B(n_1045),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1056),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_987),
.A2(n_985),
.B(n_1024),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1071),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_992),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1098),
.B(n_1101),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1066),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_985),
.A2(n_1116),
.B1(n_993),
.B2(n_1054),
.C1(n_1067),
.C2(n_1045),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1051),
.B(n_1073),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_1030),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_SL g1169 ( 
.A(n_1044),
.B(n_1059),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1068),
.B(n_1019),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_1026),
.B(n_1017),
.C(n_1038),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1079),
.A2(n_1016),
.B1(n_1028),
.B2(n_1025),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1070),
.A2(n_1080),
.B(n_1012),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1022),
.A2(n_1041),
.B1(n_1033),
.B2(n_1039),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1049),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1027),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_991),
.A2(n_1078),
.B(n_1115),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_992),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1036),
.A2(n_1059),
.B1(n_1088),
.B2(n_1046),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1032),
.A2(n_1022),
.B1(n_1053),
.B2(n_1024),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_983),
.B(n_976),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1088),
.B(n_1094),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1088),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1090),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_999),
.A2(n_1002),
.B(n_1009),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_992),
.B(n_1042),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1009),
.A2(n_1008),
.B(n_994),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1035),
.B(n_1103),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1015),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1048),
.A2(n_1020),
.B(n_1047),
.C(n_1023),
.Y(n_1190)
);

OR2x6_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_1042),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1103),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_983),
.B(n_976),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1015),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1035),
.B(n_976),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1042),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1035),
.B(n_1065),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_980),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1034),
.A2(n_980),
.B1(n_1084),
.B2(n_1094),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_998),
.A2(n_1003),
.B(n_1091),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1065),
.B(n_1117),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1084),
.A2(n_1040),
.B1(n_1114),
.B2(n_1031),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1037),
.B(n_1083),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_983),
.A2(n_996),
.B1(n_1087),
.B2(n_1117),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1082),
.B(n_1102),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1111),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1087),
.B(n_1043),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1043),
.B(n_1058),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1000),
.B(n_1062),
.Y(n_1209)
);

BUFx10_ASAP7_75t_L g1210 ( 
.A(n_1071),
.Y(n_1210)
);

AOI21xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1069),
.A2(n_741),
.B(n_458),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_984),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_988),
.B(n_938),
.Y(n_1213)
);

NAND2xp33_ASAP7_75t_L g1214 ( 
.A(n_988),
.B(n_938),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1109),
.A2(n_856),
.B1(n_912),
.B2(n_898),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_977),
.A2(n_997),
.B(n_834),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1108),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1108),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1109),
.A2(n_928),
.B1(n_929),
.B2(n_925),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_984),
.B(n_1064),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1000),
.B(n_1062),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1058),
.B(n_1076),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_992),
.Y(n_1225)
);

OAI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_989),
.A2(n_856),
.B(n_990),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_984),
.B(n_1064),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1059),
.B(n_1088),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1069),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1109),
.B(n_856),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_984),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1058),
.B(n_1076),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1081),
.A2(n_997),
.B(n_977),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_992),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_989),
.B(n_856),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1081),
.A2(n_997),
.B(n_977),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_986),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1069),
.B(n_1096),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1109),
.B(n_856),
.Y(n_1239)
);

NOR2x1_ASAP7_75t_SL g1240 ( 
.A(n_1044),
.B(n_865),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1024),
.A2(n_1020),
.B(n_1017),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1053),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1058),
.B(n_1076),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_984),
.B(n_1064),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_984),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_SL g1247 ( 
.A(n_1079),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1000),
.B(n_1062),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1058),
.B(n_1076),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_986),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_988),
.B(n_856),
.C(n_938),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_986),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1069),
.B(n_1096),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_984),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_986),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_991),
.A2(n_1082),
.B(n_1078),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_1122),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1138),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1124),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1230),
.A2(n_1239),
.B1(n_1235),
.B2(n_1215),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1155),
.B(n_1163),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1208),
.B(n_1219),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1123),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1120),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1217),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1200),
.A2(n_1187),
.B(n_1233),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1142),
.Y(n_1268)
);

INVxp67_ASAP7_75t_SL g1269 ( 
.A(n_1127),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1237),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1255),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1131),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1141),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1133),
.B(n_1139),
.Y(n_1274)
);

AOI222xp33_ASAP7_75t_L g1275 ( 
.A1(n_1213),
.A2(n_1214),
.B1(n_1226),
.B2(n_1130),
.C1(n_1251),
.C2(n_1137),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1141),
.Y(n_1276)
);

BUFx8_ASAP7_75t_SL g1277 ( 
.A(n_1132),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1238),
.Y(n_1279)
);

BUFx2_ASAP7_75t_R g1280 ( 
.A(n_1161),
.Y(n_1280)
);

AND2x4_ASAP7_75t_SL g1281 ( 
.A(n_1221),
.B(n_1227),
.Y(n_1281)
);

BUFx8_ASAP7_75t_SL g1282 ( 
.A(n_1156),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1177),
.A2(n_1256),
.B(n_1216),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1228),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1168),
.A2(n_1151),
.B1(n_1139),
.B2(n_1133),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1253),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1250),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1251),
.A2(n_1257),
.B1(n_1150),
.B2(n_1245),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1252),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1188),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1165),
.A2(n_1148),
.B1(n_1226),
.B2(n_1257),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1144),
.A2(n_1245),
.B1(n_1220),
.B2(n_1150),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1164),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1219),
.B(n_1144),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1229),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1165),
.A2(n_1220),
.B1(n_1222),
.B2(n_1249),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1141),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1175),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1146),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1125),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1222),
.A2(n_1224),
.B1(n_1121),
.B2(n_1232),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1242),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1243),
.A2(n_1167),
.B1(n_1151),
.B2(n_1223),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1241),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1180),
.A2(n_1128),
.B1(n_1171),
.B2(n_1158),
.Y(n_1305)
);

BUFx8_ASAP7_75t_L g1306 ( 
.A(n_1126),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1140),
.B(n_1160),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1143),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_SL g1309 ( 
.A(n_1210),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1203),
.Y(n_1310)
);

AO21x1_ASAP7_75t_L g1311 ( 
.A1(n_1119),
.A2(n_1170),
.B(n_1204),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1207),
.B(n_1166),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1176),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1203),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1172),
.A2(n_1171),
.B1(n_1152),
.B2(n_1211),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1129),
.A2(n_1209),
.B1(n_1248),
.B2(n_1223),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1203),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1228),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1134),
.A2(n_1173),
.B(n_1236),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1157),
.A2(n_1185),
.B(n_1173),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1153),
.B(n_1129),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1184),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1192),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1196),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1195),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1206),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1210),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1201),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1153),
.A2(n_1174),
.B1(n_1172),
.B2(n_1159),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1197),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1198),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1160),
.B(n_1174),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1186),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1170),
.B(n_1193),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1181),
.B(n_1193),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1218),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_SL g1337 ( 
.A(n_1189),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1186),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1153),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1247),
.A2(n_1169),
.B1(n_1179),
.B2(n_1240),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1186),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1233),
.A2(n_1236),
.B(n_1145),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1191),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1205),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1221),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1162),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1191),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1179),
.A2(n_1199),
.B1(n_1147),
.B2(n_1246),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1190),
.A2(n_1199),
.B(n_1202),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1191),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1162),
.B(n_1234),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1162),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1135),
.A2(n_1254),
.B1(n_1231),
.B2(n_1154),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1202),
.A2(n_1182),
.B(n_1227),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1178),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1182),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1178),
.B(n_1225),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1147),
.A2(n_1246),
.B1(n_1212),
.B2(n_1149),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1135),
.A2(n_1254),
.B(n_1154),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1212),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1225),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1231),
.A2(n_1183),
.B1(n_1244),
.B2(n_1227),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1194),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1244),
.B(n_1225),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1244),
.A2(n_1149),
.B(n_1212),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1234),
.B(n_1246),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_1187),
.B(n_1099),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1235),
.A2(n_635),
.B1(n_856),
.B2(n_571),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1230),
.A2(n_1239),
.B1(n_1215),
.B2(n_1109),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1230),
.A2(n_1239),
.B1(n_1215),
.B2(n_1109),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1155),
.B(n_1215),
.Y(n_1371)
);

AND2x2_ASAP7_75t_SL g1372 ( 
.A(n_1215),
.B(n_1213),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1155),
.B(n_1215),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1238),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_1267),
.B(n_1367),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1328),
.B(n_1332),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1304),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1292),
.B(n_1288),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1310),
.B(n_1317),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1320),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1320),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1344),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1334),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1320),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1334),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1339),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1307),
.B(n_1330),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1319),
.A2(n_1283),
.B(n_1354),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1314),
.B(n_1354),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1325),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1326),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1326),
.Y(n_1392)
);

AO21x1_ASAP7_75t_SL g1393 ( 
.A1(n_1291),
.A2(n_1370),
.B(n_1369),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1311),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1335),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1335),
.B(n_1330),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1312),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1307),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1294),
.B(n_1275),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1349),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1294),
.A2(n_1263),
.B(n_1305),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1339),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1263),
.B(n_1290),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1290),
.B(n_1329),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1296),
.B(n_1371),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1261),
.A2(n_1289),
.B(n_1287),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1272),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1278),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1269),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1359),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1303),
.B(n_1286),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1371),
.A2(n_1373),
.B(n_1298),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1373),
.B(n_1301),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1331),
.A2(n_1333),
.B(n_1350),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1279),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1372),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1374),
.B(n_1285),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1313),
.A2(n_1322),
.B(n_1323),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1259),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1268),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1270),
.Y(n_1421)
);

OAI21xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1372),
.A2(n_1262),
.B(n_1271),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1276),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1365),
.B(n_1308),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1260),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1262),
.B(n_1315),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1293),
.A2(n_1338),
.B(n_1341),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1295),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1348),
.Y(n_1429)
);

BUFx4f_ASAP7_75t_SL g1430 ( 
.A(n_1302),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1343),
.A2(n_1324),
.B(n_1362),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1274),
.B(n_1321),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1274),
.B(n_1321),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1281),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1274),
.B(n_1355),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1340),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1395),
.B(n_1412),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1412),
.B(n_1265),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1383),
.B(n_1368),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1427),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1375),
.A2(n_1361),
.B(n_1347),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_1364),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1412),
.B(n_1357),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1410),
.B(n_1281),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1385),
.B(n_1300),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1398),
.B(n_1351),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1398),
.B(n_1351),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1408),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1388),
.A2(n_1318),
.B(n_1364),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1382),
.B(n_1284),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1427),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1387),
.B(n_1352),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1387),
.B(n_1352),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1389),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1386),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1406),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1406),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1376),
.B(n_1377),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1399),
.B(n_1345),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1380),
.B(n_1346),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1396),
.B(n_1356),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1396),
.B(n_1318),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1396),
.B(n_1318),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1418),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1418),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1436),
.B(n_1345),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1284),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1418),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1400),
.B(n_1284),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1389),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1381),
.B(n_1366),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1436),
.B(n_1316),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1400),
.B(n_1353),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1381),
.B(n_1336),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1389),
.Y(n_1475)
);

AOI222xp33_ASAP7_75t_L g1476 ( 
.A1(n_1378),
.A2(n_1309),
.B1(n_1302),
.B2(n_1327),
.C1(n_1306),
.C2(n_1266),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1418),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1384),
.B(n_1363),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1476),
.A2(n_1378),
.B(n_1459),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1438),
.B(n_1411),
.Y(n_1481)
);

NOR3xp33_ASAP7_75t_L g1482 ( 
.A(n_1459),
.B(n_1429),
.C(n_1405),
.Y(n_1482)
);

OAI221xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1476),
.A2(n_1429),
.B1(n_1417),
.B2(n_1405),
.C(n_1422),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1446),
.B(n_1425),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1472),
.A2(n_1417),
.B1(n_1411),
.B2(n_1415),
.C(n_1422),
.Y(n_1485)
);

NAND4xp25_ASAP7_75t_L g1486 ( 
.A(n_1439),
.B(n_1472),
.C(n_1445),
.D(n_1466),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1439),
.B(n_1411),
.C(n_1416),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1466),
.A2(n_1416),
.B1(n_1404),
.B2(n_1426),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1445),
.A2(n_1416),
.B1(n_1404),
.B2(n_1426),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1452),
.A2(n_1416),
.B1(n_1404),
.B2(n_1426),
.Y(n_1490)
);

OAI221xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1438),
.A2(n_1413),
.B1(n_1394),
.B2(n_1415),
.C(n_1393),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_SL g1493 ( 
.A(n_1455),
.B(n_1280),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1438),
.B(n_1416),
.C(n_1431),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1442),
.B(n_1416),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1442),
.B(n_1416),
.C(n_1431),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1446),
.B(n_1425),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1442),
.B(n_1431),
.C(n_1428),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_SL g1500 ( 
.A(n_1455),
.B(n_1430),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_L g1501 ( 
.A(n_1464),
.B(n_1431),
.C(n_1465),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1431),
.C(n_1424),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1474),
.B(n_1409),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1458),
.B(n_1403),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1478),
.B(n_1401),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1449),
.B(n_1406),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1478),
.B(n_1401),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1379),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1465),
.B(n_1424),
.C(n_1413),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1468),
.B(n_1424),
.C(n_1413),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1456),
.A2(n_1393),
.B1(n_1424),
.B2(n_1402),
.C(n_1386),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1437),
.A2(n_1433),
.B(n_1432),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1468),
.B(n_1477),
.C(n_1424),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1424),
.C(n_1406),
.Y(n_1514)
);

OAI211xp5_ASAP7_75t_L g1515 ( 
.A1(n_1456),
.A2(n_1401),
.B(n_1390),
.C(n_1407),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1452),
.A2(n_1401),
.B1(n_1386),
.B2(n_1402),
.Y(n_1516)
);

AND2x2_ASAP7_75t_SL g1517 ( 
.A(n_1470),
.B(n_1401),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1473),
.A2(n_1430),
.B1(n_1402),
.B2(n_1435),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1448),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1437),
.A2(n_1390),
.B1(n_1419),
.B2(n_1420),
.C(n_1421),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1473),
.A2(n_1435),
.B1(n_1432),
.B2(n_1433),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1437),
.B(n_1379),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1453),
.A2(n_1434),
.B1(n_1358),
.B2(n_1397),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1450),
.B(n_1391),
.C(n_1392),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1481),
.B(n_1471),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1519),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1505),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1480),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1507),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1517),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1480),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1454),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1517),
.A2(n_1451),
.B(n_1440),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1503),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1522),
.Y(n_1536)
);

NAND5xp2_ASAP7_75t_L g1537 ( 
.A(n_1479),
.B(n_1435),
.C(n_1433),
.D(n_1432),
.E(n_1414),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1522),
.B(n_1454),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1508),
.B(n_1475),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1492),
.B(n_1441),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1524),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1484),
.B(n_1441),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1504),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1482),
.B(n_1258),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1506),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1457),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1498),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1467),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1520),
.B(n_1440),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1497),
.B(n_1441),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1506),
.B(n_1457),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1521),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1536),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1530),
.B(n_1521),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1543),
.B(n_1487),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1539),
.B(n_1462),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1526),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1552),
.A2(n_1494),
.B(n_1509),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1543),
.B(n_1463),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1526),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1463),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1551),
.B(n_1489),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1528),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1528),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1531),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1547),
.A2(n_1488),
.B1(n_1485),
.B2(n_1523),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1539),
.B(n_1510),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1539),
.B(n_1513),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1552),
.B(n_1499),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1539),
.B(n_1502),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1553),
.B(n_1461),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1553),
.B(n_1469),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1541),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1545),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1532),
.B(n_1490),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1532),
.B(n_1444),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1542),
.B(n_1460),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1544),
.B(n_1460),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1549),
.B(n_1541),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1525),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1558),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1529),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.B(n_1573),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1562),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1575),
.B(n_1529),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1575),
.B(n_1527),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1562),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1576),
.B(n_1573),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1560),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1590),
.B(n_1544),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1583),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1565),
.B(n_1554),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1584),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1574),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1558),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1567),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1574),
.B(n_1534),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1574),
.B(n_1534),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1584),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1564),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1568),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1556),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1590),
.B(n_1554),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1556),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.B(n_1538),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1557),
.B(n_1556),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1569),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1569),
.Y(n_1621)
);

AOI21xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1563),
.A2(n_1548),
.B(n_1483),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1570),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1570),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1571),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1572),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1630)
);

NOR3x1_ASAP7_75t_L g1631 ( 
.A(n_1587),
.B(n_1555),
.C(n_1514),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1581),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1559),
.B(n_1533),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1628),
.B(n_1277),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

INVx3_ASAP7_75t_SL g1636 ( 
.A(n_1599),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1633),
.B(n_1589),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1594),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1605),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1630),
.B(n_1587),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1555),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1633),
.B(n_1589),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1607),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1604),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1628),
.B(n_1577),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1630),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1633),
.B(n_1589),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1622),
.B(n_1578),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1605),
.B(n_1537),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1593),
.A2(n_1537),
.B1(n_1547),
.B2(n_1518),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1593),
.A2(n_1518),
.B1(n_1549),
.B2(n_1550),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1605),
.B(n_1561),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1593),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1561),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1622),
.B(n_1277),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1602),
.B(n_1578),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1596),
.B(n_1582),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1598),
.B(n_1549),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1602),
.B(n_1585),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1604),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1598),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1632),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1613),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1617),
.B(n_1585),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1598),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1596),
.Y(n_1669)
);

INVxp33_ASAP7_75t_SL g1670 ( 
.A(n_1658),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1617),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

AOI222xp33_ASAP7_75t_L g1674 ( 
.A1(n_1636),
.A2(n_1595),
.B1(n_1614),
.B2(n_1603),
.C1(n_1592),
.C2(n_1608),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1645),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

O2A1O1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1651),
.A2(n_1595),
.B(n_1614),
.C(n_1603),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1617),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1652),
.A2(n_1592),
.B(n_1608),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1656),
.A2(n_1592),
.B1(n_1609),
.B2(n_1608),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1669),
.A2(n_1616),
.B(n_1625),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1665),
.Y(n_1684)
);

NOR4xp25_ASAP7_75t_SL g1685 ( 
.A(n_1647),
.B(n_1625),
.C(n_1631),
.D(n_1511),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1634),
.B(n_1500),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1664),
.B(n_1611),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1631),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1668),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1668),
.B(n_1629),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1653),
.A2(n_1491),
.B1(n_1609),
.B2(n_1540),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1662),
.B(n_1609),
.C(n_1616),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1667),
.B(n_1613),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1648),
.A2(n_1601),
.B(n_1629),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1659),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1675),
.B(n_1667),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1684),
.B(n_1637),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1690),
.B(n_1644),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1679),
.A2(n_1689),
.B1(n_1674),
.B2(n_1692),
.C(n_1677),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1690),
.B(n_1644),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1672),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1694),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1678),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1682),
.B(n_1650),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1673),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1639),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1683),
.B(n_1642),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1693),
.B(n_1655),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1654),
.B1(n_1642),
.B2(n_1691),
.C(n_1685),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1713),
.A2(n_1642),
.B(n_1639),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1676),
.B(n_1681),
.C(n_1680),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1718)
);

AOI211x1_ASAP7_75t_L g1719 ( 
.A1(n_1703),
.A2(n_1686),
.B(n_1646),
.C(n_1635),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1713),
.A2(n_1660),
.B1(n_1666),
.B2(n_1663),
.C(n_1601),
.Y(n_1720)
);

O2A1O1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1712),
.A2(n_1666),
.B(n_1661),
.C(n_1655),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1327),
.Y(n_1722)
);

AOI222xp33_ASAP7_75t_L g1723 ( 
.A1(n_1700),
.A2(n_1657),
.B1(n_1655),
.B2(n_1661),
.C1(n_1550),
.C2(n_1613),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1698),
.A2(n_1708),
.B1(n_1696),
.B2(n_1707),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_SL g1725 ( 
.A(n_1700),
.B(n_1493),
.C(n_1615),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1701),
.A2(n_1657),
.B1(n_1661),
.B2(n_1615),
.Y(n_1726)
);

NAND4xp25_ASAP7_75t_SL g1727 ( 
.A(n_1699),
.B(n_1615),
.C(n_1620),
.D(n_1600),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1725),
.A2(n_1710),
.B1(n_1709),
.B2(n_1714),
.Y(n_1728)
);

NOR4xp25_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1711),
.C(n_1705),
.D(n_1704),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1718),
.B(n_1706),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1722),
.B(n_1702),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1721),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1724),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1719),
.B(n_1710),
.C(n_1657),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1723),
.B(n_1586),
.Y(n_1735)
);

AOI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1716),
.A2(n_1612),
.B(n_1610),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1610),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1720),
.A2(n_1266),
.B1(n_1337),
.B2(n_1258),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1728),
.A2(n_1727),
.B(n_1600),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1733),
.A2(n_1620),
.B(n_1626),
.C(n_1612),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1730),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1729),
.B(n_1306),
.C(n_1591),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1736),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1732),
.B(n_1731),
.C(n_1734),
.Y(n_1744)
);

NOR2xp67_ASAP7_75t_L g1745 ( 
.A(n_1743),
.B(n_1737),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1738),
.B1(n_1735),
.B2(n_1618),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1742),
.A2(n_1306),
.B1(n_1258),
.B2(n_1549),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1741),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1739),
.A2(n_1618),
.B(n_1619),
.C(n_1626),
.Y(n_1749)
);

AO22x2_ASAP7_75t_L g1750 ( 
.A1(n_1740),
.A2(n_1627),
.B1(n_1624),
.B2(n_1623),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1745),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1748),
.B(n_1746),
.Y(n_1752)
);

NAND4xp75_ASAP7_75t_L g1753 ( 
.A(n_1747),
.B(n_1619),
.C(n_1264),
.D(n_1282),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1749),
.B(n_1264),
.C(n_1282),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1750),
.A2(n_1606),
.B1(n_1591),
.B2(n_1624),
.C(n_1623),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1751),
.A2(n_1623),
.B(n_1621),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1627),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1754),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1757),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1759),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1760),
.B(n_1758),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1753),
.B1(n_1756),
.B2(n_1755),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1627),
.B(n_1624),
.Y(n_1763)
);

OAI22x1_ASAP7_75t_SL g1764 ( 
.A1(n_1762),
.A2(n_1264),
.B1(n_1606),
.B2(n_1591),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1764),
.B(n_1606),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1763),
.B(n_1621),
.Y(n_1766)
);

OAI21x1_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1621),
.B(n_1566),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_SL g1768 ( 
.A(n_1767),
.B(n_1765),
.C(n_1360),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1273),
.B1(n_1360),
.B2(n_1297),
.C(n_1299),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1273),
.B(n_1540),
.C(n_1423),
.Y(n_1770)
);


endmodule