module fake_jpeg_15290_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_29),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx3_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_53),
.Y(n_61)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_20),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_77),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_39),
.B1(n_45),
.B2(n_37),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_5),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_15),
.B1(n_32),
.B2(n_31),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_77),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_5),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_7),
.B(n_8),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_6),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.C(n_93),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_78),
.C(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_9),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_89),
.C(n_12),
.Y(n_99)
);

AOI321xp33_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_100),
.A3(n_33),
.B1(n_14),
.B2(n_16),
.C(n_19),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_13),
.C(n_21),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_22),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_23),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_24),
.C(n_26),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_27),
.C(n_28),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_30),
.Y(n_107)
);


endmodule