module fake_jpeg_29087_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_32),
.C(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_1),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_84),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_20),
.B1(n_19),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_20),
.B1(n_18),
.B2(n_24),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_18),
.B1(n_15),
.B2(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_76),
.B1(n_90),
.B2(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_80),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_16),
.B1(n_30),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_15),
.B1(n_22),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_15),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_92),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_35),
.B(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_30),
.B1(n_6),
.B2(n_7),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_41),
.A2(n_30),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_37),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_36),
.B(n_9),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_67),
.B(n_60),
.C(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_35),
.B(n_37),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_102),
.Y(n_144)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_108),
.Y(n_121)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_69),
.C(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_114),
.B1(n_72),
.B2(n_76),
.Y(n_126)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_84),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_84),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_112),
.B1(n_113),
.B2(n_120),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_65),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_150),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_120),
.B1(n_113),
.B2(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_154),
.B1(n_163),
.B2(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_68),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_160),
.A3(n_162),
.B1(n_126),
.B2(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_101),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_105),
.B(n_115),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_129),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_117),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_116),
.B1(n_109),
.B2(n_111),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_175),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_136),
.B1(n_127),
.B2(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_178),
.B1(n_152),
.B2(n_132),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_177),
.B(n_162),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_145),
.C(n_157),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_174),
.C(n_56),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_153),
.B(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_184),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_148),
.B(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_156),
.B(n_159),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_187),
.C(n_167),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_158),
.B(n_160),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_145),
.A3(n_147),
.B1(n_146),
.B2(n_158),
.C1(n_150),
.C2(n_125),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_132),
.A3(n_128),
.B1(n_122),
.B2(n_103),
.C1(n_106),
.C2(n_102),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_178),
.B1(n_185),
.B2(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_128),
.B1(n_122),
.B2(n_88),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_165),
.C(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_172),
.B(n_174),
.C(n_170),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.C(n_128),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_189),
.B1(n_182),
.B2(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_190),
.B1(n_196),
.B2(n_56),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_202),
.Y(n_206)
);

NAND4xp25_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_143),
.C(n_61),
.D(n_70),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_208),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_87),
.C(n_88),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_198),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_199),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_209),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_206),
.B(n_207),
.Y(n_216)
);


endmodule