module real_aes_2662_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_0), .B(n_225), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_1), .A2(n_233), .B(n_238), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g86 ( .A1(n_2), .A2(n_66), .B1(n_87), .B2(n_106), .Y(n_86) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_3), .A2(n_55), .B1(n_93), .B2(n_94), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_4), .B(n_240), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_5), .A2(n_70), .B1(n_183), .B2(n_184), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_5), .Y(n_184) );
INVx1_ASAP7_75t_L g206 ( .A(n_6), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_7), .B(n_240), .Y(n_330) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_8), .A2(n_22), .B1(n_93), .B2(n_97), .Y(n_96) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_9), .B(n_242), .Y(n_322) );
INVx2_ASAP7_75t_L g222 ( .A(n_10), .Y(n_222) );
AOI221x1_ASAP7_75t_L g264 ( .A1(n_11), .A2(n_19), .B1(n_225), .B2(n_233), .C(n_265), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_12), .A2(n_41), .B1(n_124), .B2(n_129), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_13), .B(n_225), .Y(n_318) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_14), .A2(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_15), .B(n_244), .Y(n_268) );
INVx1_ASAP7_75t_L g191 ( .A(n_16), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_16), .B(n_240), .Y(n_253) );
AO21x1_ASAP7_75t_L g274 ( .A1(n_17), .A2(n_225), .B(n_275), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_18), .A2(n_44), .B1(n_149), .B2(n_152), .Y(n_148) );
INVx1_ASAP7_75t_L g551 ( .A(n_19), .Y(n_551) );
NAND2x1_ASAP7_75t_L g296 ( .A(n_20), .B(n_240), .Y(n_296) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_21), .B(n_242), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g198 ( .A1(n_22), .A2(n_55), .B1(n_60), .B2(n_199), .C(n_201), .Y(n_198) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_23), .A2(n_67), .B(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g246 ( .A(n_23), .B(n_67), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_24), .B(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_26), .B(n_240), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_27), .B(n_242), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_28), .A2(n_233), .B(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_29), .A2(n_35), .B1(n_112), .B2(n_120), .Y(n_111) );
INVx1_ASAP7_75t_SL g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g208 ( .A(n_31), .Y(n_208) );
AND2x2_ASAP7_75t_L g231 ( .A(n_31), .B(n_206), .Y(n_231) );
AND2x2_ASAP7_75t_L g234 ( .A(n_31), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_32), .B(n_225), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_33), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_34), .B(n_242), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_36), .A2(n_233), .B(n_328), .Y(n_327) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_37), .A2(n_60), .B1(n_93), .B2(n_100), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_38), .A2(n_81), .B1(n_82), .B2(n_177), .Y(n_80) );
INVx1_ASAP7_75t_L g177 ( .A(n_38), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_39), .B(n_242), .Y(n_297) );
INVx1_ASAP7_75t_L g228 ( .A(n_40), .Y(n_228) );
INVx1_ASAP7_75t_L g237 ( .A(n_40), .Y(n_237) );
INVx1_ASAP7_75t_L g105 ( .A(n_42), .Y(n_105) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_43), .A2(n_52), .B1(n_157), .B2(n_160), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_45), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_45), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_46), .B(n_240), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_46), .A2(n_81), .B1(n_82), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_46), .Y(n_532) );
XOR2xp5_ASAP7_75t_L g538 ( .A(n_47), .B(n_81), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_48), .A2(n_233), .B(n_295), .Y(n_294) );
AO21x1_ASAP7_75t_L g276 ( .A1(n_49), .A2(n_233), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_50), .B(n_225), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_51), .A2(n_64), .B1(n_166), .B2(n_171), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_53), .A2(n_61), .B1(n_134), .B2(n_137), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_54), .B(n_225), .Y(n_331) );
INVxp33_ASAP7_75t_L g203 ( .A(n_55), .Y(n_203) );
AND2x2_ASAP7_75t_L g290 ( .A(n_56), .B(n_245), .Y(n_290) );
INVx1_ASAP7_75t_L g230 ( .A(n_57), .Y(n_230) );
INVx1_ASAP7_75t_L g235 ( .A(n_57), .Y(n_235) );
AND2x2_ASAP7_75t_L g333 ( .A(n_58), .B(n_219), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_59), .B(n_142), .Y(n_141) );
INVxp67_ASAP7_75t_L g202 ( .A(n_60), .Y(n_202) );
AND2x2_ASAP7_75t_L g218 ( .A(n_62), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_63), .B(n_225), .Y(n_255) );
AND2x2_ASAP7_75t_L g275 ( .A(n_65), .B(n_249), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_68), .B(n_242), .Y(n_254) );
AND2x2_ASAP7_75t_L g299 ( .A(n_69), .B(n_219), .Y(n_299) );
INVx1_ASAP7_75t_L g183 ( .A(n_70), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_71), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_71), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_71), .B(n_240), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_72), .A2(n_233), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_73), .B(n_242), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_74), .B(n_240), .Y(n_239) );
BUFx2_ASAP7_75t_L g187 ( .A(n_75), .Y(n_187) );
BUFx2_ASAP7_75t_SL g200 ( .A(n_76), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_77), .A2(n_233), .B(n_320), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_195), .B1(n_209), .B2(n_529), .C(n_530), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_178), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NOR2x1_ASAP7_75t_L g84 ( .A(n_85), .B(n_140), .Y(n_84) );
NAND4xp25_ASAP7_75t_L g85 ( .A(n_86), .B(n_111), .C(n_123), .D(n_133), .Y(n_85) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_98), .Y(n_90) );
AND2x4_ASAP7_75t_L g139 ( .A(n_91), .B(n_122), .Y(n_139) );
AND2x2_ASAP7_75t_L g170 ( .A(n_91), .B(n_118), .Y(n_170) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_95), .Y(n_91) );
AND2x2_ASAP7_75t_L g110 ( .A(n_92), .B(n_96), .Y(n_110) );
INVx2_ASAP7_75t_L g117 ( .A(n_92), .Y(n_117) );
INVx1_ASAP7_75t_L g94 ( .A(n_93), .Y(n_94) );
INVx2_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
INVx1_ASAP7_75t_L g100 ( .A(n_93), .Y(n_100) );
OAI22x1_ASAP7_75t_L g102 ( .A1(n_93), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_93), .Y(n_103) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_95), .Y(n_176) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
AND2x4_ASAP7_75t_L g132 ( .A(n_96), .B(n_117), .Y(n_132) );
AND2x2_ASAP7_75t_L g136 ( .A(n_98), .B(n_115), .Y(n_136) );
AND2x4_ASAP7_75t_L g151 ( .A(n_98), .B(n_132), .Y(n_151) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_101), .Y(n_98) );
BUFx2_ASAP7_75t_L g109 ( .A(n_99), .Y(n_109) );
INVx2_ASAP7_75t_L g119 ( .A(n_99), .Y(n_119) );
AND2x2_ASAP7_75t_L g147 ( .A(n_99), .B(n_102), .Y(n_147) );
AND2x4_ASAP7_75t_L g122 ( .A(n_101), .B(n_119), .Y(n_122) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g118 ( .A(n_102), .B(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_102), .Y(n_164) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx5_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g121 ( .A(n_110), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g163 ( .A(n_110), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx6_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
AND2x4_ASAP7_75t_L g128 ( .A(n_115), .B(n_122), .Y(n_128) );
AND2x2_ASAP7_75t_L g146 ( .A(n_115), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVxp67_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
AND2x2_ASAP7_75t_L g159 ( .A(n_118), .B(n_132), .Y(n_159) );
BUFx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g131 ( .A(n_122), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx8_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND4xp25_ASAP7_75t_SL g140 ( .A(n_141), .B(n_148), .C(n_156), .D(n_165), .Y(n_140) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g154 ( .A(n_147), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g174 ( .A(n_147), .B(n_175), .Y(n_174) );
BUFx4f_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_190), .B2(n_194), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B1(n_185), .B2(n_186), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_187), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_190), .Y(n_194) );
INVx1_ASAP7_75t_L g193 ( .A(n_191), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_197), .Y(n_196) );
AND3x1_ASAP7_75t_SL g197 ( .A(n_198), .B(n_204), .C(n_207), .Y(n_197) );
INVxp67_ASAP7_75t_L g537 ( .A(n_198), .Y(n_537) );
CKINVDCx8_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_204), .Y(n_535) );
AO21x1_ASAP7_75t_SL g544 ( .A1(n_204), .A2(n_545), .B(n_549), .Y(n_544) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_SL g541 ( .A(n_205), .B(n_207), .Y(n_541) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g236 ( .A(n_206), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_207), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2x1p5_ASAP7_75t_L g546 ( .A(n_208), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
NOR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_416), .Y(n_211) );
AO211x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_258), .B(n_309), .C(n_384), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND3x2_ASAP7_75t_L g465 ( .A(n_215), .B(n_346), .C(n_362), .Y(n_465) );
AND2x4_ASAP7_75t_L g468 ( .A(n_215), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_247), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_216), .B(n_324), .Y(n_323) );
INVx4_ASAP7_75t_L g377 ( .A(n_216), .Y(n_377) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_216), .B(n_371), .Y(n_462) );
AND2x2_ASAP7_75t_L g505 ( .A(n_216), .B(n_325), .Y(n_505) );
INVx5_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g354 ( .A(n_217), .Y(n_354) );
AND2x2_ASAP7_75t_L g373 ( .A(n_217), .B(n_315), .Y(n_373) );
AND2x2_ASAP7_75t_L g391 ( .A(n_217), .B(n_325), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_217), .B(n_324), .Y(n_451) );
NOR2x1_ASAP7_75t_SL g478 ( .A(n_217), .B(n_247), .Y(n_478) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_223), .Y(n_217) );
INVx3_ASAP7_75t_L g289 ( .A(n_219), .Y(n_289) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx4f_ASAP7_75t_L g316 ( .A(n_221), .Y(n_316) );
AND2x2_ASAP7_75t_SL g245 ( .A(n_222), .B(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_L g249 ( .A(n_222), .B(n_246), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_232), .B(n_244), .Y(n_223) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_225), .Y(n_529) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AND2x6_ASAP7_75t_L g242 ( .A(n_227), .B(n_235), .Y(n_242) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g240 ( .A(n_229), .B(n_237), .Y(n_240) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx5_ASAP7_75t_L g243 ( .A(n_231), .Y(n_243) );
AND2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g548 ( .A(n_235), .Y(n_548) );
INVx2_ASAP7_75t_L g550 ( .A(n_237), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_241), .B(n_243), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_243), .A2(n_253), .B(n_254), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_243), .A2(n_266), .B(n_267), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_278), .B(n_279), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_243), .A2(n_286), .B(n_287), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_243), .A2(n_296), .B(n_297), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_243), .A2(n_321), .B(n_322), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_243), .A2(n_329), .B(n_330), .Y(n_328) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_264), .B(n_268), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_244), .Y(n_332) );
OA21x2_ASAP7_75t_L g337 ( .A1(n_244), .A2(n_264), .B(n_268), .Y(n_337) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_247), .B(n_315), .Y(n_314) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_256), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_248), .B(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_248), .A2(n_250), .B(n_256), .Y(n_350) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_249), .B(n_281), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_249), .A2(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
AO21x1_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_291), .B(n_300), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_260), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_359) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
AND2x2_ASAP7_75t_L g420 ( .A(n_261), .B(n_306), .Y(n_420) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g353 ( .A(n_262), .B(n_336), .Y(n_353) );
AND2x2_ASAP7_75t_L g425 ( .A(n_262), .B(n_308), .Y(n_425) );
AND2x2_ASAP7_75t_L g444 ( .A(n_262), .B(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_263), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_269), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g404 ( .A(n_270), .B(n_303), .Y(n_404) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_282), .Y(n_270) );
AND2x2_ASAP7_75t_L g306 ( .A(n_271), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g341 ( .A(n_271), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_271), .B(n_337), .Y(n_401) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g494 ( .A(n_272), .Y(n_494) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
OAI21x1_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_276), .B(n_280), .Y(n_273) );
INVx1_ASAP7_75t_L g281 ( .A(n_275), .Y(n_281) );
INVx2_ASAP7_75t_L g342 ( .A(n_282), .Y(n_342) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_282), .Y(n_442) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_289), .B(n_290), .Y(n_282) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_283), .A2(n_289), .B(n_290), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_288), .Y(n_283) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_289), .A2(n_293), .B(n_299), .Y(n_292) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_289), .A2(n_293), .B(n_299), .Y(n_305) );
INVx2_ASAP7_75t_L g338 ( .A(n_291), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_291), .B(n_470), .Y(n_496) );
AND2x2_ASAP7_75t_L g515 ( .A(n_291), .B(n_505), .Y(n_515) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_292), .B(n_342), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g382 ( .A(n_301), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_301), .B(n_352), .Y(n_387) );
INVx1_ASAP7_75t_SL g514 ( .A(n_301), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_302), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
AND2x2_ASAP7_75t_L g526 ( .A(n_303), .B(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g402 ( .A(n_304), .B(n_307), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_304), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g456 ( .A(n_304), .B(n_308), .Y(n_456) );
AND2x2_ASAP7_75t_L g487 ( .A(n_304), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g352 ( .A(n_305), .B(n_308), .Y(n_352) );
INVxp67_ASAP7_75t_L g369 ( .A(n_305), .Y(n_369) );
BUFx3_ASAP7_75t_L g410 ( .A(n_305), .Y(n_410) );
AND2x2_ASAP7_75t_L g430 ( .A(n_306), .B(n_431), .Y(n_430) );
NAND2xp33_ASAP7_75t_L g443 ( .A(n_306), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_307), .B(n_336), .Y(n_399) );
AND2x2_ASAP7_75t_L g488 ( .A(n_307), .B(n_337), .Y(n_488) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g415 ( .A(n_308), .B(n_337), .Y(n_415) );
OR3x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_359), .C(n_374), .Y(n_309) );
OAI321xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_323), .A3(n_334), .B1(n_339), .B2(n_343), .C(n_351), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_314), .Y(n_390) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_314), .Y(n_408) );
OR2x2_ASAP7_75t_L g412 ( .A(n_314), .B(n_323), .Y(n_412) );
BUFx3_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
AND2x2_ASAP7_75t_L g363 ( .A(n_315), .B(n_349), .Y(n_363) );
INVx1_ASAP7_75t_L g380 ( .A(n_315), .Y(n_380) );
INVx2_ASAP7_75t_L g396 ( .A(n_315), .Y(n_396) );
OR2x2_ASAP7_75t_L g435 ( .A(n_315), .B(n_324), .Y(n_435) );
INVx2_ASAP7_75t_L g423 ( .A(n_323), .Y(n_423) );
AND2x2_ASAP7_75t_L g347 ( .A(n_324), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
AND2x4_ASAP7_75t_L g371 ( .A(n_324), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_324), .B(n_348), .Y(n_394) );
AND2x2_ASAP7_75t_L g501 ( .A(n_324), .B(n_396), .Y(n_501) );
INVx4_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_325), .Y(n_460) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_332), .B(n_333), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
INVx1_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x2_ASAP7_75t_L g475 ( .A(n_335), .B(n_402), .Y(n_475) );
INVx1_ASAP7_75t_SL g492 ( .A(n_335), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_335), .B(n_468), .Y(n_521) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
OR2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_337), .Y(n_364) );
AND2x2_ASAP7_75t_L g457 ( .A(n_338), .B(n_353), .Y(n_457) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_342), .B(n_353), .Y(n_480) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_344), .A2(n_493), .B1(n_498), .B2(n_500), .Y(n_497) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x2_ASAP7_75t_L g422 ( .A(n_345), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g517 ( .A(n_345), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g473 ( .A(n_346), .B(n_391), .Y(n_473) );
AND2x4_ASAP7_75t_L g427 ( .A(n_347), .B(n_373), .Y(n_427) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_349), .Y(n_525) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g358 ( .A(n_350), .Y(n_358) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .C(n_354), .D(n_355), .Y(n_351) );
AND2x2_ASAP7_75t_L g509 ( .A(n_352), .B(n_494), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_352), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_353), .B(n_429), .Y(n_428) );
OAI322xp33_ASAP7_75t_L g436 ( .A1(n_353), .A2(n_437), .A3(n_441), .B1(n_443), .B2(n_445), .C1(n_447), .C2(n_452), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_353), .B(n_402), .Y(n_452) );
INVx1_ASAP7_75t_L g520 ( .A(n_353), .Y(n_520) );
INVx2_ASAP7_75t_L g366 ( .A(n_354), .Y(n_366) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_357), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_358), .B(n_377), .Y(n_434) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
AND2x2_ASAP7_75t_L g479 ( .A(n_362), .B(n_390), .Y(n_479) );
AOI31xp33_ASAP7_75t_L g365 ( .A1(n_363), .A2(n_366), .A3(n_367), .B(n_370), .Y(n_365) );
AND2x2_ASAP7_75t_L g376 ( .A(n_363), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g504 ( .A(n_363), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_363), .B(n_391), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_363), .Y(n_512) );
INVx1_ASAP7_75t_SL g470 ( .A(n_364), .Y(n_470) );
NAND3xp33_ASAP7_75t_SL g498 ( .A(n_364), .B(n_492), .C(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g398 ( .A(n_369), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x2_ASAP7_75t_L g379 ( .A(n_371), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g440 ( .A(n_371), .Y(n_440) );
AOI322xp5_ASAP7_75t_L g522 ( .A1(n_371), .A2(n_401), .A3(n_404), .B1(n_523), .B2(n_524), .C1(n_526), .C2(n_528), .Y(n_522) );
AND2x2_ASAP7_75t_L g528 ( .A(n_371), .B(n_377), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B(n_381), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_377), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g523 ( .A(n_377), .B(n_410), .Y(n_523) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
AND2x2_ASAP7_75t_L g477 ( .A(n_380), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g524 ( .A(n_380), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g429 ( .A(n_383), .Y(n_429) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
O2A1O1Ixp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_389), .C(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g446 ( .A(n_391), .B(n_396), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_397), .B(n_403), .C(n_405), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_419), .B1(n_421), .B2(n_424), .C(n_426), .Y(n_418) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g438 ( .A(n_395), .Y(n_438) );
OR2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g503 ( .A(n_398), .Y(n_503) );
INVx1_ASAP7_75t_L g527 ( .A(n_399), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AND2x2_ASAP7_75t_L g409 ( .A(n_401), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_401), .B(n_471), .Y(n_483) );
INVx1_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_411), .B2(n_413), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_SL g471 ( .A(n_410), .Y(n_471) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND4xp75_ASAP7_75t_L g416 ( .A(n_417), .B(n_453), .C(n_481), .D(n_506), .Y(n_416) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_418), .B(n_436), .Y(n_417) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_425), .B(n_494), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_430), .B2(n_432), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_429), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx2_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
OR2x2_ASAP7_75t_L g484 ( .A(n_435), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_446), .A2(n_491), .B(n_493), .Y(n_490) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_461), .B2(n_463), .C(n_464), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_456), .A2(n_503), .B(n_504), .Y(n_502) );
INVx3_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
OAI322xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_470), .A3(n_471), .B1(n_472), .B2(n_474), .C1(n_476), .C2(n_480), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
INVx1_ASAP7_75t_L g485 ( .A(n_478), .Y(n_485) );
AND2x2_ASAP7_75t_L g500 ( .A(n_478), .B(n_501), .Y(n_500) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_495), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_486), .B2(n_489), .C(n_490), .Y(n_482) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OAI211xp5_ASAP7_75t_SL g495 ( .A1(n_489), .A2(n_496), .B(n_497), .C(n_502), .Y(n_495) );
INVx2_ASAP7_75t_SL g518 ( .A(n_505), .Y(n_518) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI211xp5_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_519), .B(n_521), .C(n_522), .Y(n_516) );
OAI222xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_533), .B1(n_538), .B2(n_539), .C1(n_542), .C2(n_551), .Y(n_530) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
endmodule