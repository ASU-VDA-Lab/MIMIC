module fake_jpeg_8384_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_57),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_48),
.B(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_24),
.B1(n_22),
.B2(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_25),
.A3(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_69),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_67),
.Y(n_103)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_26),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_74),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_81),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_40),
.B(n_38),
.C(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_88),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_39),
.B1(n_36),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_43),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_101),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_50),
.B1(n_64),
.B2(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_96),
.B1(n_25),
.B2(n_43),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_29),
.B1(n_17),
.B2(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_105),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_36),
.B1(n_65),
.B2(n_67),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_36),
.B1(n_68),
.B2(n_41),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_84),
.B(n_82),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_127),
.B(n_129),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_127),
.B1(n_126),
.B2(n_94),
.Y(n_136)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_122),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_33),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_51),
.C(n_56),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_70),
.C(n_74),
.Y(n_140)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_35),
.B(n_33),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_121),
.Y(n_139)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_135),
.B(n_138),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_164),
.B(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_144),
.C(n_116),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_98),
.B1(n_93),
.B2(n_81),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_156),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_78),
.B1(n_73),
.B2(n_77),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_95),
.B1(n_79),
.B2(n_71),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_79),
.C(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_149),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_157),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_43),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_116),
.B(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_71),
.B1(n_75),
.B2(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_73),
.B(n_53),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_169),
.Y(n_204)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_124),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_173),
.C(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_194),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_178),
.B(n_189),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_108),
.A3(n_110),
.B1(n_130),
.B2(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_108),
.B(n_110),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_87),
.B(n_115),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_182),
.Y(n_199)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_115),
.C(n_122),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_149),
.B(n_146),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_133),
.B(n_122),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_133),
.B1(n_75),
.B2(n_53),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_92),
.C(n_53),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_0),
.C(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_142),
.CI(n_155),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_176),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_154),
.C(n_138),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_135),
.B1(n_152),
.B2(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_157),
.B1(n_164),
.B2(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_162),
.B1(n_35),
.B2(n_28),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_35),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_191),
.C(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_173),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_225),
.C(n_227),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_181),
.C(n_193),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_185),
.B1(n_190),
.B2(n_189),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_237),
.B1(n_212),
.B2(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_238),
.B1(n_215),
.B2(n_196),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_185),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_218),
.C(n_217),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_235),
.B(n_236),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_182),
.B(n_174),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_165),
.B1(n_184),
.B2(n_166),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_250),
.B1(n_231),
.B2(n_230),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_206),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_200),
.B1(n_203),
.B2(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_249),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_195),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_251),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_222),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_195),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_201),
.C(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_196),
.B1(n_213),
.B2(n_216),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_237),
.B(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_216),
.B1(n_180),
.B2(n_177),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_222),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_229),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_219),
.B(n_2),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_247),
.A3(n_251),
.B1(n_241),
.B2(n_246),
.C1(n_249),
.C2(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_267),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_265),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_5),
.Y(n_267)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_243),
.C(n_266),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_243),
.B1(n_9),
.B2(n_10),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_12),
.B(n_13),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_11),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_11),
.C(n_12),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_12),
.Y(n_284)
);

AOI211xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_260),
.B(n_255),
.C(n_263),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_272),
.B(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_284),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_263),
.B1(n_13),
.B2(n_15),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_270),
.C(n_273),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_274),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_289),
.A2(n_279),
.B(n_278),
.C(n_284),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_276),
.B(n_13),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_16),
.C(n_293),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_292),
.Y(n_297)
);


endmodule