module real_jpeg_16909_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_594;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_617),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_0),
.B(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_1),
.Y(n_452)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_2),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_3),
.A2(n_72),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_3),
.A2(n_253),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_3),
.A2(n_253),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_3),
.A2(n_253),
.B1(n_525),
.B2(n_528),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_4),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_4),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_4),
.A2(n_322),
.B1(n_390),
.B2(n_395),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_4),
.A2(n_322),
.B1(n_517),
.B2(n_520),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_4),
.A2(n_322),
.B1(n_558),
.B2(n_561),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_54),
.B1(n_128),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_5),
.A2(n_131),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_5),
.A2(n_131),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_5),
.A2(n_131),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_6),
.A2(n_37),
.B1(n_105),
.B2(n_109),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_37),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_6),
.A2(n_37),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_7),
.A2(n_52),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_7),
.A2(n_52),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_52),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_8),
.A2(n_71),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_8),
.A2(n_71),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_8),
.A2(n_71),
.B1(n_241),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_9),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_9),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_9),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_10),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_10),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_11),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_11),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_11),
.A2(n_249),
.B1(n_369),
.B2(n_374),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_11),
.A2(n_249),
.B1(n_458),
.B2(n_464),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_11),
.A2(n_249),
.B1(n_540),
.B2(n_543),
.Y(n_539)
);

OAI32xp33_ASAP7_75t_L g286 ( 
.A1(n_12),
.A2(n_287),
.A3(n_291),
.B1(n_293),
.B2(n_299),
.Y(n_286)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_12),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_12),
.A2(n_38),
.B1(n_298),
.B2(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_12),
.B(n_24),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_12),
.A2(n_343),
.A3(n_438),
.B1(n_443),
.B2(n_446),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_12),
.A2(n_298),
.B1(n_473),
.B2(n_475),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_12),
.B(n_76),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_12),
.B(n_220),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_12),
.B(n_135),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_13),
.Y(n_618)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_16),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_16),
.Y(n_143)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_16),
.Y(n_267)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_168),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_22),
.B(n_65),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_23),
.A2(n_56),
.B(n_250),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

OR2x6_ASAP7_75t_SL g56 ( 
.A(n_24),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_24),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_24),
.A2(n_55),
.B1(n_318),
.B2(n_325),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_26),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_30),
.Y(n_182)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_31),
.Y(n_345)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_36),
.Y(n_420)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_46),
.A2(n_127),
.B(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_55),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_50),
.Y(n_321)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_67),
.B(n_74),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_67),
.B1(n_127),
.B2(n_132),
.Y(n_126)
);

OAI22x1_ASAP7_75t_SL g244 ( 
.A1(n_56),
.A2(n_132),
.B1(n_245),
.B2(n_250),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_56),
.A2(n_132),
.B1(n_319),
.B2(n_362),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_56),
.A2(n_74),
.B(n_420),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_61),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_61),
.Y(n_366)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_62),
.Y(n_292)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_65),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_65),
.B(n_173),
.Y(n_616)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_75),
.CI(n_111),
.CON(n_65),
.SN(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_72),
.B(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_89),
.B(n_103),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_76),
.B(n_114),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_76),
.A2(n_89),
.B1(n_179),
.B2(n_413),
.Y(n_412)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_81),
.Y(n_240)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_83),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_83),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_83),
.Y(n_521)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_114),
.B(n_123),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_89),
.A2(n_179),
.B(n_188),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_89),
.A2(n_123),
.B(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_90),
.A2(n_104),
.B(n_189),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_90),
.A2(n_124),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_90),
.A2(n_124),
.B1(n_279),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_90),
.A2(n_124),
.B1(n_368),
.B2(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_90),
.A2(n_124),
.B1(n_389),
.B2(n_472),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_98),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_98),
.Y(n_297)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_101),
.Y(n_284)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_108),
.Y(n_373)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_125),
.C(n_133),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_112),
.A2(n_113),
.B1(n_133),
.B2(n_134),
.Y(n_175)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_114),
.Y(n_341)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_176),
.C(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_134),
.B(n_178),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_146),
.B(n_157),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_135),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_135),
.B(n_229),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_135),
.A2(n_146),
.B1(n_513),
.B2(n_516),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_135),
.A2(n_146),
.B1(n_457),
.B2(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_136),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_136),
.B(n_158),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_136),
.A2(n_271),
.B1(n_456),
.B2(n_465),
.Y(n_455)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_139),
.Y(n_530)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_143),
.Y(n_499)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_143),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_146),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_146),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_146),
.A2(n_416),
.B(n_480),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_148),
.Y(n_507)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_150),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_150),
.Y(n_515)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g360 ( 
.A1(n_158),
.A2(n_271),
.B(n_335),
.Y(n_360)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21x1_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_190),
.B(n_615),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_174),
.A2(n_176),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_174),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_176),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_176),
.A2(n_594),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_177),
.B(n_592),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_181),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_187),
.Y(n_281)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_187),
.Y(n_377)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_589),
.B(n_612),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_426),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_352),
.B(n_403),
.C(n_404),
.D(n_425),
.Y(n_192)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_326),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_326),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_255),
.C(n_276),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_196),
.A2(n_255),
.B1(n_256),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_196),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_243),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_197),
.B(n_244),
.C(n_254),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_227),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_198),
.B(n_227),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_210),
.B(n_217),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_199),
.A2(n_210),
.B1(n_304),
.B2(n_312),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_199),
.A2(n_217),
.B(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_199),
.A2(n_538),
.B1(n_548),
.B2(n_549),
.Y(n_537)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_200),
.B(n_222),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_200),
.A2(n_262),
.B(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_200),
.A2(n_524),
.B(n_531),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_200),
.A2(n_220),
.B1(n_298),
.B2(n_557),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_200),
.A2(n_539),
.B1(n_557),
.B2(n_571),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_203),
.Y(n_542)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_204),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_205),
.Y(n_547)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_206),
.Y(n_572)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_216),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_226),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_228),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_231),
.Y(n_445)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_242),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_254),
.Y(n_243)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_269),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_257),
.B(n_269),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_268),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_258),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_259),
.Y(n_402)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_262),
.Y(n_454)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_267),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_268),
.A2(n_304),
.B(n_402),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_271),
.A2(n_272),
.B(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_276),
.B(n_354),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.C(n_317),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_277),
.B(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_303),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_286),
.B(n_303),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_290),
.Y(n_394)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_297),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_298),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_298),
.B(n_506),
.Y(n_505)
);

OAI21xp33_ASAP7_75t_SL g513 ( 
.A1(n_298),
.A2(n_505),
.B(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_311),
.Y(n_527)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_316),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_327),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_337),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_328),
.B(n_337),
.C(n_349),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_329),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_329),
.A2(n_336),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_334),
.Y(n_422)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g603 ( 
.A1(n_336),
.A2(n_421),
.B(n_604),
.Y(n_603)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_338),
.B(n_348),
.C(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.C(n_379),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_353),
.B(n_356),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.C(n_378),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_378),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.C(n_367),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_367),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_382),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_385),
.C(n_387),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_383),
.B(n_586),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_387),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_399),
.C(n_401),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_388),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_390),
.Y(n_475)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_399),
.A2(n_400),
.B1(n_401),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR3xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_428),
.C(n_431),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_407),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_408),
.B(n_423),
.C(n_607),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_417),
.B1(n_423),
.B2(n_424),
.Y(n_410)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_411),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_412),
.B(n_414),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_417),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_417),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_422),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_419),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g604 ( 
.A(n_422),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_583),
.B(n_588),
.Y(n_432)
);

AOI21x1_ASAP7_75t_SL g433 ( 
.A1(n_434),
.A2(n_486),
.B(n_582),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_476),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_435),
.B(n_476),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_455),
.C(n_471),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_436),
.B(n_579),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_453),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_453),
.Y(n_478)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_455),
.B(n_471),
.Y(n_579)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_481),
.B1(n_482),
.B2(n_485),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_478),
.B(n_479),
.C(n_481),
.Y(n_584)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_577),
.B(n_581),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_535),
.B(n_576),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_522),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_489),
.B(n_522),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_511),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_490),
.A2(n_511),
.B1(n_512),
.B2(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_490),
.Y(n_553)
);

OAI32xp33_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_496),
.A3(n_500),
.B1(n_505),
.B2(n_508),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_532),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_523),
.B(n_533),
.C(n_534),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_524),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_554),
.B(n_575),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_552),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_552),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_555),
.A2(n_569),
.B(n_574),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_556),
.B(n_564),
.Y(n_555)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_565),
.B(n_566),
.Y(n_564)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_570),
.B(n_573),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_573),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_SL g577 ( 
.A(n_578),
.B(n_580),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_578),
.B(n_580),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_585),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_584),
.B(n_585),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_590),
.B(n_605),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_590),
.A2(n_613),
.B(n_614),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_SL g590 ( 
.A(n_591),
.B(n_595),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_595),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_600),
.C(n_602),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_597),
.A2(n_600),
.B1(n_601),
.B2(n_611),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_597),
.Y(n_611)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_598),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_602),
.A2(n_603),
.B1(n_609),
.B2(n_610),
.Y(n_608)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_608),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_608),
.Y(n_613)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);


endmodule