module real_jpeg_7019_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_0),
.A2(n_137),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_0),
.A2(n_188),
.B1(n_195),
.B2(n_217),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_0),
.A2(n_217),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_0),
.A2(n_36),
.B1(n_143),
.B2(n_217),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_1),
.A2(n_56),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_1),
.A2(n_56),
.B1(n_175),
.B2(n_396),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_1),
.A2(n_56),
.B1(n_99),
.B2(n_410),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_104),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_104),
.B1(n_141),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_2),
.A2(n_104),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_3),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_95),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_3),
.A2(n_95),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_3),
.A2(n_95),
.B1(n_289),
.B2(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_4),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_174),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_4),
.A2(n_93),
.B1(n_103),
.B2(n_174),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_4),
.A2(n_152),
.B1(n_174),
.B2(n_346),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_5),
.Y(n_206)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_5),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_6),
.Y(n_340)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_6),
.Y(n_347)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_7),
.Y(n_343)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_19)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_14),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_14),
.A2(n_64),
.B1(n_354),
.B2(n_358),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_14),
.A2(n_64),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_14),
.A2(n_64),
.B1(n_312),
.B2(n_449),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_15),
.A2(n_188),
.B1(n_194),
.B2(n_195),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_15),
.A2(n_134),
.B1(n_194),
.B2(n_257),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_15),
.A2(n_194),
.B1(n_344),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_15),
.A2(n_194),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_17),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_17),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_17),
.B(n_183),
.C(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_17),
.B(n_81),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_17),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_17),
.B(n_132),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_17),
.B(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_18),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_18),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_18),
.A2(n_175),
.B1(n_281),
.B2(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_18),
.A2(n_281),
.B1(n_287),
.B2(n_405),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g462 ( 
.A1(n_18),
.A2(n_281),
.B1(n_340),
.B2(n_463),
.Y(n_462)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_538),
.B(n_541),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_155),
.B(n_537),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_147),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_26),
.B(n_147),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_139),
.C(n_144),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_27),
.A2(n_28),
.B1(n_533),
.B2(n_534),
.Y(n_532)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_65),
.C(n_105),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_29),
.B(n_525),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_50),
.B1(n_57),
.B2(n_59),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_30),
.A2(n_57),
.B1(n_59),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_30),
.A2(n_57),
.B1(n_140),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_30),
.A2(n_368),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_30),
.A2(n_40),
.B1(n_412),
.B2(n_437),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_30),
.A2(n_50),
.B1(n_57),
.B2(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_31),
.A2(n_366),
.B(n_367),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_31),
.B(n_369),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_31),
.A2(n_58),
.B(n_540),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_36),
.Y(n_413)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_37),
.Y(n_143)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_37),
.Y(n_463)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_40),
.B(n_169),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_43),
.Y(n_288)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_44),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_44),
.Y(n_374)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_46),
.Y(n_338)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g334 ( 
.A1(n_48),
.A2(n_335),
.A3(n_339),
.B1(n_341),
.B2(n_345),
.Y(n_334)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_57),
.A2(n_437),
.B(n_464),
.Y(n_474)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_58),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_58),
.B(n_462),
.Y(n_461)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_65),
.A2(n_105),
.B1(n_106),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_65),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_65)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_66),
.A2(n_96),
.B1(n_309),
.B2(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_66),
.A2(n_96),
.B1(n_404),
.B2(n_409),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_66),
.A2(n_90),
.B1(n_96),
.B2(n_514),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_81),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_75),
.B2(n_80),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_69),
.Y(n_294)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_70),
.Y(n_298)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_74),
.Y(n_272)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_74),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_74),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g438 ( 
.A1(n_81),
.A2(n_145),
.B1(n_315),
.B2(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_81),
.A2(n_145),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_89),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_85),
.Y(n_401)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_87),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_87),
.Y(n_396)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_88),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_88),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_96),
.B(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_96),
.A2(n_309),
.B(n_314),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_105),
.A2(n_106),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_105),
.B(n_509),
.C(n_512),
.Y(n_520)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_131),
.B(n_133),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_165),
.B(n_170),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_107),
.A2(n_131),
.B1(n_216),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_107),
.A2(n_170),
.B(n_256),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_107),
.A2(n_131),
.B1(n_376),
.B2(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_108),
.B(n_171),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_108),
.A2(n_132),
.B1(n_395),
.B2(n_397),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_108),
.A2(n_132),
.B1(n_397),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_108),
.A2(n_132),
.B1(n_419),
.B2(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_112),
.Y(n_422)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_121),
.A2(n_216),
.B(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_126),
.Y(n_282)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_126),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_126),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_127),
.Y(n_323)
);

BUFx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_128),
.Y(n_280)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_128),
.Y(n_357)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_131),
.A2(n_220),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_133),
.Y(n_453)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_136),
.B(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_139),
.B(n_144),
.Y(n_534)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_145),
.A2(n_264),
.B(n_273),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_145),
.B(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_145),
.A2(n_273),
.B(n_477),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_147),
.B(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_147),
.B(n_539),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_148),
.Y(n_540)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_154),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_531),
.B(n_536),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_503),
.B(n_528),
.Y(n_156)
);

OAI311xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_381),
.A3(n_479),
.B1(n_497),
.C1(n_502),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_328),
.B(n_380),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_300),
.B(n_327),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_250),
.B(n_299),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_223),
.B(n_249),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_185),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_163),
.B(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_178),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_164),
.A2(n_178),
.B1(n_179),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_169),
.A2(n_198),
.B(n_204),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_169),
.A2(n_265),
.B(n_269),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_169),
.B(n_346),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_SL g366 ( 
.A1(n_169),
.A2(n_345),
.B(n_346),
.Y(n_366)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_213),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_214),
.C(n_222),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_198),
.B(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_197),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_198),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_198),
.A2(n_351),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_198),
.A2(n_390),
.B(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_207),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_199),
.A2(n_278),
.B1(n_319),
.B2(n_324),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_199),
.A2(n_353),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_205),
.Y(n_351)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_221),
.B2(n_222),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_239),
.B(n_248),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_238),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_237),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B(n_236),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_277),
.B(n_283),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_246),
.Y(n_248)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_252),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_275),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_262),
.B2(n_263),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_262),
.C(n_275),
.Y(n_301)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx5_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_265),
.Y(n_410)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_268),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI32xp33_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_287),
.A3(n_289),
.B1(n_292),
.B2(n_295),
.Y(n_286)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_301),
.B(n_302),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_326),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_306),
.C(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_316),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_317),
.C(n_318),
.Y(n_360)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_329),
.B(n_330),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_363),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_348),
.B2(n_349),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_334),
.B(n_348),
.Y(n_475)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_360),
.B(n_361),
.C(n_363),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_370),
.B2(n_379),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_364),
.B(n_371),
.C(n_375),
.Y(n_488)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_370),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

INVx6_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_465),
.Y(n_381)
);

A2O1A1Ixp33_ASAP7_75t_SL g497 ( 
.A1(n_382),
.A2(n_465),
.B(n_498),
.C(n_501),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_440),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_383),
.B(n_440),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_416),
.C(n_428),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_384),
.B(n_416),
.CI(n_428),
.CON(n_478),
.SN(n_478)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_402),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_385),
.B(n_403),
.C(n_411),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_386),
.B(n_394),
.Y(n_471)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_411),
.Y(n_402)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_423),
.B2(n_427),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_423),
.Y(n_457)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_423),
.A2(n_427),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_423),
.A2(n_457),
.B(n_460),
.Y(n_506)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_435),
.C(n_438),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_432),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_432),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_435),
.A2(n_436),
.B1(n_438),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_441),
.B(n_444),
.C(n_455),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_455),
.B2(n_456),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_451),
.B(n_454),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_452),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g505 ( 
.A(n_454),
.B(n_506),
.CI(n_507),
.CON(n_505),
.SN(n_505)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_506),
.C(n_507),
.Y(n_527)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_478),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_478),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.C(n_472),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_467),
.A2(n_468),
.B1(n_471),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_471),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.C(n_476),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_473),
.A2(n_474),
.B1(n_476),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_478),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_492),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_481),
.A2(n_499),
.B(n_500),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_489),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.C(n_488),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_495),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_494),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_517),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_516),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_516),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_505),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_511),
.B2(n_515),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_508),
.A2(n_509),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_519),
.C(n_523),
.Y(n_535)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_511),
.Y(n_515)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_517),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_527),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_527),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_535),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);


endmodule