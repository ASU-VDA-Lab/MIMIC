module real_jpeg_6447_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_5),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_21),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_33),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_8),
.B(n_28),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_20),
.B(n_23),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_12),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_14),
.B(n_18),
.Y(n_12)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_17),
.A2(n_40),
.B(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

OR2x4_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_49),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);


endmodule