module fake_netlist_1_11086_n_641 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_641, n_602);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_641;
output n_602;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_63), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_52), .Y(n_75) );
INVx2_ASAP7_75t_SL g76 ( .A(n_19), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_59), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_47), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_40), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_48), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_8), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_5), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_25), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_66), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_37), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_5), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_7), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_10), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_22), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_60), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_49), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_4), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_54), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_35), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_62), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_58), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_55), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_23), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_36), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_51), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_18), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_61), .Y(n_118) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_101), .A2(n_31), .B(n_71), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_88), .A2(n_95), .B1(n_82), .B2(n_83), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_104), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_88), .B(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_74), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_101), .B(n_76), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_102), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_76), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_75), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_108), .B(n_1), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_108), .B(n_2), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_100), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_78), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_114), .B(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_100), .Y(n_144) );
BUFx12f_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_80), .B(n_6), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_92), .B(n_34), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_103), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_105), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_106), .B(n_8), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_121), .B(n_118), .C(n_117), .Y(n_161) );
INVx2_ASAP7_75t_SL g162 ( .A(n_158), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_158), .B(n_118), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_128), .B(n_109), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_132), .B(n_116), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_128), .B(n_117), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_145), .B(n_112), .Y(n_168) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_123), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_134), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_120), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx5_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_137), .B(n_85), .Y(n_174) );
INVxp67_ASAP7_75t_SL g175 ( .A(n_123), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_123), .B(n_85), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_132), .B(n_115), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_135), .A2(n_98), .B1(n_94), .B2(n_111), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_127), .B(n_115), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_147), .B(n_109), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_127), .B(n_93), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_149), .A2(n_110), .B1(n_112), .B2(n_93), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_147), .B(n_90), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_145), .B(n_90), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_120), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_133), .B(n_84), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_124), .B(n_9), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_133), .B(n_110), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_138), .B(n_38), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_144), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g204 ( .A(n_138), .B(n_33), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_141), .B(n_39), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_120), .Y(n_207) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_119), .A2(n_32), .B(n_68), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_129), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_131), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_142), .B(n_9), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_203), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_199), .B(n_157), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_174), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_173), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_212), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_165), .B(n_157), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_162), .B(n_142), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_182), .B(n_152), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_173), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_195), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_162), .B(n_150), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_191), .A2(n_149), .B1(n_136), .B2(n_154), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_198), .B(n_150), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_182), .B(n_152), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_191), .B(n_154), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_167), .B(n_153), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_203), .Y(n_232) );
AND2x6_ASAP7_75t_SL g233 ( .A(n_168), .B(n_155), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_167), .B(n_153), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_173), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_168), .A2(n_122), .B1(n_125), .B2(n_148), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_159), .A2(n_156), .B1(n_151), .B2(n_148), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_187), .B(n_156), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_188), .B(n_151), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_187), .A2(n_139), .B1(n_131), .B2(n_122), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_159), .A2(n_139), .B1(n_125), .B2(n_140), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_196), .B(n_140), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_187), .B(n_140), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_159), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_177), .B(n_119), .Y(n_249) );
AND3x1_ASAP7_75t_L g250 ( .A(n_190), .B(n_11), .C(n_12), .Y(n_250) );
CKINVDCx14_ASAP7_75t_R g251 ( .A(n_168), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_170), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_170), .A2(n_130), .B1(n_120), .B2(n_146), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_163), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_178), .B(n_146), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_178), .A2(n_146), .B1(n_130), .B2(n_120), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_192), .B(n_146), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_170), .A2(n_130), .B1(n_120), .B2(n_146), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_183), .B(n_146), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_166), .A2(n_130), .B1(n_12), .B2(n_13), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_193), .Y(n_264) );
AND2x6_ASAP7_75t_L g265 ( .A(n_189), .B(n_130), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_166), .A2(n_130), .B1(n_13), .B2(n_14), .Y(n_266) );
NOR2x2_ASAP7_75t_L g267 ( .A(n_205), .B(n_11), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
OAI22xp5_ASAP7_75t_SL g269 ( .A1(n_181), .A2(n_202), .B1(n_161), .B2(n_197), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g270 ( .A1(n_251), .A2(n_205), .B1(n_166), .B2(n_180), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_263), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_217), .B(n_181), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_220), .A2(n_192), .B(n_186), .C(n_164), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_249), .A2(n_160), .B(n_179), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_222), .B(n_166), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_180), .B(n_204), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_214), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_225), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_222), .B(n_166), .Y(n_279) );
INVxp67_ASAP7_75t_SL g280 ( .A(n_263), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_254), .B(n_180), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_218), .B(n_205), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_SL g283 ( .A1(n_221), .A2(n_200), .B(n_204), .C(n_210), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_226), .B(n_205), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_226), .B(n_200), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_267), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_225), .Y(n_287) );
O2A1O1Ixp5_ASAP7_75t_L g288 ( .A1(n_231), .A2(n_210), .B(n_172), .C(n_201), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_259), .A2(n_208), .B(n_185), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_228), .B(n_208), .Y(n_290) );
NOR2xp67_ASAP7_75t_L g291 ( .A(n_232), .B(n_17), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_221), .A2(n_201), .B(n_185), .C(n_184), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_264), .B(n_184), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_215), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_241), .B(n_172), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_230), .A2(n_207), .B(n_194), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
BUFx5_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_263), .B(n_207), .Y(n_301) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_230), .A2(n_207), .B(n_194), .Y(n_303) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_250), .B(n_24), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_248), .A2(n_207), .B(n_194), .Y(n_305) );
NOR2xp33_ASAP7_75t_R g306 ( .A(n_233), .B(n_26), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_216), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_225), .B(n_194), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_269), .B(n_27), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_223), .A2(n_171), .B(n_30), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_238), .B(n_29), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_227), .B(n_43), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_229), .A2(n_171), .B(n_45), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_241), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_296), .B(n_235), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_244), .B1(n_261), .B2(n_260), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_299), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_SL g318 ( .A1(n_290), .A2(n_255), .B(n_257), .C(n_242), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_307), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_283), .A2(n_256), .B(n_266), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_272), .A2(n_247), .B(n_236), .C(n_234), .Y(n_322) );
NOR2xp33_ASAP7_75t_SL g323 ( .A(n_277), .B(n_265), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_276), .A2(n_246), .B(n_268), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_286), .A2(n_243), .B1(n_239), .B2(n_252), .Y(n_325) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_271), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_294), .A2(n_262), .B(n_240), .C(n_219), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_272), .B(n_239), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_274), .A2(n_245), .B(n_258), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_302), .B(n_213), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_286), .B(n_245), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_305), .A2(n_258), .B(n_253), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_270), .A2(n_213), .B1(n_237), .B2(n_224), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_312), .A2(n_253), .B(n_265), .C(n_171), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_314), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_306), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_273), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_309), .A2(n_265), .B(n_46), .C(n_50), .Y(n_342) );
AO31x2_ASAP7_75t_L g343 ( .A1(n_289), .A2(n_265), .A3(n_171), .B(n_56), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_336), .A2(n_313), .B(n_310), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_324), .A2(n_305), .B(n_298), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_318), .A2(n_303), .B(n_285), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_343), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_339), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_333), .A2(n_301), .B(n_308), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_330), .A2(n_284), .B(n_282), .Y(n_352) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_335), .A2(n_292), .B(n_287), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_328), .A2(n_279), .B(n_275), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_337), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_340), .A2(n_280), .B(n_311), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_315), .B(n_304), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_322), .A2(n_302), .B(n_271), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_322), .A2(n_271), .B(n_278), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_327), .B(n_278), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_332), .B(n_291), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_343), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_341), .A2(n_300), .B1(n_53), .B2(n_57), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_326), .B(n_44), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_325), .A2(n_64), .B1(n_72), .B2(n_300), .C(n_316), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_317), .Y(n_369) );
AOI21x1_ASAP7_75t_L g370 ( .A1(n_348), .A2(n_334), .B(n_343), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_349), .B(n_338), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_360), .B(n_326), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_356), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_360), .B(n_331), .Y(n_374) );
INVx6_ASAP7_75t_SL g375 ( .A(n_366), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_363), .B(n_342), .C(n_323), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_348), .A2(n_321), .B(n_342), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_349), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_366), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_351), .B(n_321), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_358), .B(n_331), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_351), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_348), .Y(n_388) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_358), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_369), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_362), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_300), .B1(n_365), .B2(n_363), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_300), .B(n_359), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_365), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_300), .B(n_346), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_389), .B(n_357), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_376), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_376), .B(n_357), .Y(n_405) );
AND4x1_ASAP7_75t_L g406 ( .A(n_377), .B(n_361), .C(n_352), .D(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_378), .B(n_357), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_384), .B(n_357), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_399), .A2(n_367), .B1(n_352), .B2(n_353), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_390), .B(n_353), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_392), .B(n_353), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_390), .B(n_345), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_384), .B(n_345), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_388), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_397), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_370), .A2(n_350), .B(n_345), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_381), .B(n_345), .Y(n_422) );
INVx5_ASAP7_75t_SL g423 ( .A(n_375), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_344), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_375), .A2(n_344), .B1(n_350), .B2(n_393), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_386), .B(n_344), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_400), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_391), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_373), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_386), .B(n_344), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
OR2x6_ASAP7_75t_L g441 ( .A(n_382), .B(n_383), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_387), .B(n_382), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_394), .A2(n_383), .A3(n_374), .B(n_385), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_402), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_402), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_383), .B(n_372), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_383), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_372), .B(n_380), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g450 ( .A(n_436), .B(n_371), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_417), .B(n_380), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_430), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_380), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_380), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_410), .B(n_385), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_418), .B(n_374), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_430), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_422), .B(n_398), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_401), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_447), .B(n_398), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_418), .B(n_401), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_419), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_447), .B(n_401), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_430), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_419), .B(n_401), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_414), .B(n_370), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_426), .B(n_375), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_420), .B(n_431), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_431), .B(n_442), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_411), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_426), .B(n_449), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_441), .B(n_443), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_442), .B(n_424), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_427), .B(n_434), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_449), .B(n_429), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_429), .B(n_439), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_445), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
OR2x6_ASAP7_75t_SL g489 ( .A(n_403), .B(n_424), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_439), .B(n_443), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_424), .B(n_409), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_446), .B(n_432), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_428), .B(n_434), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_425), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_427), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_409), .B(n_405), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_432), .B(n_440), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_441), .B(n_434), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_446), .B(n_440), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_433), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_405), .B(n_438), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_415), .B(n_438), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_480), .B(n_415), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_463), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_438), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_485), .B(n_437), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_485), .B(n_437), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_497), .B(n_413), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_497), .B(n_413), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_486), .B(n_403), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_486), .B(n_448), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_452), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_491), .B(n_437), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_491), .B(n_408), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_490), .B(n_448), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_456), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_489), .B(n_435), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_490), .B(n_408), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_453), .B(n_435), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_453), .B(n_435), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_489), .Y(n_528) );
OAI21xp33_ASAP7_75t_L g529 ( .A1(n_473), .A2(n_412), .B(n_441), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_455), .B(n_441), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_455), .B(n_441), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_503), .B(n_425), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_458), .B(n_444), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_503), .B(n_472), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_465), .B(n_425), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_487), .B(n_444), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_504), .B(n_425), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_434), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_462), .B(n_421), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_488), .B(n_427), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_462), .B(n_421), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_504), .B(n_421), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_477), .A2(n_427), .B1(n_421), .B2(n_406), .C(n_423), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_468), .B(n_406), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_484), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_450), .B(n_423), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_468), .B(n_423), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_459), .B(n_423), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_459), .B(n_423), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_528), .B(n_551), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_539), .B(n_457), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_539), .B(n_457), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_548), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_548), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_541), .B(n_474), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_514), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_516), .B(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_541), .B(n_474), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_529), .A2(n_493), .B(n_461), .C(n_470), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_546), .B(n_481), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_522), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_546), .B(n_505), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_550), .B(n_494), .Y(n_569) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_551), .B(n_494), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_505), .B(n_481), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_534), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_520), .B(n_492), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_530), .B(n_499), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_514), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_520), .B(n_500), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_517), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_512), .B(n_482), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_533), .A2(n_481), .B1(n_499), .B2(n_454), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_512), .B(n_502), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_513), .B(n_536), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_515), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_521), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_554), .B(n_513), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_569), .B(n_544), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_575), .Y(n_590) );
NAND2x1_ASAP7_75t_SL g591 ( .A(n_554), .B(n_535), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_566), .A2(n_530), .B1(n_531), .B2(n_538), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_580), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_581), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_569), .B(n_494), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_584), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_587), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_564), .A2(n_493), .B(n_483), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_585), .B(n_523), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_574), .A2(n_525), .B1(n_524), .B2(n_508), .C(n_531), .Y(n_601) );
UNKNOWN g602 ( );
INVx1_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_560), .A2(n_538), .B1(n_535), .B2(n_532), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_571), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_570), .A2(n_554), .B(n_578), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_582), .B(n_523), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_589), .A2(n_565), .B1(n_567), .B2(n_559), .Y(n_609) );
OAI32xp33_ASAP7_75t_L g610 ( .A1(n_606), .A2(n_567), .A3(n_565), .B1(n_537), .B2(n_568), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_601), .A2(n_600), .B1(n_592), .B2(n_604), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_605), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_601), .A2(n_570), .B1(n_561), .B2(n_576), .C(n_579), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_608), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_599), .A2(n_559), .B1(n_562), .B2(n_555), .C(n_556), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_602), .A2(n_540), .B(n_454), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_599), .A2(n_577), .B(n_499), .C(n_537), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_591), .A2(n_562), .B(n_572), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_595), .A2(n_511), .B1(n_510), .B2(n_509), .C(n_542), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g620 ( .A(n_588), .B(n_552), .C(n_553), .D(n_496), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_617), .A2(n_603), .B1(n_598), .B2(n_590), .C(n_593), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_615), .A2(n_555), .A3(n_556), .B1(n_596), .B2(n_584), .C1(n_572), .C2(n_577), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_611), .B(n_553), .C(n_577), .D(n_542), .Y(n_623) );
NAND4xp75_ASAP7_75t_L g624 ( .A(n_609), .B(n_597), .C(n_594), .D(n_532), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_610), .A2(n_607), .B(n_478), .C(n_475), .Y(n_625) );
NAND3xp33_ASAP7_75t_SL g626 ( .A(n_618), .B(n_519), .C(n_479), .Y(n_626) );
AOI222xp33_ASAP7_75t_L g627 ( .A1(n_613), .A2(n_507), .B1(n_527), .B2(n_526), .C1(n_586), .C2(n_563), .Y(n_627) );
OAI211xp5_ASAP7_75t_SL g628 ( .A1(n_622), .A2(n_616), .B(n_619), .C(n_612), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_626), .B(n_620), .Y(n_629) );
NAND4xp75_ASAP7_75t_L g630 ( .A(n_623), .B(n_614), .C(n_526), .D(n_527), .Y(n_630) );
OAI321xp33_ASAP7_75t_L g631 ( .A1(n_625), .A2(n_519), .A3(n_518), .B1(n_586), .B2(n_563), .C(n_464), .Y(n_631) );
NOR5xp2_ASAP7_75t_L g632 ( .A(n_628), .B(n_621), .C(n_624), .D(n_627), .E(n_501), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_629), .B(n_547), .C(n_545), .Y(n_633) );
XOR2x2_ASAP7_75t_L g634 ( .A(n_633), .B(n_630), .Y(n_634) );
NOR2x2_ASAP7_75t_L g635 ( .A(n_632), .B(n_631), .Y(n_635) );
INVxp33_ASAP7_75t_SL g636 ( .A(n_635), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_636), .A2(n_634), .B1(n_543), .B2(n_545), .Y(n_637) );
AOI21xp33_ASAP7_75t_SL g638 ( .A1(n_637), .A2(n_498), .B(n_547), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_638), .A2(n_543), .B(n_549), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_639), .A2(n_549), .B1(n_495), .B2(n_471), .C(n_466), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_640), .A2(n_464), .B1(n_466), .B2(n_471), .Y(n_641) );
endmodule