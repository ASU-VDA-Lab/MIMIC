module real_jpeg_21766_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_334, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_334;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_0),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_96),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_96),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_96),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_1),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_86),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_86),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_86),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_29),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_2),
.A2(n_43),
.B(n_46),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_101),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_80),
.B1(n_81),
.B2(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_2),
.B(n_57),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_2),
.A2(n_31),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_23),
.B1(n_46),
.B2(n_47),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_3),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_4),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_103),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_103),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_103),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_6),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_98),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_98),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_237)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_257)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_11),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_11),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_12),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_92),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_253)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_31),
.A3(n_42),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx3_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_327),
.B(n_330),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_70),
.B(n_326),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_35),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_21),
.B(n_35),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_21),
.B(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_21),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_27),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_24),
.B(n_101),
.CON(n_100),
.SN(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_26),
.A2(n_29),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_26),
.A2(n_29),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_26),
.A2(n_29),
.B(n_33),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_27),
.B(n_31),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_28),
.A2(n_30),
.B1(n_100),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_30),
.B(n_101),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_66),
.C(n_68),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_36),
.A2(n_37),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_49),
.C(n_58),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_38),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_38),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_38),
.A2(n_49),
.B1(n_296),
.B2(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B(n_48),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_45),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_39),
.A2(n_45),
.B1(n_85),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_39),
.A2(n_45),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_39),
.A2(n_45),
.B1(n_155),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_39),
.A2(n_45),
.B1(n_176),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_39),
.A2(n_45),
.B1(n_91),
.B2(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_39),
.A2(n_45),
.B1(n_87),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_39),
.A2(n_45),
.B1(n_230),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_39),
.A2(n_45),
.B1(n_48),
.B2(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_41),
.B(n_53),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_42),
.A2(n_44),
.B(n_101),
.C(n_151),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_45),
.B(n_101),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_47),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_56),
.B(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_51),
.A2(n_57),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_51),
.A2(n_57),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_55),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_52),
.A2(n_55),
.B1(n_97),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_52),
.A2(n_55),
.B1(n_128),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_52),
.A2(n_55),
.B1(n_111),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_52),
.A2(n_55),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_58),
.A2(n_59),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_60),
.A2(n_63),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_60),
.A2(n_63),
.B1(n_109),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_60),
.A2(n_63),
.B1(n_237),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_68),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_319),
.B(n_325),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_288),
.A3(n_311),
.B1(n_317),
.B2(n_318),
.C(n_334),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_267),
.B(n_287),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_243),
.B(n_266),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_134),
.B(n_219),
.C(n_242),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_119),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_76),
.B(n_119),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_104),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_88),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_78),
.B(n_88),
.C(n_104),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_79),
.B(n_84),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_82),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_80),
.A2(n_117),
.B1(n_118),
.B2(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_80),
.A2(n_144),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_80),
.A2(n_81),
.B1(n_147),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_80),
.A2(n_133),
.B1(n_160),
.B2(n_178),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_80),
.A2(n_83),
.B1(n_160),
.B2(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_80),
.A2(n_160),
.B(n_228),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_101),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.C(n_99),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_106),
.B(n_112),
.C(n_113),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.C(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_218),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_213),
.B(n_217),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_199),
.B(n_212),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_180),
.B(n_198),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_168),
.B(n_179),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_156),
.B(n_167),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_148),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_162),
.B(n_166),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_182),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_185),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_201),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_209),
.C(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_221),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_241),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_232),
.C(n_241),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_235),
.C(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_245),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_265),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_258),
.B2(n_259),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_259),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_251),
.C(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_253),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_261),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_262),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_279),
.B(n_282),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_285),
.B2(n_286),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_278),
.C(n_286),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_277),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_290),
.C(n_301),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_290),
.B1(n_291),
.B2(n_316),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_277),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_303),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_303),
.Y(n_318)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_297),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_297),
.A2(n_300),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_305),
.C(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_302),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule