module fake_jpeg_31064_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_10),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

XOR2x1_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_20),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_17),
.B1(n_18),
.B2(n_12),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_13),
.B1(n_14),
.B2(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_19),
.B(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_37),
.B1(n_29),
.B2(n_13),
.Y(n_40)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_41),
.B1(n_42),
.B2(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_25),
.B1(n_28),
.B2(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_48),
.B1(n_43),
.B2(n_39),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_33),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_43),
.B(n_45),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_48),
.A3(n_45),
.B1(n_47),
.B2(n_46),
.C1(n_39),
.C2(n_5),
.Y(n_53)
);

AOI322xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_49),
.A3(n_51),
.B1(n_4),
.B2(n_5),
.C1(n_0),
.C2(n_3),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_52),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_3),
.Y(n_56)
);


endmodule