module fake_jpeg_16561_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_19),
.A2(n_6),
.B(n_1),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_48),
.B(n_33),
.C(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_18),
.B1(n_21),
.B2(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_7),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_9),
.C(n_3),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_11),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_12),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_0),
.C(n_3),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_32),
.C(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_18),
.B1(n_21),
.B2(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_38),
.B1(n_51),
.B2(n_5),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_56),
.B1(n_47),
.B2(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_28),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_77),
.Y(n_97)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_76),
.Y(n_107)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_10),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_11),
.Y(n_84)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_68),
.B(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_103),
.B1(n_59),
.B2(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_32),
.C(n_22),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_92),
.C(n_102),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_22),
.C(n_14),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_95),
.B1(n_64),
.B2(n_86),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_49),
.B(n_40),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_44),
.B1(n_49),
.B2(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_44),
.B1(n_79),
.B2(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_58),
.B1(n_57),
.B2(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_78),
.C(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.C(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_62),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_82),
.B(n_78),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_121),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_106),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_122),
.B(n_127),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_103),
.B1(n_105),
.B2(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_57),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_132),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_97),
.B1(n_120),
.B2(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_58),
.B(n_71),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_129),
.B1(n_116),
.B2(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_97),
.B1(n_102),
.B2(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_91),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_138),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_103),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_108),
.B1(n_89),
.B2(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_111),
.A3(n_103),
.B1(n_92),
.B2(n_101),
.C1(n_88),
.C2(n_96),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_147),
.B(n_133),
.C(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_126),
.B1(n_128),
.B2(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_121),
.B1(n_131),
.B2(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_114),
.C(n_132),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_119),
.C(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_143),
.B1(n_144),
.B2(n_138),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_146),
.C(n_134),
.Y(n_163)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_145),
.B1(n_137),
.B2(n_147),
.C(n_124),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_148),
.C(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_148),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_156),
.C(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_163),
.C(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_154),
.C(n_164),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_174),
.Y(n_178)
);


endmodule