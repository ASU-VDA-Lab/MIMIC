module fake_jpeg_20944_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_15),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_52),
.B1(n_59),
.B2(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_26),
.B1(n_18),
.B2(n_15),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_20),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_51),
.B1(n_58),
.B2(n_56),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_27),
.B1(n_19),
.B2(n_24),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_31),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_14),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_0),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_62),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_69),
.C(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_71),
.B1(n_76),
.B2(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_32),
.B1(n_40),
.B2(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_25),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_45),
.C(n_44),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_57),
.B1(n_1),
.B2(n_3),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_64),
.B(n_61),
.C(n_75),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_43),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_89),
.C(n_78),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_48),
.C(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_5),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_60),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_63),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_103),
.B(n_108),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_78),
.B(n_71),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_71),
.B(n_77),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_88),
.B(n_84),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_67),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_86),
.C(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_63),
.B(n_5),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_96),
.B(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_103),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_122),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_124),
.Y(n_130)
);

FAx1_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_104),
.CI(n_102),
.CON(n_122),
.SN(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_111),
.C(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.C(n_113),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_111),
.C(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_127),
.C(n_132),
.Y(n_137)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_122),
.A3(n_105),
.B1(n_121),
.B2(n_101),
.C(n_10),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_87),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_122),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_138),
.A3(n_87),
.B1(n_10),
.B2(n_7),
.C1(n_8),
.C2(n_11),
.Y(n_139)
);

AO221x1_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_11),
.B1(n_12),
.B2(n_73),
.C(n_6),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_5),
.Y(n_142)
);


endmodule