module real_jpeg_24618_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_8),
.B1(n_38),
.B2(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_38),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_45),
.C(n_47),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_44),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_34),
.C(n_71),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_22),
.C(n_31),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_4),
.B(n_62),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_74),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_53),
.B1(n_68),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_22),
.B1(n_25),
.B2(n_68),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_64)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_35),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_114),
.B1(n_255),
.B2(n_256),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_14),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_113),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_96),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_16),
.B(n_96),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_57),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_27),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_18),
.A2(n_41),
.B1(n_42),
.B2(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_18),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_18),
.A2(n_28),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_24),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_20),
.B(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_24),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_21),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_22),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_23),
.A2(n_104),
.B(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_27),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_28),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_36),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_29),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_29),
.A2(n_36),
.B(n_130),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

OA22x2_ASAP7_75t_SL g73 ( 
.A1(n_33),
.A2(n_34),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_34),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_37),
.A2(n_39),
.B1(n_62),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_37),
.B(n_89),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_50),
.B1(n_55),
.B2(n_110),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_47),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_47),
.B(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_55),
.Y(n_83)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_52),
.B(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_76),
.B2(n_77),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_60),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_65),
.A2(n_109),
.B1(n_119),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_65),
.B(n_171),
.C(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_65),
.A2(n_161),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_65),
.B(n_109),
.C(n_150),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_73),
.B(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_69),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_92),
.B(n_94),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_111),
.C(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_78),
.A2(n_79),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_78),
.A2(n_79),
.B1(n_131),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_123),
.C(n_131),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_83),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_95),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_101),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_100),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_109),
.C(n_111),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_103),
.Y(n_246)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_106),
.A2(n_107),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_106),
.A2(n_107),
.B1(n_184),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_107),
.B(n_178),
.C(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_107),
.B(n_155),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_111),
.A2(n_112),
.B1(n_146),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_111),
.A2(n_112),
.B1(n_129),
.B2(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_112),
.B(n_129),
.C(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_114),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_136),
.B(n_254),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_134),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_116),
.B(n_134),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_117),
.B(n_120),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_122),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_123),
.A2(n_124),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_129),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_157),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_129),
.A2(n_143),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_131),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_249),
.B(n_253),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_174),
.B(n_235),
.C(n_248),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_163),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_139),
.B(n_163),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_149),
.B2(n_162),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_142),
.B(n_148),
.C(n_162),
.Y(n_236)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_154),
.A2(n_155),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_209),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_170),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_165),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_173),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_234),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_193),
.B(n_233),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_190),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_177),
.B(n_190),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_179),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_226),
.B(n_232),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_220),
.B(n_225),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_212),
.B(n_219),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_202),
.B(n_211),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_210),
.Y(n_202)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_244),
.B2(n_245),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_245),
.C(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);


endmodule