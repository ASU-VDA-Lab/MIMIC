module fake_jpeg_26515_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_3),
.Y(n_64)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_42),
.B1(n_34),
.B2(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_40),
.B1(n_35),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_39),
.B1(n_17),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_39),
.C(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_16),
.C(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_6),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_67),
.CON(n_82),
.SN(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_6),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_7),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_59),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_73),
.B1(n_20),
.B2(n_22),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_21),
.B1(n_27),
.B2(n_10),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_8),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_9),
.B(n_30),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_11),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_13),
.C(n_15),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_78),
.C(n_68),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_72),
.B(n_76),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_89),
.B(n_86),
.Y(n_91)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_86),
.C(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_75),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_81),
.B(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_71),
.B(n_80),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_73),
.C(n_90),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_24),
.Y(n_98)
);


endmodule