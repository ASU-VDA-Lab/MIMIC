module fake_jpeg_27111_n_274 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_20;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_24),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_21),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_45),
.Y(n_53)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_42),
.B1(n_48),
.B2(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_34),
.B1(n_28),
.B2(n_32),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_37),
.B1(n_42),
.B2(n_47),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_13),
.B1(n_25),
.B2(n_17),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_34),
.B1(n_32),
.B2(n_25),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_62),
.B1(n_39),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_25),
.B1(n_13),
.B2(n_16),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_49),
.B1(n_59),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_62),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_39),
.CI(n_27),
.CON(n_77),
.SN(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_81),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_64),
.B1(n_57),
.B2(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_49),
.B1(n_55),
.B2(n_13),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_85),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_43),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_92),
.B1(n_80),
.B2(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_101),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_63),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_83),
.B1(n_79),
.B2(n_77),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_57),
.B(n_51),
.C(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_50),
.C(n_56),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_98),
.C(n_65),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_67),
.B1(n_73),
.B2(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_61),
.B1(n_40),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_100),
.B1(n_69),
.B2(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_31),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_31),
.C(n_27),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_25),
.B1(n_13),
.B2(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_73),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_106),
.B(n_117),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_68),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_116),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_86),
.B1(n_101),
.B2(n_93),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_123),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_26),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_82),
.C(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_136),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_134),
.B1(n_143),
.B2(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_86),
.B1(n_103),
.B2(n_101),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_88),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_109),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_114),
.C(n_107),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_156),
.C(n_165),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_116),
.C(n_100),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_141),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_122),
.C(n_109),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_147),
.B1(n_143),
.B2(n_127),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_121),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_10),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_75),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_65),
.C(n_66),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_0),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_97),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_35),
.C(n_29),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_171),
.C(n_165),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_97),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_147),
.B1(n_125),
.B2(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_180),
.B1(n_153),
.B2(n_16),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_131),
.B1(n_128),
.B2(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_131),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_190),
.B(n_12),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_102),
.B1(n_97),
.B2(n_72),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_191),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_174),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_14),
.B1(n_26),
.B2(n_16),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_169),
.B1(n_154),
.B2(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_163),
.B1(n_159),
.B2(n_155),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_192),
.C(n_188),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_180),
.C(n_35),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_160),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_14),
.B(n_26),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_203),
.B1(n_209),
.B2(n_23),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_205),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_202),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_15),
.B1(n_20),
.B2(n_23),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_208),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_15),
.B1(n_20),
.B2(n_23),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_16),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_15),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_185),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_223),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_172),
.B(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_175),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_225),
.C(n_19),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_14),
.B(n_23),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_29),
.C(n_19),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_24),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_24),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_199),
.B1(n_196),
.B2(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_210),
.C(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_220),
.C(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_236),
.C(n_18),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_18),
.B1(n_20),
.B2(n_15),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_224),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_225),
.B(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_242),
.C(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

NOR2x1_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_12),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_22),
.C(n_11),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_12),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_226),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_18),
.C(n_22),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_8),
.C(n_1),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_244),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_234),
.B(n_237),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_256),
.B(n_246),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_9),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_257),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_249),
.C(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_261),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_8),
.C(n_1),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_264),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_256),
.C(n_8),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_0),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_263),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_266),
.B(n_5),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_3),
.C(n_7),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_272),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_3),
.B(n_7),
.Y(n_274)
);


endmodule