module fake_netlist_5_1796_n_1757 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1757);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1757;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1705;
wire n_659;
wire n_1294;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_2),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_32),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_52),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_52),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_62),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_122),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_27),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_97),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_32),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_54),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_19),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_36),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_76),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_34),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_58),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_107),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_17),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_23),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_45),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_26),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_1),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_85),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_45),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_41),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_72),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_117),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_38),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_46),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_88),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_89),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_93),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_22),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_24),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_86),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_90),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_34),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_144),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_96),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_2),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_44),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_44),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_28),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_160),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_73),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_75),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_53),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_74),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_101),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_113),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_47),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_69),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_61),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_40),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_12),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_31),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_25),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_55),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_99),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_6),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_87),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_66),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_29),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_57),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_46),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_41),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_138),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_33),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_81),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_94),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_130),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_134),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_38),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_112),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_42),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_18),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_4),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_33),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_79),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_106),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_71),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_43),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_115),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_145),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_237),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_177),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_198),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_177),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_201),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_202),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_167),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_205),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_208),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_207),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_177),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_213),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_174),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_221),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_224),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_174),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_177),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_239),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_177),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_241),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_247),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_249),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_181),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_245),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_258),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_237),
.B(n_0),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_166),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_245),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_245),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_245),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_204),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_204),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_1),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_251),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_303),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_252),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_193),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_255),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_297),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_256),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_263),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_214),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_293),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_232),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_264),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_184),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_265),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_270),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_273),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_274),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_279),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_232),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_197),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_194),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_174),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_275),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_242),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_184),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_234),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_234),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_283),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_176),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_299),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_299),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_199),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_162),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_276),
.B(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_324),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_326),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_162),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_322),
.B(n_165),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_352),
.B(n_163),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_329),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_275),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_344),
.B(n_359),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_228),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_345),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_350),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_331),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_371),
.B(n_194),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_334),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_347),
.B(n_356),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_334),
.B(n_185),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_333),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_381),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_335),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_392),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_360),
.B(n_163),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_362),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_360),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_336),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_R g453 ( 
.A(n_379),
.B(n_164),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_164),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_328),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_334),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_337),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_368),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_339),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_341),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_383),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_348),
.B(n_244),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_342),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_165),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_343),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_337),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_357),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_361),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_363),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_392),
.B1(n_364),
.B2(n_200),
.Y(n_475)
);

OAI221xp5_ASAP7_75t_L g476 ( 
.A1(n_442),
.A2(n_200),
.B1(n_169),
.B2(n_227),
.C(n_250),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_470),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_418),
.Y(n_478)
);

NOR2x1p5_ASAP7_75t_L g479 ( 
.A(n_402),
.B(n_300),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_366),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_412),
.B(n_170),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_445),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_367),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_450),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_170),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_450),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_428),
.B(n_373),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_418),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_448),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_448),
.B(n_375),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_376),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_463),
.B(n_464),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_427),
.B(n_377),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_374),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_407),
.B(n_378),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_421),
.B(n_374),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_380),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_470),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_421),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_407),
.B(n_419),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_449),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_425),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_425),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_470),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_424),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_421),
.B(n_372),
.C(n_209),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_403),
.B(n_370),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_449),
.B(n_291),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_454),
.B(n_318),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_454),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_463),
.B(n_194),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_466),
.A2(n_300),
.B1(n_168),
.B2(n_212),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g536 ( 
.A(n_405),
.B(n_211),
.Y(n_536)
);

BUFx8_ASAP7_75t_SL g537 ( 
.A(n_456),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_SL g538 ( 
.A(n_438),
.B(n_172),
.Y(n_538)
);

HB1xp67_ASAP7_75t_SL g539 ( 
.A(n_441),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_440),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_387),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_405),
.B(n_178),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_415),
.B(n_211),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_431),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

AND3x2_ASAP7_75t_L g547 ( 
.A(n_441),
.B(n_219),
.C(n_218),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_422),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_423),
.B(n_387),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_423),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_426),
.A2(n_271),
.B1(n_222),
.B2(n_233),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_410),
.B(n_383),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_429),
.B(n_388),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_429),
.A2(n_173),
.B1(n_259),
.B2(n_284),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_430),
.B(n_388),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_420),
.B(n_210),
.C(n_203),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_445),
.B(n_196),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_434),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_446),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_424),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_444),
.B(n_319),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_447),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_409),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_435),
.B(n_437),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_452),
.A2(n_225),
.B1(n_243),
.B2(n_235),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_437),
.B(n_389),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_440),
.B(n_206),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_461),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_462),
.B(n_253),
.C(n_240),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_465),
.B(n_196),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_473),
.B(n_196),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_446),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_451),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_409),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_467),
.B(n_383),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_471),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_166),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_401),
.B(n_218),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_433),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_451),
.B(n_389),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_433),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_443),
.B(n_175),
.Y(n_595)
);

INVx6_ASAP7_75t_L g596 ( 
.A(n_433),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_455),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_440),
.Y(n_598)
);

AO21x2_ASAP7_75t_L g599 ( 
.A1(n_443),
.A2(n_217),
.B(n_215),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_455),
.A2(n_246),
.B1(n_257),
.B2(n_260),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_459),
.B(n_383),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_459),
.B(n_399),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_460),
.B(n_219),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_468),
.B(n_321),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_468),
.B(n_399),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_433),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_457),
.B(n_226),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_457),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_469),
.B(n_242),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_458),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_458),
.B(n_231),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_458),
.B(n_390),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_458),
.B(n_236),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_469),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_469),
.B(n_238),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_469),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_401),
.B(n_175),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_401),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_514),
.B(n_404),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_512),
.B(n_330),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_404),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_507),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_474),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_404),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_577),
.B(n_306),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_485),
.B(n_408),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_532),
.B(n_408),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_532),
.B(n_408),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_529),
.B(n_416),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_489),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_531),
.B(n_506),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_480),
.B(n_416),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_474),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_480),
.B(n_242),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_489),
.B(n_174),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_480),
.B(n_416),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_536),
.B(n_242),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_489),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_505),
.B(n_494),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_505),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_483),
.B(n_417),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_498),
.B(n_417),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_536),
.A2(n_353),
.B1(n_346),
.B2(n_308),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_502),
.B(n_417),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_487),
.B(n_272),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_540),
.B(n_277),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_602),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_602),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_560),
.B(n_278),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_494),
.B(n_302),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_507),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_611),
.B(n_242),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_482),
.B(n_307),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_492),
.A2(n_384),
.B(n_337),
.C(n_310),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_611),
.B(n_254),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_606),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_495),
.B(n_254),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_491),
.B(n_179),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_521),
.B(n_179),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_598),
.B(n_254),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_476),
.A2(n_312),
.B1(n_267),
.B2(n_191),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_609),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_475),
.A2(n_180),
.B1(n_182),
.B2(n_290),
.Y(n_669)
);

BUFx4_ASAP7_75t_L g670 ( 
.A(n_539),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_545),
.B(n_254),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_545),
.B(n_254),
.Y(n_672)
);

AOI221xp5_ASAP7_75t_L g673 ( 
.A1(n_538),
.A2(n_171),
.B1(n_186),
.B2(n_188),
.C(n_189),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_516),
.B(n_232),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_510),
.A2(n_171),
.B1(n_288),
.B2(n_186),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_500),
.B(n_320),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_489),
.B(n_174),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_524),
.B(n_320),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_497),
.B(n_573),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_609),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_489),
.A2(n_320),
.B1(n_174),
.B2(n_286),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_541),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_528),
.B(n_174),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_543),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_489),
.B(n_576),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_541),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_543),
.B(n_180),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_541),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_559),
.B(n_285),
.C(n_282),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_610),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_501),
.B(n_182),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_527),
.B(n_183),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_534),
.B(n_183),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_546),
.B(n_187),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_567),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_591),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_488),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_548),
.A2(n_604),
.B(n_551),
.C(n_550),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_567),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_579),
.B(n_220),
.C(n_281),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_528),
.B(n_174),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_484),
.B(n_187),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_479),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_484),
.B(n_190),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_556),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_503),
.B(n_190),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_195),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_504),
.B(n_561),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_519),
.A2(n_384),
.B(n_290),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_580),
.B(n_582),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_504),
.B(n_195),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_SL g714 ( 
.A(n_481),
.B(n_305),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_561),
.B(n_305),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_569),
.B(n_581),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_569),
.B(n_309),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_612),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_528),
.B(n_311),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_519),
.A2(n_384),
.B(n_316),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_576),
.B(n_311),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_486),
.B(n_188),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_584),
.B(n_316),
.Y(n_723)
);

OAI221xp5_ASAP7_75t_L g724 ( 
.A1(n_552),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.C(n_248),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_570),
.B(n_317),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_547),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_516),
.B(n_396),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_522),
.B(n_261),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_538),
.A2(n_262),
.B1(n_266),
.B2(n_269),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_517),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_590),
.A2(n_280),
.B1(n_189),
.B2(n_294),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_612),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_390),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_549),
.A2(n_298),
.B(n_286),
.C(n_287),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_585),
.B(n_396),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_597),
.B(n_394),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_597),
.B(n_393),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_613),
.B(n_391),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_517),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_599),
.A2(n_296),
.B1(n_315),
.B2(n_314),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_490),
.B(n_296),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_556),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_533),
.B(n_192),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_570),
.B(n_294),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_570),
.B(n_391),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_558),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_558),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_558),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_593),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_481),
.B(n_315),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_562),
.B(n_314),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_593),
.B(n_80),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_555),
.B(n_313),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_588),
.B(n_313),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_593),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_599),
.A2(n_301),
.B1(n_298),
.B2(n_292),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_587),
.B(n_301),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_587),
.B(n_292),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

AO22x1_ASAP7_75t_L g760 ( 
.A1(n_601),
.A2(n_289),
.B1(n_288),
.B2(n_287),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_599),
.A2(n_289),
.B1(n_192),
.B2(n_7),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_496),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_549),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_158),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_621),
.A2(n_156),
.B1(n_155),
.B2(n_153),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_572),
.B(n_148),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_574),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_568),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_574),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_614),
.B(n_146),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_136),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_600),
.B(n_8),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_135),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_526),
.B(n_10),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_478),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_496),
.B(n_129),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_595),
.B(n_11),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_576),
.B(n_126),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_591),
.B(n_120),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_589),
.B(n_15),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_535),
.A2(n_116),
.B1(n_105),
.B2(n_103),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_622),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_509),
.B(n_15),
.Y(n_784)
);

O2A1O1Ixp5_ASAP7_75t_L g785 ( 
.A1(n_519),
.A2(n_102),
.B(n_100),
.C(n_98),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_635),
.B(n_607),
.Y(n_787)
);

BUFx8_ASAP7_75t_SL g788 ( 
.A(n_670),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_720),
.A2(n_509),
.B(n_511),
.Y(n_789)
);

AND2x4_ASAP7_75t_SL g790 ( 
.A(n_624),
.B(n_537),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_686),
.A2(n_509),
.B(n_511),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_627),
.B(n_589),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_680),
.A2(n_605),
.B1(n_603),
.B2(n_544),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_685),
.B(n_486),
.Y(n_794)
);

AND2x4_ASAP7_75t_SL g795 ( 
.A(n_637),
.B(n_537),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_680),
.A2(n_557),
.B1(n_619),
.B2(n_617),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_477),
.Y(n_797)
);

NOR2x2_ASAP7_75t_L g798 ( 
.A(n_629),
.B(n_563),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_628),
.A2(n_511),
.B(n_615),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_701),
.C(n_696),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_663),
.B(n_594),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_631),
.A2(n_496),
.B(n_518),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_651),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_630),
.A2(n_608),
.B(n_620),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_632),
.A2(n_496),
.B(n_518),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_634),
.A2(n_496),
.B(n_518),
.Y(n_806)
);

OAI21xp33_ASAP7_75t_L g807 ( 
.A1(n_688),
.A2(n_499),
.B(n_478),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_634),
.A2(n_640),
.B(n_636),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_699),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_663),
.B(n_594),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_673),
.B(n_499),
.C(n_583),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_634),
.A2(n_518),
.B(n_592),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_638),
.A2(n_518),
.B1(n_571),
.B2(n_575),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_649),
.B(n_571),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_SL g816 ( 
.A1(n_641),
.A2(n_493),
.B(n_508),
.C(n_583),
.Y(n_816)
);

NAND2x1_ASAP7_75t_L g817 ( 
.A(n_762),
.B(n_596),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_638),
.A2(n_575),
.B1(n_493),
.B2(n_553),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_684),
.A2(n_554),
.B(n_508),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_634),
.A2(n_586),
.B(n_520),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_683),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_687),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_739),
.B(n_563),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_689),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_645),
.A2(n_586),
.B(n_520),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_633),
.A2(n_586),
.B(n_520),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_668),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_623),
.A2(n_525),
.B(n_592),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_741),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_625),
.A2(n_525),
.B(n_592),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_657),
.A2(n_660),
.B(n_684),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_641),
.A2(n_542),
.B(n_553),
.C(n_554),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_646),
.A2(n_525),
.B(n_530),
.Y(n_833)
);

CKINVDCx8_ASAP7_75t_R g834 ( 
.A(n_629),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_707),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_744),
.A2(n_578),
.B(n_564),
.C(n_542),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_629),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_648),
.A2(n_530),
.B(n_565),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_742),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_643),
.A2(n_596),
.B1(n_591),
.B2(n_530),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_688),
.B(n_565),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_761),
.A2(n_643),
.B1(n_749),
.B2(n_746),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_626),
.B(n_565),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_676),
.B(n_578),
.C(n_564),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_656),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_764),
.A2(n_745),
.B(n_679),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_710),
.B(n_523),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_657),
.A2(n_660),
.B(n_703),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_755),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_642),
.B(n_477),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_596),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_716),
.B(n_763),
.Y(n_852)
);

OA21x2_ASAP7_75t_L g853 ( 
.A1(n_703),
.A2(n_513),
.B(n_523),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_727),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_712),
.A2(n_596),
.B1(n_591),
.B2(n_618),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_767),
.B(n_513),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_769),
.B(n_477),
.Y(n_857)
);

NOR2x1_ASAP7_75t_L g858 ( 
.A(n_712),
.B(n_618),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_758),
.B(n_477),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_681),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_761),
.A2(n_566),
.B1(n_591),
.B2(n_91),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_642),
.B(n_566),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_675),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_777),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_762),
.A2(n_83),
.B(n_68),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_698),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_744),
.A2(n_22),
.B(n_23),
.C(n_28),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_753),
.B(n_29),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_747),
.B(n_35),
.Y(n_870)
);

AND2x2_ASAP7_75t_SL g871 ( 
.A(n_682),
.B(n_772),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_748),
.B(n_37),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_762),
.A2(n_63),
.B(n_49),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_753),
.B(n_754),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_762),
.A2(n_48),
.B(n_49),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_642),
.B(n_48),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_771),
.A2(n_50),
.B(n_51),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_718),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_732),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_773),
.A2(n_50),
.B(n_51),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_781),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_759),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_738),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_750),
.B(n_57),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_754),
.B(n_54),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_757),
.B(n_55),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_700),
.A2(n_757),
.B(n_725),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_667),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_642),
.B(n_752),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_639),
.A2(n_678),
.B(n_719),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_752),
.A2(n_664),
.B1(n_692),
.B2(n_719),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_733),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_637),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_766),
.B(n_682),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_652),
.B(n_653),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_772),
.A2(n_751),
.B(n_743),
.C(n_664),
.Y(n_896)
);

NOR2x1p5_ASAP7_75t_L g897 ( 
.A(n_702),
.B(n_661),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_674),
.B(n_672),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_725),
.A2(n_783),
.B(n_780),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_705),
.B(n_726),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_775),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_728),
.B(n_751),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_743),
.B(n_760),
.C(n_728),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_671),
.B(n_672),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_774),
.B(n_697),
.Y(n_905)
);

AOI22x1_ASAP7_75t_L g906 ( 
.A1(n_722),
.A2(n_711),
.B1(n_671),
.B2(n_665),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_650),
.A2(n_654),
.B(n_655),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_704),
.B(n_717),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_721),
.A2(n_778),
.B(n_776),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_740),
.A2(n_756),
.B(n_692),
.C(n_666),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_666),
.B(n_756),
.C(n_740),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_706),
.A2(n_723),
.B1(n_715),
.B2(n_713),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_734),
.A2(n_784),
.B(n_785),
.C(n_729),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_708),
.B(n_709),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_658),
.B(n_693),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_778),
.A2(n_770),
.B(n_665),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_694),
.B(n_695),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_735),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_736),
.Y(n_919)
);

AOI21xp33_ASAP7_75t_L g920 ( 
.A1(n_669),
.A2(n_724),
.B(n_690),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_765),
.A2(n_784),
.B1(n_782),
.B2(n_770),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_737),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_779),
.A2(n_697),
.B(n_662),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_677),
.A2(n_731),
.B1(n_697),
.B2(n_659),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_697),
.A2(n_480),
.B1(n_485),
.B2(n_635),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_768),
.A2(n_480),
.B1(n_485),
.B2(n_635),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_635),
.B(n_510),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_635),
.A2(n_480),
.B(n_442),
.C(n_680),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_680),
.A2(n_480),
.B1(n_635),
.B2(n_485),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_696),
.B(n_701),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_772),
.A2(n_480),
.B(n_442),
.C(n_761),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_699),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_635),
.B(n_510),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_699),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_762),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_699),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_643),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_635),
.A2(n_480),
.B1(n_485),
.B2(n_483),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_699),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_772),
.A2(n_480),
.B(n_442),
.C(n_761),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_638),
.A2(n_641),
.B(n_657),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_668),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_627),
.B(n_626),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_668),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_635),
.B(n_510),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_772),
.A2(n_480),
.B(n_442),
.C(n_761),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_699),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_635),
.B(n_480),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_644),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_635),
.B(n_514),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_644),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_699),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_684),
.A2(n_703),
.B(n_679),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_635),
.B(n_514),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_668),
.Y(n_962)
);

OAI21xp33_ASAP7_75t_L g963 ( 
.A1(n_688),
.A2(n_464),
.B(n_442),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_720),
.A2(n_686),
.B(n_519),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_628),
.A2(n_480),
.B(n_630),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_684),
.A2(n_703),
.B(n_679),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_929),
.A2(n_874),
.B(n_965),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_819),
.A2(n_791),
.B(n_802),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_953),
.B(n_961),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_805),
.A2(n_966),
.B(n_959),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_830),
.B(n_828),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_789),
.A2(n_935),
.B(n_927),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_874),
.A2(n_902),
.B(n_896),
.C(n_928),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_893),
.B(n_797),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_902),
.A2(n_934),
.B(n_928),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_896),
.A2(n_934),
.B(n_948),
.C(n_910),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_948),
.B(n_914),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_954),
.A2(n_958),
.B(n_955),
.Y(n_978)
);

AOI21x1_ASAP7_75t_SL g979 ( 
.A1(n_859),
.A2(n_886),
.B(n_908),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_914),
.B(n_963),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_960),
.A2(n_964),
.B(n_951),
.Y(n_981)
);

OA21x2_ASAP7_75t_L g982 ( 
.A1(n_887),
.A2(n_848),
.B(n_831),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_951),
.A2(n_890),
.B(n_894),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_809),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_940),
.A2(n_930),
.B(n_913),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_883),
.B(n_852),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_946),
.B(n_900),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_892),
.B(n_871),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_894),
.A2(n_799),
.B(n_909),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_833),
.A2(n_838),
.B(n_836),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_822),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_871),
.A2(n_911),
.B1(n_885),
.B2(n_869),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_932),
.B(n_942),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_804),
.A2(n_899),
.B(n_913),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_923),
.A2(n_825),
.B(n_826),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_932),
.B(n_942),
.Y(n_996)
);

OAI21x1_ASAP7_75t_SL g997 ( 
.A1(n_868),
.A2(n_877),
.B(n_880),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_925),
.A2(n_921),
.B(n_916),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_793),
.A2(n_904),
.B(n_891),
.Y(n_999)
);

AO31x2_ASAP7_75t_L g1000 ( 
.A1(n_910),
.A2(n_949),
.A3(n_885),
.B(n_869),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_938),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_787),
.A2(n_808),
.B(n_846),
.Y(n_1002)
);

AND3x4_ASAP7_75t_L g1003 ( 
.A(n_800),
.B(n_903),
.C(n_933),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_813),
.A2(n_806),
.B(n_820),
.Y(n_1004)
);

CKINVDCx11_ASAP7_75t_R g1005 ( 
.A(n_810),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_801),
.A2(n_811),
.B(n_907),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_SL g1007 ( 
.A1(n_842),
.A2(n_906),
.B(n_857),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_950),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_949),
.A2(n_889),
.B1(n_926),
.B2(n_841),
.Y(n_1009)
);

AO31x2_ASAP7_75t_L g1010 ( 
.A1(n_796),
.A2(n_862),
.A3(n_818),
.B(n_924),
.Y(n_1010)
);

AO31x2_ASAP7_75t_L g1011 ( 
.A1(n_841),
.A2(n_912),
.A3(n_814),
.B(n_865),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_824),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_938),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_844),
.A2(n_812),
.B(n_917),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_854),
.B(n_881),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_SL g1016 ( 
.A(n_893),
.B(n_834),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_853),
.A2(n_863),
.B(n_817),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_915),
.A2(n_847),
.B(n_920),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_792),
.B(n_794),
.Y(n_1019)
);

AO21x1_ASAP7_75t_L g1020 ( 
.A1(n_903),
.A2(n_876),
.B(n_905),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_797),
.B(n_889),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_856),
.A2(n_858),
.B(n_850),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_815),
.A2(n_816),
.B(n_919),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_898),
.A2(n_839),
.B(n_849),
.C(n_835),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_807),
.A2(n_816),
.B(n_855),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_L g1026 ( 
.A1(n_895),
.A2(n_800),
.B1(n_875),
.B2(n_864),
.C(n_922),
.Y(n_1026)
);

O2A1O1Ixp5_ASAP7_75t_L g1027 ( 
.A1(n_870),
.A2(n_872),
.B(n_861),
.C(n_843),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_SL g1028 ( 
.A1(n_866),
.A2(n_873),
.B(n_840),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_946),
.B(n_900),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_829),
.A2(n_794),
.B(n_931),
.Y(n_1030)
);

OAI22x1_ASAP7_75t_L g1031 ( 
.A1(n_837),
.A2(n_897),
.B1(n_957),
.B2(n_941),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_888),
.A2(n_962),
.B(n_878),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_827),
.A2(n_879),
.B(n_947),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_937),
.A2(n_843),
.B(n_918),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_786),
.A2(n_803),
.B(n_956),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_937),
.A2(n_851),
.B(n_939),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_939),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_941),
.B(n_957),
.C(n_884),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_952),
.B(n_845),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_851),
.A2(n_945),
.B(n_882),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_860),
.A2(n_867),
.B(n_901),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_845),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_936),
.B(n_792),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_795),
.B(n_790),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_823),
.A2(n_798),
.B(n_788),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_809),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_953),
.B(n_961),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_819),
.A2(n_791),
.B(n_802),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_854),
.B(n_928),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_797),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_871),
.A2(n_911),
.B1(n_874),
.B2(n_902),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_953),
.B(n_961),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_809),
.B(n_933),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_874),
.B(n_928),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_797),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_809),
.B(n_933),
.Y(n_1056)
);

AO31x2_ASAP7_75t_L g1057 ( 
.A1(n_943),
.A2(n_913),
.A3(n_921),
.B(n_940),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_953),
.B(n_961),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_819),
.A2(n_791),
.B(n_802),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_874),
.B(n_928),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_902),
.B(n_928),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_854),
.B(n_928),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_902),
.B(n_928),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_953),
.B(n_961),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_854),
.B(n_928),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_953),
.B(n_961),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_936),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_797),
.Y(n_1068)
);

INVx6_ASAP7_75t_L g1069 ( 
.A(n_810),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_929),
.A2(n_480),
.B(n_874),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_789),
.A2(n_964),
.B(n_935),
.Y(n_1071)
);

BUFx2_ASAP7_75t_SL g1072 ( 
.A(n_809),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_953),
.B(n_961),
.Y(n_1073)
);

INVx8_ASAP7_75t_L g1074 ( 
.A(n_810),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_953),
.B(n_961),
.Y(n_1075)
);

NAND2x1p5_ASAP7_75t_L g1076 ( 
.A(n_893),
.B(n_797),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_927),
.A2(n_944),
.B(n_935),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_950),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_797),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_819),
.A2(n_791),
.B(n_802),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_821),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_854),
.B(n_928),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_789),
.A2(n_964),
.B(n_935),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_874),
.A2(n_902),
.B1(n_934),
.B2(n_928),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_809),
.Y(n_1085)
);

NAND2x1_ASAP7_75t_L g1086 ( 
.A(n_939),
.B(n_762),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_929),
.A2(n_480),
.B(n_874),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_874),
.A2(n_902),
.B(n_896),
.C(n_928),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_854),
.B(n_928),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_874),
.A2(n_902),
.B(n_896),
.C(n_928),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_927),
.A2(n_944),
.B(n_935),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_821),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_809),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_SL g1094 ( 
.A1(n_910),
.A2(n_896),
.B1(n_963),
.B2(n_942),
.C(n_949),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_797),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_874),
.A2(n_902),
.B(n_928),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_965),
.A2(n_887),
.B(n_848),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_902),
.B(n_928),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_874),
.B(n_928),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_953),
.B(n_961),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_896),
.A2(n_932),
.B(n_949),
.C(n_942),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_874),
.B(n_928),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_874),
.B(n_928),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_953),
.B(n_961),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_854),
.B(n_928),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_938),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_946),
.B(n_627),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_977),
.B(n_1061),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1054),
.A2(n_1103),
.B1(n_1099),
.B2(n_1102),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1093),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1053),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_1005),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_991),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_L g1115 ( 
.A(n_969),
.B(n_1047),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1012),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_1008),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1072),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1078),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1054),
.A2(n_1060),
.B1(n_1099),
.B2(n_1103),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1084),
.A2(n_1060),
.B1(n_1102),
.B2(n_1104),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1065),
.B(n_1082),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1107),
.B(n_987),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1052),
.B(n_1058),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1081),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1079),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1089),
.B(n_1105),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1107),
.B(n_987),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1064),
.A2(n_1075),
.B1(n_1066),
.B2(n_1073),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1053),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_984),
.B(n_1046),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1096),
.A2(n_975),
.B1(n_1051),
.B2(n_992),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1053),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1063),
.B(n_1098),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1001),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1100),
.B(n_1013),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1092),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1029),
.B(n_1050),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1017),
.A2(n_1004),
.B(n_970),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1056),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_973),
.A2(n_1090),
.B(n_1088),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1033),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1051),
.A2(n_992),
.B1(n_976),
.B2(n_980),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1001),
.Y(n_1144)
);

INVx3_ASAP7_75t_SL g1145 ( 
.A(n_1056),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

OAI31xp33_ASAP7_75t_L g1147 ( 
.A1(n_1009),
.A2(n_1038),
.A3(n_1030),
.B(n_986),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1067),
.B(n_988),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1029),
.B(n_1050),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1079),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1039),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1079),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1003),
.A2(n_993),
.B1(n_996),
.B2(n_1070),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1015),
.B(n_1106),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1056),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1003),
.A2(n_1019),
.B1(n_1026),
.B2(n_1043),
.Y(n_1156)
);

BUFx4_ASAP7_75t_SL g1157 ( 
.A(n_1074),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_1055),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1032),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1055),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1018),
.B(n_1094),
.Y(n_1161)
);

OAI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1042),
.A2(n_1106),
.B(n_1026),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1085),
.B(n_1031),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1035),
.B(n_1095),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1055),
.B(n_1068),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1074),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_1095),
.B(n_1037),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1055),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1024),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_1068),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_967),
.A2(n_1101),
.B(n_999),
.C(n_985),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1068),
.B(n_1037),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1000),
.B(n_1014),
.Y(n_1173)
);

OAI321xp33_ASAP7_75t_L g1174 ( 
.A1(n_998),
.A2(n_1087),
.A3(n_1101),
.B1(n_1071),
.B2(n_972),
.C(n_1083),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1068),
.B(n_1016),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_978),
.A2(n_1091),
.B(n_1077),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1000),
.B(n_1006),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1040),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1069),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1040),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1069),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1000),
.B(n_1006),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1020),
.A2(n_1044),
.B1(n_1069),
.B2(n_1021),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1000),
.B(n_1045),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_974),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1036),
.B(n_1034),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_1086),
.B(n_1036),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1074),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_982),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_982),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1077),
.A2(n_1091),
.B(n_989),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1034),
.B(n_1057),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_974),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1076),
.A2(n_1097),
.B1(n_994),
.B2(n_981),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1057),
.B(n_1011),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1076),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1011),
.B(n_1057),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1027),
.B(n_983),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1057),
.B(n_1011),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_997),
.A2(n_1027),
.B(n_1007),
.C(n_1025),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1022),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_989),
.A2(n_981),
.B(n_1002),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1002),
.A2(n_983),
.B(n_1097),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_994),
.B(n_1010),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_979),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1028),
.A2(n_1023),
.B(n_1010),
.C(n_990),
.Y(n_1206)
);

INVx6_ASAP7_75t_SL g1207 ( 
.A(n_1023),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_995),
.A2(n_971),
.B(n_1048),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1010),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_1010),
.B(n_968),
.Y(n_1210)
);

INVx3_ASAP7_75t_SL g1211 ( 
.A(n_1059),
.Y(n_1211)
);

OR2x6_ASAP7_75t_L g1212 ( 
.A(n_1080),
.B(n_1072),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1107),
.B(n_987),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1001),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_874),
.B1(n_902),
.B2(n_510),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1067),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_969),
.B(n_1047),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1093),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1001),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1054),
.A2(n_874),
.B1(n_902),
.B2(n_911),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1054),
.A2(n_874),
.B(n_902),
.C(n_1060),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1072),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1067),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1107),
.B(n_987),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_969),
.B(n_1047),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1084),
.A2(n_977),
.B1(n_1060),
.B2(n_1054),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1013),
.Y(n_1228)
);

BUFx4_ASAP7_75t_SL g1229 ( 
.A(n_1053),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_991),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1093),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1013),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1055),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1017),
.A2(n_1004),
.B(n_970),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1055),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_969),
.B(n_1047),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_969),
.B(n_1047),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_874),
.B(n_902),
.C(n_1060),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1001),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1107),
.B(n_987),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1093),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1167),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1113),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1215),
.A2(n_1120),
.B1(n_1156),
.B2(n_1121),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1144),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1125),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1137),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1157),
.Y(n_1248)
);

AO21x1_ASAP7_75t_L g1249 ( 
.A1(n_1143),
.A2(n_1171),
.B(n_1200),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1114),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1198),
.A2(n_1208),
.B(n_1203),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1221),
.A2(n_1238),
.B1(n_1217),
.B2(n_1236),
.Y(n_1252)
);

INVx3_ASAP7_75t_SL g1253 ( 
.A(n_1118),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_SL g1254 ( 
.A(n_1110),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1139),
.A2(n_1234),
.B(n_1208),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1178),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1154),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1124),
.A2(n_1226),
.B1(n_1237),
.B2(n_1236),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1203),
.A2(n_1194),
.B(n_1176),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.Y(n_1260)
);

INVx5_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1141),
.A2(n_1129),
.B1(n_1184),
.B2(n_1148),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1144),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1220),
.A2(n_1109),
.B1(n_1227),
.B2(n_1115),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1230),
.Y(n_1265)
);

BUFx4f_ASAP7_75t_SL g1266 ( 
.A(n_1117),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1214),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1170),
.B(n_1164),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1214),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1170),
.B(n_1111),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1167),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1170),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1216),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1224),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1207),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1228),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1157),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1151),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_SL g1279 ( 
.A(n_1145),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1219),
.Y(n_1280)
);

AO21x1_ASAP7_75t_L g1281 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1227),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1132),
.A2(n_1153),
.B1(n_1147),
.B2(n_1134),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1124),
.A2(n_1237),
.B1(n_1217),
.B2(n_1226),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1219),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1202),
.A2(n_1191),
.B(n_1206),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1222),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1132),
.B(n_1209),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1206),
.A2(n_1146),
.B(n_1159),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1135),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1174),
.A2(n_1192),
.B(n_1182),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1232),
.Y(n_1292)
);

BUFx2_ASAP7_75t_R g1293 ( 
.A(n_1166),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_1170),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1126),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1108),
.A2(n_1183),
.B1(n_1145),
.B2(n_1119),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1131),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1239),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_1112),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1136),
.A2(n_1122),
.B1(n_1127),
.B2(n_1223),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1189),
.A2(n_1239),
.B1(n_1162),
.B2(n_1140),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1180),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1142),
.A2(n_1187),
.B(n_1201),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1165),
.Y(n_1304)
);

INVx6_ASAP7_75t_SL g1305 ( 
.A(n_1123),
.Y(n_1305)
);

BUFx2_ASAP7_75t_SL g1306 ( 
.A(n_1218),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1130),
.B(n_1155),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1207),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1186),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1186),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1126),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1177),
.A2(n_1182),
.B(n_1195),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1212),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1205),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1229),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1173),
.B(n_1177),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1205),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1172),
.Y(n_1318)
);

AOI21xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1231),
.A2(n_1241),
.B(n_1133),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1190),
.Y(n_1320)
);

BUFx8_ASAP7_75t_L g1321 ( 
.A(n_1168),
.Y(n_1321)
);

AO21x1_ASAP7_75t_L g1322 ( 
.A1(n_1161),
.A2(n_1195),
.B(n_1199),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1199),
.A2(n_1197),
.B(n_1204),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1190),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1172),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1185),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1210),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1210),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1229),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1163),
.A2(n_1175),
.B1(n_1128),
.B2(n_1225),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1212),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1212),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1188),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1150),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1160),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1158),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1193),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1211),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1175),
.B(n_1196),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1233),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1138),
.A2(n_1149),
.B(n_1128),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1123),
.A2(n_1225),
.B1(n_1213),
.B2(n_1240),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1188),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1138),
.A2(n_1179),
.B1(n_1181),
.B2(n_1158),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1235),
.A2(n_1158),
.B1(n_1150),
.B2(n_1152),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1152),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1152),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1167),
.Y(n_1349)
);

CKINVDCx14_ASAP7_75t_R g1350 ( 
.A(n_1113),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1139),
.A2(n_1234),
.B(n_1208),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1121),
.A2(n_902),
.B1(n_1060),
.B2(n_1054),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1173),
.B(n_1177),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1116),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1154),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1139),
.A2(n_1234),
.B(n_1208),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1215),
.A2(n_874),
.B1(n_902),
.B2(n_1054),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1215),
.A2(n_874),
.B1(n_902),
.B2(n_1054),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1256),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1320),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1312),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1331),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1285),
.A2(n_1251),
.B(n_1259),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1245),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1268),
.Y(n_1366)
);

INVx4_ASAP7_75t_SL g1367 ( 
.A(n_1272),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1268),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1245),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1299),
.B(n_1273),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1324),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1316),
.B(n_1353),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1322),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1316),
.B(n_1353),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1322),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1291),
.B(n_1323),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1263),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1243),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1291),
.B(n_1323),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1249),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1281),
.A2(n_1249),
.B(n_1255),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1352),
.A2(n_1358),
.B1(n_1357),
.B2(n_1282),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1261),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1263),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1299),
.B(n_1274),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1243),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1261),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1267),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1244),
.A2(n_1262),
.B1(n_1264),
.B2(n_1287),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1331),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1324),
.B(n_1291),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1331),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1287),
.B(n_1309),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1310),
.B(n_1309),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1313),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1267),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1252),
.B(n_1302),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1310),
.B(n_1313),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1351),
.A2(n_1356),
.B(n_1303),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1266),
.B(n_1300),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1332),
.B(n_1338),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1344),
.B(n_1292),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1261),
.B(n_1275),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1278),
.B(n_1260),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1269),
.B(n_1250),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1350),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1314),
.A2(n_1265),
.B(n_1337),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1269),
.B(n_1280),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1284),
.B(n_1257),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1314),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1289),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1355),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1296),
.A2(n_1301),
.B1(n_1330),
.B2(n_1308),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1317),
.A2(n_1242),
.B(n_1349),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1290),
.B(n_1298),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1354),
.B(n_1246),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1247),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1304),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1275),
.B(n_1308),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1326),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1275),
.B(n_1349),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1339),
.B(n_1276),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1339),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1271),
.B(n_1341),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1408),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1372),
.B(n_1340),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1372),
.B(n_1325),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1408),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1408),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1374),
.B(n_1276),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1374),
.B(n_1318),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1374),
.B(n_1347),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1365),
.B(n_1307),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1392),
.B(n_1307),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1382),
.A2(n_1345),
.B1(n_1329),
.B2(n_1342),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1390),
.A2(n_1329),
.B1(n_1297),
.B2(n_1315),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1359),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1371),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1370),
.B(n_1253),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1413),
.B(n_1412),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1413),
.B(n_1321),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1415),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1388),
.A2(n_1297),
.B1(n_1279),
.B2(n_1293),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1360),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1423),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1388),
.A2(n_1270),
.B(n_1319),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1415),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1360),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1396),
.Y(n_1451)
);

INVxp67_ASAP7_75t_SL g1452 ( 
.A(n_1412),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1396),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1321),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1387),
.B(n_1402),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1387),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1364),
.Y(n_1457)
);

NAND2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1407),
.B(n_1333),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1364),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1373),
.B(n_1348),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1425),
.B(n_1335),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1423),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1377),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1375),
.B(n_1336),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1377),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1425),
.B(n_1336),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1398),
.A2(n_1253),
.B1(n_1305),
.B2(n_1333),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1414),
.A2(n_1254),
.B1(n_1350),
.B2(n_1343),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1410),
.B(n_1321),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1401),
.A2(n_1254),
.B1(n_1343),
.B2(n_1306),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1467),
.B(n_1420),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1468),
.A2(n_1398),
.B(n_1379),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1468),
.A2(n_1379),
.B(n_1376),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_SL g1474 ( 
.A(n_1470),
.B(n_1376),
.C(n_1379),
.D(n_1384),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1448),
.A2(n_1385),
.B1(n_1403),
.B2(n_1378),
.C(n_1386),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1470),
.A2(n_1394),
.B1(n_1387),
.B2(n_1383),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1426),
.A2(n_1363),
.B(n_1400),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1457),
.B(n_1384),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1459),
.B(n_1397),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1463),
.B(n_1397),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1465),
.B(n_1409),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1448),
.B(n_1424),
.C(n_1419),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1438),
.B(n_1424),
.C(n_1437),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1441),
.B(n_1420),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1443),
.A2(n_1376),
.B1(n_1394),
.B2(n_1375),
.C(n_1416),
.Y(n_1485)
);

NAND4xp25_ASAP7_75t_L g1486 ( 
.A(n_1442),
.B(n_1416),
.C(n_1406),
.D(n_1417),
.Y(n_1486)
);

OAI221xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1436),
.A2(n_1402),
.B1(n_1399),
.B2(n_1417),
.C(n_1391),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1438),
.B(n_1419),
.C(n_1393),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1447),
.B(n_1402),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1452),
.B(n_1409),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1434),
.B(n_1406),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1460),
.B(n_1393),
.C(n_1391),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1434),
.B(n_1406),
.Y(n_1493)
);

OA211x2_ASAP7_75t_L g1494 ( 
.A1(n_1454),
.A2(n_1405),
.B(n_1367),
.C(n_1346),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1455),
.A2(n_1387),
.B(n_1383),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1402),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1399),
.C(n_1420),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1445),
.B(n_1420),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1462),
.B(n_1362),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1445),
.A2(n_1422),
.B1(n_1404),
.B2(n_1395),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1429),
.B(n_1369),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1418),
.C(n_1421),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1429),
.B(n_1369),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1433),
.B(n_1432),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1439),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1433),
.B(n_1369),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1469),
.B(n_1254),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1458),
.B(n_1286),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1435),
.B(n_1286),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1466),
.B(n_1361),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1436),
.A2(n_1368),
.B1(n_1366),
.B2(n_1405),
.C(n_1418),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1427),
.B(n_1389),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1461),
.B(n_1404),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1464),
.B(n_1411),
.C(n_1425),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1427),
.B(n_1389),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1510),
.B(n_1444),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1505),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1505),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1510),
.B(n_1428),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1502),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1514),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1477),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1502),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1492),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1499),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1481),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1478),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1495),
.B(n_1455),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1479),
.Y(n_1531)
);

NAND2x1_ASAP7_75t_L g1532 ( 
.A(n_1495),
.B(n_1426),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1480),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1482),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1483),
.A2(n_1380),
.B1(n_1381),
.B2(n_1395),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1491),
.B(n_1440),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1493),
.B(n_1451),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1497),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1486),
.B(n_1430),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1512),
.B(n_1430),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1431),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1521),
.B(n_1444),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1518),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_SL g1546 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_1444),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1521),
.B(n_1444),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1541),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1517),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1517),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1520),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1520),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1473),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1538),
.B(n_1513),
.Y(n_1557)
);

AND2x2_ASAP7_75t_SL g1558 ( 
.A(n_1535),
.B(n_1540),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1541),
.B(n_1485),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1522),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1532),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1542),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1542),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1449),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1568)
);

NAND2x1_ASAP7_75t_L g1569 ( 
.A(n_1530),
.B(n_1455),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1534),
.B(n_1472),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1529),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1506),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1534),
.A2(n_1474),
.B(n_1488),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1522),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1543),
.Y(n_1576)
);

NOR2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1524),
.B(n_1248),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1522),
.Y(n_1578)
);

NAND2x1_ASAP7_75t_SL g1579 ( 
.A(n_1562),
.B(n_1526),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1543),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1516),
.Y(n_1581)
);

OAI221xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1570),
.A2(n_1535),
.B1(n_1475),
.B2(n_1500),
.C(n_1530),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1545),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1557),
.B(n_1516),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1550),
.B(n_1543),
.Y(n_1586)
);

OAI322xp33_ASAP7_75t_L g1587 ( 
.A1(n_1546),
.A2(n_1528),
.A3(n_1531),
.B1(n_1533),
.B2(n_1527),
.C1(n_1532),
.C2(n_1537),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1547),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1547),
.Y(n_1589)
);

OAI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1570),
.A2(n_1476),
.A3(n_1498),
.B(n_1471),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1563),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1558),
.B(n_1528),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1562),
.Y(n_1594)
);

AND3x1_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1508),
.C(n_1509),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.B(n_1526),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1558),
.A2(n_1573),
.B1(n_1577),
.B2(n_1556),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1553),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1553),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1563),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1556),
.B(n_1539),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1554),
.B(n_1539),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1577),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1572),
.B(n_1507),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1551),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1562),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1555),
.B(n_1527),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1572),
.B(n_1538),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1555),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1532),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1559),
.B(n_1525),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1561),
.B(n_1525),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1564),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1564),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1566),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1538),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_L g1620 ( 
.A(n_1544),
.B(n_1530),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1569),
.B(n_1456),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1597),
.B(n_1561),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1620),
.B(n_1544),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1592),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1544),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1583),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1591),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1596),
.B(n_1566),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1575),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1575),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1619),
.B(n_1548),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1619),
.B(n_1548),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1602),
.B(n_1576),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1608),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1580),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1601),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1595),
.A2(n_1530),
.B1(n_1500),
.B2(n_1569),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1612),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1579),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1616),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1607),
.B(n_1576),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1580),
.Y(n_1652)
);

AOI222xp33_ASAP7_75t_L g1653 ( 
.A1(n_1593),
.A2(n_1549),
.B1(n_1571),
.B2(n_1537),
.C1(n_1568),
.C2(n_1536),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1604),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1594),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1598),
.Y(n_1657)
);

INVx3_ASAP7_75t_SL g1658 ( 
.A(n_1630),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1625),
.A2(n_1606),
.B1(n_1611),
.B2(n_1530),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1585),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1625),
.A2(n_1582),
.B(n_1611),
.Y(n_1661)
);

INVxp33_ASAP7_75t_L g1662 ( 
.A(n_1622),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1657),
.B(n_1590),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1615),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1655),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1626),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1648),
.A2(n_1605),
.B(n_1610),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1645),
.A2(n_1530),
.B1(n_1618),
.B2(n_1617),
.Y(n_1668)
);

AOI31xp33_ASAP7_75t_L g1669 ( 
.A1(n_1651),
.A2(n_1248),
.A3(n_1277),
.B(n_1621),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1653),
.A2(n_1586),
.B(n_1609),
.C(n_1594),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1643),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1626),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1586),
.Y(n_1673)
);

AOI222xp33_ASAP7_75t_L g1674 ( 
.A1(n_1633),
.A2(n_1549),
.B1(n_1585),
.B2(n_1609),
.C1(n_1484),
.C2(n_1551),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1628),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1529),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1621),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1652),
.B(n_1529),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1648),
.A2(n_1494),
.B1(n_1530),
.B2(n_1380),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1628),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1629),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1652),
.B(n_1529),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1658),
.B(n_1636),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1671),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1671),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1678),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1662),
.B(n_1637),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1677),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1663),
.B(n_1637),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1631),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1666),
.B(n_1629),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1670),
.A2(n_1638),
.B1(n_1623),
.B2(n_1641),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1641),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1678),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1672),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1659),
.A2(n_1638),
.B1(n_1623),
.B2(n_1650),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1675),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1681),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1665),
.B(n_1664),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1660),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1697),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1691),
.A2(n_1667),
.B(n_1668),
.Y(n_1705)
);

OAI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1699),
.A2(n_1674),
.B(n_1680),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1682),
.Y(n_1707)
);

NAND4xp75_ASAP7_75t_L g1708 ( 
.A(n_1691),
.B(n_1656),
.C(n_1679),
.D(n_1676),
.Y(n_1708)
);

AOI322xp5_ASAP7_75t_L g1709 ( 
.A1(n_1702),
.A2(n_1680),
.A3(n_1640),
.B1(n_1650),
.B2(n_1649),
.C1(n_1639),
.C2(n_1647),
.Y(n_1709)
);

AOI31xp33_ASAP7_75t_L g1710 ( 
.A1(n_1686),
.A2(n_1277),
.A3(n_1635),
.B(n_1656),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1684),
.A2(n_1702),
.B(n_1693),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1695),
.A2(n_1683),
.B1(n_1649),
.B2(n_1647),
.C(n_1646),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1693),
.B(n_1635),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1704),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1706),
.A2(n_1689),
.B1(n_1703),
.B2(n_1696),
.C(n_1692),
.Y(n_1716)
);

NAND4xp75_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1694),
.C(n_1712),
.D(n_1687),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1711),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1707),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1714),
.A2(n_1690),
.B1(n_1708),
.B2(n_1688),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1710),
.B(n_1698),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1709),
.B(n_1700),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1639),
.C(n_1632),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1716),
.A2(n_1646),
.B(n_1644),
.C(n_1632),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_SL g1726 ( 
.A(n_1720),
.B(n_1644),
.C(n_1627),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1722),
.B(n_1642),
.C(n_1627),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1723),
.B(n_1642),
.C(n_1627),
.Y(n_1728)
);

NOR2x2_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1624),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_L g1730 ( 
.A(n_1721),
.B(n_1634),
.C(n_1624),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1728),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1727),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1718),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1719),
.B1(n_1624),
.B2(n_1642),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1729),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1729),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_SL g1738 ( 
.A(n_1734),
.B(n_1724),
.C(n_1487),
.Y(n_1738)
);

NAND4xp75_ASAP7_75t_L g1739 ( 
.A(n_1736),
.B(n_1634),
.C(n_1640),
.D(n_1494),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1737),
.B(n_1634),
.Y(n_1740)
);

NOR2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1733),
.B(n_1334),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1732),
.B(n_1567),
.Y(n_1742)
);

XNOR2x1_ASAP7_75t_L g1743 ( 
.A(n_1741),
.B(n_1731),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1740),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1742),
.Y(n_1745)
);

AOI22x1_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1731),
.B1(n_1735),
.B2(n_1738),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1746),
.B(n_1745),
.C(n_1744),
.D(n_1743),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_SL g1748 ( 
.A1(n_1747),
.A2(n_1739),
.B(n_1565),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1747),
.A2(n_1578),
.B1(n_1560),
.B2(n_1565),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1748),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1749),
.A2(n_1565),
.B(n_1560),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1750),
.A2(n_1574),
.B(n_1560),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1751),
.B(n_1578),
.C(n_1574),
.Y(n_1753)
);

XNOR2xp5_ASAP7_75t_L g1754 ( 
.A(n_1752),
.B(n_1404),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_R g1755 ( 
.A1(n_1754),
.A2(n_1753),
.B1(n_1453),
.B2(n_1446),
.C(n_1450),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_R g1756 ( 
.A1(n_1755),
.A2(n_1294),
.B1(n_1578),
.B2(n_1574),
.C(n_1552),
.Y(n_1756)
);

AOI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1272),
.B(n_1311),
.C(n_1295),
.Y(n_1757)
);


endmodule