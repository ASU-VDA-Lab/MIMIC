module fake_jpeg_29335_n_398 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_398);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_398;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_44),
.B(n_48),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_77),
.Y(n_103)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_51),
.B(n_58),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_19),
.B(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_13),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_15),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_15),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_21),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_29),
.CON(n_87),
.SN(n_87)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_27),
.B1(n_39),
.B2(n_33),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_85),
.A2(n_93),
.B1(n_96),
.B2(n_112),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_27),
.B1(n_39),
.B2(n_33),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_59),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_117),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_22),
.B1(n_42),
.B2(n_40),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_39),
.B1(n_43),
.B2(n_31),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_29),
.B(n_31),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_108),
.A2(n_52),
.B(n_66),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_50),
.A2(n_17),
.B1(n_40),
.B2(n_37),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_119),
.B1(n_122),
.B2(n_69),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_47),
.A2(n_42),
.B1(n_22),
.B2(n_35),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_54),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_55),
.A2(n_41),
.B1(n_36),
.B2(n_20),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_127),
.B1(n_4),
.B2(n_5),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_61),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_62),
.B1(n_77),
.B2(n_79),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_137),
.B(n_147),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_91),
.CI(n_96),
.CON(n_140),
.SN(n_140)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_140),
.B(n_176),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_87),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_142),
.B(n_159),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_58),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_63),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_68),
.B1(n_67),
.B2(n_70),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_166),
.B1(n_100),
.B2(n_124),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx10_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_69),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_64),
.C(n_46),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_129),
.C(n_92),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_98),
.B(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_121),
.B(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_106),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_80),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_164),
.B(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_85),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_172),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_104),
.A2(n_80),
.B1(n_52),
.B2(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_108),
.B(n_1),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_131),
.B(n_1),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_3),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_3),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_179),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_105),
.Y(n_174)
);

INVx2_ASAP7_75t_R g218 ( 
.A(n_174),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_177),
.B1(n_123),
.B2(n_95),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_100),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_88),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_88),
.B(n_7),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_8),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_8),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_104),
.B(n_9),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_156),
.B(n_176),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_182),
.A2(n_187),
.B1(n_192),
.B2(n_208),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_200),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_97),
.B1(n_130),
.B2(n_129),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_95),
.B1(n_123),
.B2(n_97),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_203),
.C(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_92),
.C(n_9),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_219),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_147),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_10),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_171),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_11),
.B1(n_12),
.B2(n_138),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_137),
.B1(n_163),
.B2(n_172),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_140),
.B(n_158),
.C(n_144),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_140),
.B(n_167),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_136),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_221),
.B(n_223),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_222),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_253),
.B1(n_214),
.B2(n_204),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_159),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_146),
.B1(n_138),
.B2(n_176),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_231),
.A2(n_251),
.B1(n_255),
.B2(n_199),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_173),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_181),
.B1(n_216),
.B2(n_190),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_234),
.A2(n_231),
.B1(n_255),
.B2(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_143),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_236),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_138),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_184),
.B(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_237),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_250),
.B(n_252),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_134),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_183),
.B(n_150),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_244),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_160),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_249),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_168),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_247),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_170),
.B(n_162),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_203),
.B(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_184),
.B(n_157),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_216),
.A2(n_169),
.B(n_145),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_145),
.B1(n_174),
.B2(n_154),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_202),
.A2(n_151),
.B(n_153),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_212),
.A2(n_174),
.B1(n_155),
.B2(n_135),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_153),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_236),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_182),
.A2(n_153),
.B1(n_208),
.B2(n_190),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_222),
.B1(n_240),
.B2(n_226),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_260),
.B(n_273),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_193),
.B(n_205),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_263),
.B(n_268),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_211),
.B1(n_209),
.B2(n_189),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_209),
.B(n_189),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_245),
.C(n_254),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_234),
.A2(n_201),
.B(n_199),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_197),
.B(n_201),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_234),
.A2(n_197),
.B(n_220),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_196),
.B(n_220),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_224),
.A2(n_191),
.B1(n_215),
.B2(n_196),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_277),
.B1(n_223),
.B2(n_239),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_237),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_283),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_234),
.A2(n_252),
.B(n_232),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_286),
.B(n_249),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_232),
.A2(n_253),
.B(n_248),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_288),
.A2(n_261),
.B1(n_277),
.B2(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_262),
.B(n_235),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_259),
.B(n_264),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_297),
.C(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_289),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_269),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_226),
.C(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_303),
.B1(n_306),
.B2(n_256),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_229),
.B1(n_242),
.B2(n_224),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_233),
.B1(n_230),
.B2(n_228),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_307),
.Y(n_317)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_225),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_221),
.C(n_227),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_241),
.Y(n_311)
);

OA21x2_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_259),
.B(n_264),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_312),
.B(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_314),
.B(n_316),
.Y(n_345)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_315),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_295),
.B(n_285),
.C(n_266),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_304),
.B(n_301),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_302),
.B(n_280),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_311),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_280),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_325),
.B(n_326),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_287),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_330),
.B1(n_303),
.B2(n_260),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_286),
.B1(n_273),
.B2(n_266),
.Y(n_330)
);

OAI322xp33_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_306),
.A3(n_275),
.B1(n_283),
.B2(n_292),
.C1(n_310),
.C2(n_297),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_335),
.B(n_349),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_324),
.Y(n_359)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_301),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_338),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_289),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_258),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_318),
.B(n_304),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_257),
.C(n_271),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.C(n_350),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_263),
.C(n_307),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_347),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_323),
.A2(n_300),
.B1(n_317),
.B2(n_330),
.Y(n_348)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_313),
.B(n_308),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_261),
.C(n_270),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_317),
.B1(n_323),
.B2(n_261),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_343),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_353),
.B(n_359),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_361),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_282),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_355),
.A2(n_334),
.B1(n_342),
.B2(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_340),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_366),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_345),
.B(n_334),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_368),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_346),
.C(n_345),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_344),
.C(n_336),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_371),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_363),
.B(n_320),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_320),
.Y(n_373)
);

AOI221xp5_ASAP7_75t_L g375 ( 
.A1(n_373),
.A2(n_351),
.B1(n_352),
.B2(n_357),
.C(n_329),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_350),
.C(n_341),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_372),
.C(n_369),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_375),
.B(n_378),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_366),
.A2(n_353),
.B(n_352),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_365),
.A2(n_355),
.B1(n_332),
.B2(n_331),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_374),
.A2(n_328),
.B1(n_290),
.B2(n_293),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_379),
.B(n_360),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_387),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_372),
.C(n_369),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_377),
.B(n_294),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_382),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_385),
.A2(n_376),
.A3(n_380),
.B1(n_382),
.B2(n_381),
.C1(n_298),
.C2(n_282),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_L g395 ( 
.A1(n_390),
.A2(n_393),
.A3(n_384),
.B1(n_284),
.B2(n_278),
.C1(n_282),
.C2(n_241),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_284),
.B(n_393),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_SL g397 ( 
.A(n_396),
.B(n_394),
.C(n_391),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_359),
.Y(n_398)
);


endmodule