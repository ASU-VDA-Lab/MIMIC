module fake_jpeg_25237_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_2),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

NAND2x1_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_18),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_20),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_17),
.B1(n_27),
.B2(n_22),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_26),
.B1(n_19),
.B2(n_21),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_20),
.C(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_31),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_42),
.B1(n_27),
.B2(n_22),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_79),
.B1(n_46),
.B2(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_22),
.B1(n_27),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_78),
.B1(n_81),
.B2(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_23),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_85),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_38),
.B1(n_30),
.B2(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_47),
.C(n_52),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_62),
.C(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_100),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_18),
.B(n_44),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_98),
.B(n_66),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_97),
.B1(n_109),
.B2(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_49),
.B1(n_46),
.B2(n_51),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_48),
.B(n_2),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_80),
.B1(n_61),
.B2(n_10),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_1),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_4),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_5),
.B(n_6),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_48),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_77),
.B1(n_74),
.B2(n_62),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_130),
.B1(n_96),
.B2(n_105),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_120),
.B(n_96),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_89),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_122),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_102),
.B1(n_99),
.B2(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_113),
.C(n_122),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_87),
.B(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_125),
.C(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_101),
.B1(n_91),
.B2(n_87),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_142),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_91),
.B1(n_87),
.B2(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_127),
.B1(n_123),
.B2(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_148),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_143),
.B1(n_139),
.B2(n_133),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_131),
.B(n_134),
.Y(n_174)
);

BUFx12f_ASAP7_75t_SL g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_164),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_163),
.C(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_165),
.B1(n_147),
.B2(n_134),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_125),
.C(n_90),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_90),
.B1(n_8),
.B2(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_177),
.C(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_161),
.B1(n_141),
.B2(n_146),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_165),
.B(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_136),
.C(n_133),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_177),
.C(n_167),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_180),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_175),
.B(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_158),
.B1(n_164),
.B2(n_153),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_158),
.B1(n_136),
.B2(n_135),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.C(n_61),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_191),
.B(n_7),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_146),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_151),
.B1(n_186),
.B2(n_183),
.C(n_176),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_141),
.B(n_159),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_184),
.A3(n_179),
.B1(n_185),
.B2(n_189),
.C1(n_178),
.C2(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_196),
.C(n_8),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_13),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_8),
.B(n_11),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_11),
.C(n_12),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_195),
.A2(n_14),
.B(n_15),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_202),
.B1(n_194),
.B2(n_12),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);


endmodule