module fake_jpeg_12865_n_405 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_405);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_62),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_9),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_36),
.B(n_0),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_9),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_34),
.B1(n_39),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_27),
.B1(n_68),
.B2(n_67),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_34),
.B1(n_39),
.B2(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_27),
.B1(n_39),
.B2(n_33),
.Y(n_121)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_39),
.B1(n_33),
.B2(n_27),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_69),
.C(n_71),
.Y(n_119)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_31),
.B1(n_26),
.B2(n_32),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_113),
.B1(n_44),
.B2(n_51),
.Y(n_115)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_32),
.B1(n_26),
.B2(n_17),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_116),
.B(n_126),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_54),
.B1(n_63),
.B2(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_117),
.A2(n_137),
.B1(n_87),
.B2(n_110),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_70),
.B(n_29),
.C(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_132),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_119),
.B(n_43),
.Y(n_179)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_124),
.B1(n_147),
.B2(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_40),
.C(n_18),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_131),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_129),
.B(n_134),
.Y(n_166)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_58),
.CON(n_129),
.SN(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_48),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_138),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_82),
.B(n_59),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_50),
.B1(n_46),
.B2(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_57),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_29),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_29),
.A3(n_43),
.B1(n_18),
.B2(n_52),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_47),
.CI(n_94),
.CON(n_165),
.SN(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_148),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_41),
.B1(n_26),
.B2(n_32),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_55),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_37),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_37),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_163),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_86),
.B(n_92),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_99),
.B1(n_83),
.B2(n_127),
.Y(n_202)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_183),
.Y(n_214)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_121),
.B1(n_76),
.B2(n_80),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_134),
.Y(n_203)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_140),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_133),
.A2(n_105),
.B(n_79),
.Y(n_183)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_132),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_138),
.C(n_135),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_212),
.C(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_143),
.B1(n_139),
.B2(n_124),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_202),
.B1(n_210),
.B2(n_155),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_116),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_190),
.B(n_199),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_195),
.B1(n_196),
.B2(n_182),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_118),
.B1(n_122),
.B2(n_114),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_114),
.B1(n_120),
.B2(n_123),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_144),
.B1(n_136),
.B2(n_142),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_176),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_128),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_161),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_110),
.B1(n_106),
.B2(n_80),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_128),
.C(n_105),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_23),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_222),
.B1(n_229),
.B2(n_192),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_242),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_165),
.B1(n_168),
.B2(n_170),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_225),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_200),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_179),
.B1(n_173),
.B2(n_154),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_184),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_173),
.C(n_154),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_240),
.B1(n_191),
.B2(n_184),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_152),
.B1(n_160),
.B2(n_176),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_246),
.B1(n_235),
.B2(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_155),
.B1(n_152),
.B2(n_160),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_241),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g243 ( 
.A1(n_186),
.A2(n_213),
.A3(n_198),
.B1(n_195),
.B2(n_203),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_215),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_185),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_174),
.B(n_158),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_198),
.A2(n_106),
.B1(n_87),
.B2(n_180),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_251),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_270),
.C(n_250),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_206),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_252),
.A2(n_263),
.B(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_275),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_259),
.B1(n_274),
.B2(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_226),
.B(n_201),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_164),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_269),
.B(n_157),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_164),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_215),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_187),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_242),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_285),
.C(n_290),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_218),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_283),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_220),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_222),
.B1(n_229),
.B2(n_225),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_301),
.B1(n_274),
.B2(n_267),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_220),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_241),
.B(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_288),
.B(n_302),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.Y(n_290)
);

XNOR2x2_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_239),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_295),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_253),
.B(n_241),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_217),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_297),
.C(n_299),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_246),
.C(n_216),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_187),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_201),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_140),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_35),
.B1(n_23),
.B2(n_146),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_248),
.C(n_276),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_306),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_260),
.B(n_266),
.Y(n_305)
);

AO22x1_ASAP7_75t_L g334 ( 
.A1(n_305),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_247),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_251),
.B1(n_257),
.B2(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_313),
.A2(n_35),
.B1(n_111),
.B2(n_81),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_289),
.A2(n_255),
.B1(n_35),
.B2(n_94),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_320),
.Y(n_328)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_255),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_322),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_111),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_12),
.Y(n_326)
);

AO221x1_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_291),
.B1(n_16),
.B2(n_15),
.C(n_10),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_282),
.C(n_278),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_333),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_283),
.C(n_285),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_12),
.B(n_16),
.C(n_15),
.Y(n_358)
);

BUFx12_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_293),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_339),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_340),
.A2(n_311),
.B1(n_305),
.B2(n_307),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_11),
.B(n_16),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_342),
.A2(n_310),
.B(n_320),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_321),
.B(n_322),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_354),
.B(n_358),
.Y(n_371)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_346),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_343),
.Y(n_349)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_304),
.B1(n_324),
.B2(n_309),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_359),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_309),
.C(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_356),
.C(n_357),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_316),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_325),
.C(n_316),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_37),
.C(n_21),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_336),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_37),
.C(n_21),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_357),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_355),
.A2(n_335),
.B(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_361),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_352),
.A2(n_335),
.B(n_342),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_358),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_344),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_356),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_353),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_355),
.A2(n_332),
.B(n_340),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_373),
.B1(n_358),
.B2(n_360),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_13),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_0),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_374),
.B(n_384),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_376),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_380),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_379),
.A2(n_371),
.B(n_369),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_22),
.C(n_21),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_22),
.C(n_21),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_1),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_361),
.A2(n_2),
.B(n_3),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_383),
.A2(n_362),
.B(n_373),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_368),
.B(n_363),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_391),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_388),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_366),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_375),
.B(n_6),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_3),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_379),
.C(n_381),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_398),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_387),
.B(n_380),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_396),
.A2(n_397),
.B(n_393),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_2),
.B(n_3),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_390),
.C(n_5),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_401),
.C(n_400),
.Y(n_402)
);

AOI311xp33_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_4),
.A3(n_5),
.B(n_6),
.C(n_378),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_4),
.C(n_6),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_4),
.Y(n_405)
);


endmodule