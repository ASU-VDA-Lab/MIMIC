module fake_netlist_6_3356_n_15804 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_15804);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_15804;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_2542;
wire n_1671;
wire n_14428;
wire n_2817;
wire n_13611;
wire n_15214;
wire n_801;
wire n_4452;
wire n_6566;
wire n_2576;
wire n_5172;
wire n_13045;
wire n_11173;
wire n_15268;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_10487;
wire n_6872;
wire n_13998;
wire n_1351;
wire n_5254;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_14769;
wire n_2157;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_10587;
wire n_5019;
wire n_2332;
wire n_8713;
wire n_15450;
wire n_10960;
wire n_6141;
wire n_7111;
wire n_3849;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_578;
wire n_5138;
wire n_13522;
wire n_10931;
wire n_4395;
wire n_4388;
wire n_6960;
wire n_1061;
wire n_15609;
wire n_3089;
wire n_12265;
wire n_8169;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_783;
wire n_7180;
wire n_11574;
wire n_5653;
wire n_4978;
wire n_13530;
wire n_8604;
wire n_15049;
wire n_5409;
wire n_5301;
wire n_13125;
wire n_7263;
wire n_188;
wire n_1854;
wire n_15181;
wire n_3088;
wire n_8168;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_8186;
wire n_7504;
wire n_677;
wire n_6126;
wire n_6725;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_12322;
wire n_14318;
wire n_8899;
wire n_14196;
wire n_2317;
wire n_5524;
wire n_10236;
wire n_442;
wire n_5345;
wire n_11205;
wire n_11678;
wire n_11776;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_1975;
wire n_11650;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_2179;
wire n_8534;
wire n_5963;
wire n_12179;
wire n_13942;
wire n_5055;
wire n_15294;
wire n_14439;
wire n_1547;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_11905;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_893;
wire n_14825;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_4249;
wire n_11536;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_9104;
wire n_1844;
wire n_14914;
wire n_6999;
wire n_14741;
wire n_15295;
wire n_15665;
wire n_11046;
wire n_11079;
wire n_1555;
wire n_5548;
wire n_10283;
wire n_5057;
wire n_15581;
wire n_11065;
wire n_15445;
wire n_8339;
wire n_8272;
wire n_14215;
wire n_13997;
wire n_14402;
wire n_7161;
wire n_3030;
wire n_830;
wire n_7868;
wire n_14882;
wire n_5838;
wire n_15764;
wire n_5725;
wire n_6324;
wire n_13437;
wire n_447;
wire n_15623;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_3427;
wire n_852;
wire n_11214;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_7000;
wire n_8561;
wire n_14944;
wire n_14998;
wire n_11954;
wire n_7398;
wire n_2926;
wire n_1078;
wire n_544;
wire n_14232;
wire n_10392;
wire n_14341;
wire n_12882;
wire n_5900;
wire n_4273;
wire n_15074;
wire n_5545;
wire n_12617;
wire n_8411;
wire n_2321;
wire n_8499;
wire n_2019;
wire n_8236;
wire n_5102;
wire n_15253;
wire n_15356;
wire n_13137;
wire n_3345;
wire n_13221;
wire n_2074;
wire n_6882;
wire n_2919;
wire n_4501;
wire n_9626;
wire n_10775;
wire n_11163;
wire n_2129;
wire n_9526;
wire n_13657;
wire n_15571;
wire n_9840;
wire n_4724;
wire n_6325;
wire n_945;
wire n_14099;
wire n_5598;
wire n_15632;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_10719;
wire n_4997;
wire n_2399;
wire n_7389;
wire n_9018;
wire n_4843;
wire n_11419;
wire n_1232;
wire n_8070;
wire n_12095;
wire n_13663;
wire n_13990;
wire n_4696;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_14939;
wire n_11740;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_13993;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_3877;
wire n_12392;
wire n_15353;
wire n_3929;
wire n_8366;
wire n_3048;
wire n_1455;
wire n_9362;
wire n_11979;
wire n_8102;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_567;
wire n_1781;
wire n_1971;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_15797;
wire n_9962;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_10373;
wire n_3077;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_8913;
wire n_9525;
wire n_3107;
wire n_10816;
wire n_9725;
wire n_155;
wire n_4956;
wire n_11537;
wire n_14699;
wire n_13814;
wire n_12707;
wire n_454;
wire n_14861;
wire n_7686;
wire n_1421;
wire n_3664;
wire n_6914;
wire n_1936;
wire n_5337;
wire n_10335;
wire n_15194;
wire n_15362;
wire n_5129;
wire n_11301;
wire n_12424;
wire n_13681;
wire n_14121;
wire n_15101;
wire n_5420;
wire n_15572;
wire n_1660;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_713;
wire n_11703;
wire n_11699;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_6374;
wire n_2843;
wire n_7651;
wire n_11543;
wire n_10947;
wire n_6628;
wire n_13483;
wire n_8125;
wire n_3760;
wire n_6015;
wire n_14662;
wire n_11261;
wire n_14811;
wire n_10226;
wire n_13247;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_6526;
wire n_13929;
wire n_1894;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_3347;
wire n_10767;
wire n_15421;
wire n_5136;
wire n_907;
wire n_8040;
wire n_8535;
wire n_14646;
wire n_11821;
wire n_14095;
wire n_5638;
wire n_13121;
wire n_13989;
wire n_9100;
wire n_14864;
wire n_15069;
wire n_4110;
wire n_6784;
wire n_1658;
wire n_12107;
wire n_14520;
wire n_10755;
wire n_4950;
wire n_14780;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_6323;
wire n_9614;
wire n_14431;
wire n_15200;
wire n_13515;
wire n_10682;
wire n_6110;
wire n_1967;
wire n_11684;
wire n_3999;
wire n_12652;
wire n_3928;
wire n_6371;
wire n_14410;
wire n_8079;
wire n_10699;
wire n_2613;
wire n_15507;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_2708;
wire n_15800;
wire n_1648;
wire n_9400;
wire n_5151;
wire n_1911;
wire n_8142;
wire n_11627;
wire n_2011;
wire n_5684;
wire n_13139;
wire n_8598;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_13803;
wire n_281;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_14066;
wire n_7856;
wire n_7774;
wire n_15600;
wire n_564;
wire n_5680;
wire n_6674;
wire n_13606;
wire n_6148;
wire n_6951;
wire n_11659;
wire n_13501;
wire n_279;
wire n_686;
wire n_7625;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_9106;
wire n_13509;
wire n_12775;
wire n_2735;
wire n_13729;
wire n_4662;
wire n_8869;
wire n_7863;
wire n_4671;
wire n_6989;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14813;
wire n_4314;
wire n_9520;
wire n_2080;
wire n_14791;
wire n_8958;
wire n_14485;
wire n_14931;
wire n_12833;
wire n_323;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_14628;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_13687;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_1381;
wire n_331;
wire n_1699;
wire n_2093;
wire n_12371;
wire n_4296;
wire n_10114;
wire n_12203;
wire n_10357;
wire n_14540;
wire n_15762;
wire n_7147;
wire n_2770;
wire n_8115;
wire n_608;
wire n_2101;
wire n_4507;
wire n_9398;
wire n_8389;
wire n_5902;
wire n_11497;
wire n_512;
wire n_14900;
wire n_15320;
wire n_3484;
wire n_12359;
wire n_4677;
wire n_792;
wire n_12915;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_1328;
wire n_2917;
wire n_13149;
wire n_13711;
wire n_13454;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_12742;
wire n_3923;
wire n_14091;
wire n_9042;
wire n_15755;
wire n_11768;
wire n_3900;
wire n_8412;
wire n_9267;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_14478;
wire n_8987;
wire n_11805;
wire n_14461;
wire n_6485;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_1910;
wire n_13958;
wire n_1075;
wire n_3980;
wire n_14935;
wire n_2998;
wire n_15332;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_237;
wire n_6863;
wire n_6282;
wire n_6994;
wire n_12770;
wire n_1895;
wire n_10012;
wire n_14570;
wire n_4294;
wire n_13754;
wire n_12985;
wire n_4698;
wire n_13797;
wire n_4445;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_7564;
wire n_11635;
wire n_3859;
wire n_14989;
wire n_15434;
wire n_2692;
wire n_175;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_14171;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_10296;
wire n_8119;
wire n_3397;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_15212;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_9718;
wire n_9128;
wire n_2469;
wire n_10281;
wire n_13344;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_14380;
wire n_8748;
wire n_3927;
wire n_13984;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_14239;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_8718;
wire n_7110;
wire n_764;
wire n_5476;
wire n_2764;
wire n_12831;
wire n_13920;
wire n_9935;
wire n_2895;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_14045;
wire n_733;
wire n_14288;
wire n_14824;
wire n_2922;
wire n_10097;
wire n_3882;
wire n_4856;
wire n_8223;
wire n_15767;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_15635;
wire n_4331;
wire n_7297;
wire n_9866;
wire n_10018;
wire n_15183;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_7298;
wire n_15118;
wire n_5536;
wire n_9129;
wire n_10141;
wire n_9858;
wire n_2072;
wire n_12427;
wire n_1354;
wire n_7533;
wire n_14162;
wire n_13771;
wire n_586;
wire n_423;
wire n_7221;
wire n_4375;
wire n_1701;
wire n_13977;
wire n_10656;
wire n_15159;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_2678;
wire n_11295;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_11662;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_1726;
wire n_8246;
wire n_4613;
wire n_8952;
wire n_15679;
wire n_13014;
wire n_2434;
wire n_9070;
wire n_2878;
wire n_11708;
wire n_3875;
wire n_3012;
wire n_10266;
wire n_15629;
wire n_14401;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_10897;
wire n_10827;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_15154;
wire n_14922;
wire n_210;
wire n_10449;
wire n_7569;
wire n_2641;
wire n_7823;
wire n_7861;
wire n_7734;
wire n_8955;
wire n_9680;
wire n_5658;
wire n_4731;
wire n_9477;
wire n_7062;
wire n_12147;
wire n_12172;
wire n_3052;
wire n_12923;
wire n_178;
wire n_7039;
wire n_355;
wire n_8577;
wire n_12384;
wire n_14961;
wire n_11349;
wire n_8594;
wire n_5046;
wire n_13227;
wire n_8428;
wire n_9829;
wire n_15438;
wire n_2749;
wire n_11260;
wire n_3298;
wire n_8848;
wire n_12825;
wire n_2254;
wire n_13341;
wire n_5058;
wire n_10685;
wire n_1926;
wire n_11351;
wire n_3273;
wire n_4467;
wire n_15185;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_14803;
wire n_1747;
wire n_195;
wire n_5667;
wire n_780;
wire n_8259;
wire n_12540;
wire n_15611;
wire n_10607;
wire n_14388;
wire n_2624;
wire n_15490;
wire n_5865;
wire n_15182;
wire n_12249;
wire n_8349;
wire n_6836;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_14977;
wire n_11998;
wire n_4681;
wire n_13239;
wire n_8164;
wire n_4072;
wire n_10628;
wire n_4752;
wire n_4220;
wire n_13429;
wire n_835;
wire n_928;
wire n_5281;
wire n_7905;
wire n_11775;
wire n_8776;
wire n_15100;
wire n_9143;
wire n_10769;
wire n_2092;
wire n_10256;
wire n_8287;
wire n_10368;
wire n_1654;
wire n_6771;
wire n_14732;
wire n_7753;
wire n_7950;
wire n_9947;
wire n_1750;
wire n_1462;
wire n_13999;
wire n_9088;
wire n_8607;
wire n_2514;
wire n_14037;
wire n_10138;
wire n_12117;
wire n_604;
wire n_11706;
wire n_6248;
wire n_11800;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_1588;
wire n_10452;
wire n_11464;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_12960;
wire n_14878;
wire n_14094;
wire n_13033;
wire n_11642;
wire n_15046;
wire n_2468;
wire n_4381;
wire n_11143;
wire n_15703;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_515;
wire n_2096;
wire n_3968;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_12131;
wire n_12851;
wire n_5795;
wire n_11934;
wire n_12349;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_14282;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_514;
wire n_6714;
wire n_15518;
wire n_687;
wire n_11308;
wire n_890;
wire n_13550;
wire n_14217;
wire n_10903;
wire n_7677;
wire n_13348;
wire n_5457;
wire n_8416;
wire n_10396;
wire n_13919;
wire n_2812;
wire n_190;
wire n_4518;
wire n_10724;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_15574;
wire n_11084;
wire n_14062;
wire n_9988;
wire n_1709;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_14167;
wire n_12740;
wire n_2393;
wire n_2657;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_10363;
wire n_2409;
wire n_2252;
wire n_13240;
wire n_3237;
wire n_949;
wire n_8949;
wire n_10831;
wire n_3500;
wire n_3834;
wire n_9131;
wire n_11553;
wire n_10517;
wire n_12578;
wire n_12795;
wire n_4589;
wire n_2075;
wire n_10323;
wire n_12194;
wire n_13623;
wire n_2972;
wire n_10842;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_10876;
wire n_2763;
wire n_11511;
wire n_2762;
wire n_9137;
wire n_15649;
wire n_11180;
wire n_14043;
wire n_9724;
wire n_11146;
wire n_9281;
wire n_3192;
wire n_8995;
wire n_10883;
wire n_760;
wire n_10101;
wire n_1546;
wire n_9393;
wire n_4394;
wire n_6581;
wire n_13845;
wire n_12709;
wire n_2279;
wire n_161;
wire n_6010;
wire n_13432;
wire n_1296;
wire n_3352;
wire n_8711;
wire n_3073;
wire n_7013;
wire n_12771;
wire n_14150;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_7290;
wire n_12278;
wire n_13721;
wire n_595;
wire n_1779;
wire n_524;
wire n_10820;
wire n_13514;
wire n_4921;
wire n_9687;
wire n_1858;
wire n_14787;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_2558;
wire n_7315;
wire n_13194;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_1164;
wire n_4697;
wire n_13244;
wire n_4288;
wire n_4289;
wire n_11866;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_5529;
wire n_3733;
wire n_15659;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_9102;
wire n_1487;
wire n_11526;
wire n_13404;
wire n_9578;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_14785;
wire n_7438;
wire n_14355;
wire n_14128;
wire n_2145;
wire n_7268;
wire n_7337;
wire n_11851;
wire n_898;
wire n_4964;
wire n_9489;
wire n_12804;
wire n_14123;
wire n_5957;
wire n_6965;
wire n_12116;
wire n_10728;
wire n_4228;
wire n_3423;
wire n_10094;
wire n_925;
wire n_1932;
wire n_1101;
wire n_9144;
wire n_13755;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_14105;
wire n_14126;
wire n_7461;
wire n_8285;
wire n_13870;
wire n_4322;
wire n_10655;
wire n_13791;
wire n_3644;
wire n_9797;
wire n_15133;
wire n_6955;
wire n_8483;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_9521;
wire n_15288;
wire n_9932;
wire n_9478;
wire n_1451;
wire n_8332;
wire n_13040;
wire n_320;
wire n_639;
wire n_963;
wire n_2767;
wire n_11370;
wire n_6509;
wire n_7278;
wire n_13900;
wire n_4576;
wire n_7454;
wire n_11253;
wire n_14652;
wire n_11379;
wire n_15527;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_11981;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_9895;
wire n_1521;
wire n_8741;
wire n_12918;
wire n_1366;
wire n_4000;
wire n_11585;
wire n_9351;
wire n_5445;
wire n_2897;
wire n_13140;
wire n_13962;
wire n_14556;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_6839;
wire n_7232;
wire n_13753;
wire n_4345;
wire n_7377;
wire n_5501;
wire n_996;
wire n_532;
wire n_173;
wire n_6646;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_1376;
wire n_12102;
wire n_9189;
wire n_413;
wire n_15149;
wire n_15365;
wire n_4664;
wire n_13716;
wire n_2170;
wire n_4156;
wire n_14844;
wire n_14701;
wire n_948;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_14391;
wire n_7904;
wire n_11691;
wire n_6033;
wire n_977;
wire n_11541;
wire n_15495;
wire n_13610;
wire n_536;
wire n_3158;
wire n_1788;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_13332;
wire n_2643;
wire n_5748;
wire n_14408;
wire n_3782;
wire n_9356;
wire n_15293;
wire n_12865;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_1835;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_5076;
wire n_581;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_432;
wire n_3700;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_10959;
wire n_3104;
wire n_6809;
wire n_11233;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_7840;
wire n_10972;
wire n_4310;
wire n_7782;
wire n_6359;
wire n_1432;
wire n_13213;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_989;
wire n_8800;
wire n_13385;
wire n_15695;
wire n_10845;
wire n_7080;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_2191;
wire n_8229;
wire n_1246;
wire n_4528;
wire n_8410;
wire n_14756;
wire n_14863;
wire n_5811;
wire n_14156;
wire n_899;
wire n_13992;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_1035;
wire n_4914;
wire n_7624;
wire n_4939;
wire n_7629;
wire n_499;
wire n_13790;
wire n_1426;
wire n_3418;
wire n_705;
wire n_14384;
wire n_9735;
wire n_9186;
wire n_10818;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_12552;
wire n_13304;
wire n_2069;
wire n_14633;
wire n_11069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_9941;
wire n_7003;
wire n_11951;
wire n_12222;
wire n_15178;
wire n_11900;
wire n_15699;
wire n_3119;
wire n_14711;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_3735;
wire n_2297;
wire n_11369;
wire n_4379;
wire n_10563;
wire n_14210;
wire n_486;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_1448;
wire n_15788;
wire n_5901;
wire n_13362;
wire n_6538;
wire n_14373;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_8107;
wire n_648;
wire n_11108;
wire n_7010;
wire n_9728;
wire n_12883;
wire n_11004;
wire n_12992;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_6519;
wire n_2103;
wire n_15752;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_3770;
wire n_9818;
wire n_2772;
wire n_7219;
wire n_6530;
wire n_9662;
wire n_12896;
wire n_4440;
wire n_15694;
wire n_8774;
wire n_4402;
wire n_14518;
wire n_10566;
wire n_927;
wire n_13397;
wire n_10178;
wire n_5052;
wire n_7299;
wire n_12367;
wire n_4541;
wire n_12104;
wire n_5009;
wire n_15360;
wire n_4872;
wire n_929;
wire n_6402;
wire n_12469;
wire n_13526;
wire n_9936;
wire n_12563;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_13132;
wire n_7326;
wire n_6609;
wire n_7243;
wire n_10115;
wire n_13321;
wire n_9530;
wire n_14692;
wire n_15042;
wire n_5326;
wire n_7471;
wire n_10455;
wire n_7067;
wire n_1183;
wire n_11778;
wire n_12793;
wire n_14722;
wire n_13427;
wire n_15488;
wire n_15519;
wire n_4627;
wire n_14835;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_15391;
wire n_9909;
wire n_11393;
wire n_14871;
wire n_12406;
wire n_8691;
wire n_8620;
wire n_14907;
wire n_3342;
wire n_6748;
wire n_15264;
wire n_7741;
wire n_998;
wire n_5035;
wire n_9466;
wire n_13270;
wire n_717;
wire n_11719;
wire n_7790;
wire n_6149;
wire n_10052;
wire n_10109;
wire n_1383;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_1424;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_15358;
wire n_1000;
wire n_11963;
wire n_12428;
wire n_14636;
wire n_9571;
wire n_8424;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_8026;
wire n_7528;
wire n_9470;
wire n_3810;
wire n_552;
wire n_4798;
wire n_9638;
wire n_2532;
wire n_15516;
wire n_1388;
wire n_3006;
wire n_216;
wire n_10265;
wire n_12655;
wire n_8174;
wire n_7941;
wire n_13524;
wire n_912;
wire n_11175;
wire n_13792;
wire n_5010;
wire n_15756;
wire n_11483;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_15067;
wire n_11995;
wire n_14378;
wire n_5089;
wire n_13356;
wire n_2849;
wire n_11371;
wire n_14912;
wire n_1201;
wire n_1398;
wire n_884;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_1395;
wire n_14191;
wire n_6264;
wire n_2199;
wire n_2661;
wire n_8861;
wire n_731;
wire n_5359;
wire n_13480;
wire n_8644;
wire n_1955;
wire n_8907;
wire n_931;
wire n_474;
wire n_312;
wire n_1791;
wire n_12304;
wire n_13571;
wire n_15156;
wire n_11080;
wire n_10984;
wire n_958;
wire n_5137;
wire n_6902;
wire n_3331;
wire n_5104;
wire n_14079;
wire n_10100;
wire n_15168;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_15411;
wire n_15743;
wire n_2773;
wire n_6205;
wire n_10906;
wire n_6380;
wire n_9441;
wire n_7478;
wire n_7913;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_589;
wire n_15144;
wire n_3606;
wire n_1310;
wire n_12692;
wire n_819;
wire n_13600;
wire n_13715;
wire n_1334;
wire n_3591;
wire n_7939;
wire n_13602;
wire n_2788;
wire n_964;
wire n_14224;
wire n_8503;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_14919;
wire n_6449;
wire n_2797;
wire n_6723;
wire n_9108;
wire n_7458;
wire n_9787;
wire n_10846;
wire n_7436;
wire n_6440;
wire n_4746;
wire n_13363;
wire n_15186;
wire n_14101;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_211;
wire n_2748;
wire n_9376;
wire n_5194;
wire n_9786;
wire n_14682;
wire n_1834;
wire n_8446;
wire n_14908;
wire n_9033;
wire n_2331;
wire n_13810;
wire n_14403;
wire n_12933;
wire n_2292;
wire n_7435;
wire n_12908;
wire n_15031;
wire n_3441;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_3534;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_13893;
wire n_3964;
wire n_12996;
wire n_2416;
wire n_311;
wire n_15171;
wire n_14201;
wire n_5947;
wire n_8923;
wire n_13625;
wire n_12643;
wire n_1877;
wire n_13315;
wire n_13473;
wire n_3944;
wire n_7685;
wire n_6124;
wire n_6736;
wire n_7363;
wire n_8192;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_14597;
wire n_5985;
wire n_8197;
wire n_556;
wire n_15663;
wire n_2209;
wire n_14353;
wire n_3605;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_1602;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_14950;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_3306;
wire n_12827;
wire n_12678;
wire n_13795;
wire n_276;
wire n_9115;
wire n_3026;
wire n_12235;
wire n_14547;
wire n_221;
wire n_4584;
wire n_15416;
wire n_3090;
wire n_5232;
wire n_11833;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_14386;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_9938;
wire n_11285;
wire n_12098;
wire n_8082;
wire n_4428;
wire n_8730;
wire n_1533;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_15533;
wire n_266;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_2274;
wire n_9203;
wire n_14415;
wire n_9977;
wire n_15073;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_15165;
wire n_5761;
wire n_13982;
wire n_13475;
wire n_518;
wire n_9242;
wire n_15079;
wire n_6773;
wire n_4618;
wire n_12611;
wire n_13859;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_4679;
wire n_13569;
wire n_1745;
wire n_914;
wire n_3479;
wire n_11262;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_12713;
wire n_317;
wire n_12880;
wire n_13144;
wire n_7455;
wire n_4805;
wire n_1679;
wire n_8651;
wire n_13959;
wire n_3454;
wire n_2160;
wire n_9141;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_2146;
wire n_6531;
wire n_10952;
wire n_2131;
wire n_488;
wire n_10851;
wire n_11027;
wire n_13628;
wire n_11852;
wire n_10660;
wire n_10221;
wire n_5472;
wire n_3547;
wire n_7430;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_11803;
wire n_15738;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_13685;
wire n_2575;
wire n_5100;
wire n_9286;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_1933;
wire n_8281;
wire n_10819;
wire n_1179;
wire n_324;
wire n_3816;
wire n_14693;
wire n_4807;
wire n_15613;
wire n_8842;
wire n_14786;
wire n_4411;
wire n_14521;
wire n_9184;
wire n_3214;
wire n_1243;
wire n_9704;
wire n_301;
wire n_2928;
wire n_13585;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_1917;
wire n_14486;
wire n_8024;
wire n_1580;
wire n_12562;
wire n_7730;
wire n_8814;
wire n_8530;
wire n_11428;
wire n_2822;
wire n_11592;
wire n_4180;
wire n_15090;
wire n_9193;
wire n_1281;
wire n_11677;
wire n_8467;
wire n_7281;
wire n_15385;
wire n_3109;
wire n_9717;
wire n_13577;
wire n_3354;
wire n_2572;
wire n_7711;
wire n_1520;
wire n_3126;
wire n_11090;
wire n_8984;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_9290;
wire n_6417;
wire n_351;
wire n_13281;
wire n_5740;
wire n_259;
wire n_1731;
wire n_13769;
wire n_14870;
wire n_5648;
wire n_5820;
wire n_13266;
wire n_13957;
wire n_14580;
wire n_15627;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_13672;
wire n_14028;
wire n_9875;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_858;
wire n_2049;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_14772;
wire n_8676;
wire n_956;
wire n_5534;
wire n_8003;
wire n_663;
wire n_4880;
wire n_13827;
wire n_8785;
wire n_9853;
wire n_13192;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_15681;
wire n_2781;
wire n_4126;
wire n_410;
wire n_14542;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_6556;
wire n_1594;
wire n_15048;
wire n_8692;
wire n_664;
wire n_1869;
wire n_6889;
wire n_9183;
wire n_7230;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_9778;
wire n_14326;
wire n_5196;
wire n_6199;
wire n_2016;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_15739;
wire n_10852;
wire n_15003;
wire n_4470;
wire n_14665;
wire n_6726;
wire n_12374;
wire n_13200;
wire n_9529;
wire n_580;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_8998;
wire n_465;
wire n_10538;
wire n_1790;
wire n_7011;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_4014;
wire n_13342;
wire n_4704;
wire n_11066;
wire n_341;
wire n_1744;
wire n_828;
wire n_10315;
wire n_2142;
wire n_4252;
wire n_607;
wire n_13886;
wire n_9123;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_2448;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_15545;
wire n_4048;
wire n_4596;
wire n_14924;
wire n_12368;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_3406;
wire n_820;
wire n_13193;
wire n_951;
wire n_12796;
wire n_6100;
wire n_6516;
wire n_952;
wire n_3919;
wire n_14489;
wire n_8462;
wire n_13774;
wire n_6977;
wire n_9380;
wire n_13847;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_12529;
wire n_2263;
wire n_15708;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_974;
wire n_6522;
wire n_8979;
wire n_14053;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_10514;
wire n_8930;
wire n_8429;
wire n_14581;
wire n_628;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_7890;
wire n_12785;
wire n_3973;
wire n_2756;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_9347;
wire n_6024;
wire n_807;
wire n_4761;
wire n_15312;
wire n_6675;
wire n_6270;
wire n_14155;
wire n_12461;
wire n_1275;
wire n_2884;
wire n_6808;
wire n_485;
wire n_13603;
wire n_1510;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_6207;
wire n_5783;
wire n_7006;
wire n_6931;
wire n_3120;
wire n_5821;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_238;
wire n_9082;
wire n_10925;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_202;
wire n_9879;
wire n_1749;
wire n_11158;
wire n_3474;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_2549;
wire n_4690;
wire n_11669;
wire n_14390;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_8264;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_12078;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_248;
wire n_2302;
wire n_8135;
wire n_10618;
wire n_15647;
wire n_1667;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_1037;
wire n_8545;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_3592;
wire n_11739;
wire n_468;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_10497;
wire n_14561;
wire n_9445;
wire n_14978;
wire n_2637;
wire n_1639;
wire n_7627;
wire n_13301;
wire n_183;
wire n_9803;
wire n_13293;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_3195;
wire n_466;
wire n_2526;
wire n_6346;
wire n_14381;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_15709;
wire n_15729;
wire n_8408;
wire n_12639;
wire n_3277;
wire n_14212;
wire n_2548;
wire n_5386;
wire n_991;
wire n_10661;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_3817;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_7811;
wire n_340;
wire n_13158;
wire n_1108;
wire n_14649;
wire n_11676;
wire n_11044;
wire n_14737;
wire n_11771;
wire n_12266;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_12175;
wire n_5003;
wire n_15530;
wire n_13536;
wire n_10512;
wire n_13833;
wire n_14714;
wire n_11384;
wire n_4827;
wire n_1601;
wire n_12287;
wire n_1960;
wire n_2694;
wire n_11679;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_1686;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_12353;
wire n_14441;
wire n_3042;
wire n_14129;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_12398;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_13485;
wire n_9087;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_9043;
wire n_6075;
wire n_12991;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_10789;
wire n_11134;
wire n_12705;
wire n_13735;
wire n_15333;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_11828;
wire n_14470;
wire n_12326;
wire n_15497;
wire n_1586;
wire n_14264;
wire n_7847;
wire n_8506;
wire n_14115;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_380;
wire n_13830;
wire n_13178;
wire n_6133;
wire n_3723;
wire n_11548;
wire n_13041;
wire n_1190;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_14184;
wire n_7822;
wire n_397;
wire n_4380;
wire n_6453;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_6127;
wire n_14183;
wire n_10762;
wire n_11452;
wire n_4398;
wire n_2498;
wire n_11342;
wire n_11362;
wire n_15734;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_14200;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_10797;
wire n_7289;
wire n_4193;
wire n_11266;
wire n_3570;
wire n_14110;
wire n_12309;
wire n_7926;
wire n_14806;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_12479;
wire n_172;
wire n_7354;
wire n_15568;
wire n_8352;
wire n_12502;
wire n_13824;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_10360;
wire n_239;
wire n_7960;
wire n_15620;
wire n_9450;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_5689;
wire n_13953;
wire n_7482;
wire n_1043;
wire n_12912;
wire n_14847;
wire n_10312;
wire n_4090;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_4165;
wire n_12454;
wire n_10480;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_9223;
wire n_8143;
wire n_13191;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_10131;
wire n_352;
wire n_12537;
wire n_6838;
wire n_15464;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_11988;
wire n_12600;
wire n_12921;
wire n_14536;
wire n_2169;
wire n_13226;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_13567;
wire n_1361;
wire n_6139;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_13686;
wire n_662;
wire n_6256;
wire n_7965;
wire n_13645;
wire n_15645;
wire n_3262;
wire n_6613;
wire n_11438;
wire n_11244;
wire n_4008;
wire n_12919;
wire n_3356;
wire n_14432;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_1642;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_3210;
wire n_6361;
wire n_937;
wire n_9880;
wire n_13253;
wire n_4689;
wire n_14321;
wire n_8183;
wire n_1682;
wire n_14981;
wire n_11348;
wire n_4547;
wire n_11245;
wire n_9685;
wire n_11685;
wire n_11169;
wire n_7474;
wire n_12422;
wire n_5731;
wire n_12467;
wire n_13354;
wire n_11607;
wire n_8650;
wire n_6085;
wire n_6329;
wire n_6678;
wire n_11546;
wire n_15259;
wire n_14654;
wire n_3329;
wire n_15460;
wire n_10503;
wire n_330;
wire n_8662;
wire n_14422;
wire n_15058;
wire n_9694;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_14664;
wire n_13215;
wire n_1406;
wire n_13400;
wire n_4601;
wire n_14971;
wire n_9905;
wire n_962;
wire n_9948;
wire n_10465;
wire n_14630;
wire n_12429;
wire n_10590;
wire n_3647;
wire n_3681;
wire n_13782;
wire n_14734;
wire n_15476;
wire n_14494;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_8526;
wire n_13331;
wire n_1186;
wire n_14956;
wire n_4623;
wire n_7325;
wire n_13751;
wire n_10887;
wire n_14866;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_14019;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_2518;
wire n_5883;
wire n_13743;
wire n_7166;
wire n_13812;
wire n_14970;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_13378;
wire n_3988;
wire n_6560;
wire n_14055;
wire n_11319;
wire n_1720;
wire n_3476;
wire n_7028;
wire n_4842;
wire n_204;
wire n_482;
wire n_7838;
wire n_9890;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_11492;
wire n_7873;
wire n_2688;
wire n_394;
wire n_1845;
wire n_1489;
wire n_6535;
wire n_12731;
wire n_12399;
wire n_942;
wire n_7518;
wire n_12342;
wire n_2798;
wire n_7414;
wire n_9744;
wire n_9817;
wire n_6147;
wire n_2852;
wire n_9199;
wire n_10063;
wire n_12640;
wire n_1524;
wire n_11160;
wire n_8973;
wire n_9548;
wire n_6448;
wire n_13544;
wire n_7791;
wire n_14292;
wire n_1964;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_1920;
wire n_2753;
wire n_12533;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_9862;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_1225;
wire n_12616;
wire n_11385;
wire n_1544;
wire n_1485;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_1846;
wire n_12535;
wire n_3437;
wire n_12178;
wire n_4111;
wire n_14375;
wire n_12653;
wire n_6643;
wire n_533;
wire n_12327;
wire n_7146;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_11346;
wire n_2506;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_14896;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_2626;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_14810;
wire n_9069;
wire n_13110;
wire n_15719;
wire n_14879;
wire n_3562;
wire n_5852;
wire n_14030;
wire n_2973;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_15164;
wire n_8249;
wire n_7052;
wire n_11343;
wire n_12348;
wire n_3665;
wire n_273;
wire n_10496;
wire n_3007;
wire n_12257;
wire n_3528;
wire n_15590;
wire n_15770;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_14149;
wire n_13394;
wire n_4571;
wire n_10843;
wire n_13391;
wire n_3698;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_13384;
wire n_3355;
wire n_14680;
wire n_2454;
wire n_8234;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_9960;
wire n_1066;
wire n_10997;
wire n_1948;
wire n_157;
wire n_4215;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_10998;
wire n_15422;
wire n_9003;
wire n_2154;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_1484;
wire n_12418;
wire n_14216;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_14837;
wire n_13498;
wire n_3752;
wire n_7312;
wire n_13263;
wire n_7919;
wire n_2283;
wire n_14877;
wire n_5145;
wire n_15203;
wire n_4219;
wire n_1229;
wire n_11269;
wire n_10800;
wire n_7085;
wire n_1373;
wire n_11491;
wire n_12065;
wire n_3958;
wire n_13950;
wire n_9341;
wire n_7848;
wire n_6939;
wire n_11408;
wire n_14048;
wire n_3985;
wire n_2427;
wire n_11772;
wire n_4196;
wire n_1447;
wire n_14103;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_13183;
wire n_6689;
wire n_13732;
wire n_14968;
wire n_10993;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12519;
wire n_9172;
wire n_12769;
wire n_14985;
wire n_15542;
wire n_14653;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_5149;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_2680;
wire n_11311;
wire n_10112;
wire n_14443;
wire n_1047;
wire n_10765;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_15263;
wire n_11792;
wire n_14285;
wire n_1385;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_9734;
wire n_502;
wire n_2668;
wire n_7288;
wire n_8558;
wire n_13242;
wire n_10489;
wire n_1257;
wire n_7707;
wire n_3197;
wire n_12421;
wire n_7223;
wire n_13282;
wire n_14436;
wire n_7833;
wire n_12113;
wire n_14868;
wire n_4987;
wire n_14599;
wire n_2128;
wire n_5512;
wire n_7274;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_14351;
wire n_3743;
wire n_6206;
wire n_9068;
wire n_13352;
wire n_8136;
wire n_834;
wire n_5033;
wire n_9808;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_14812;
wire n_3124;
wire n_10612;
wire n_11086;
wire n_1741;
wire n_7466;
wire n_1002;
wire n_6529;
wire n_10260;
wire n_11293;
wire n_1949;
wire n_14728;
wire n_3759;
wire n_545;
wire n_2671;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_12285;
wire n_2715;
wire n_1804;
wire n_13310;
wire n_11710;
wire n_8619;
wire n_251;
wire n_2508;
wire n_11568;
wire n_3511;
wire n_2054;
wire n_10253;
wire n_6290;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_1337;
wire n_9150;
wire n_10134;
wire n_14508;
wire n_15122;
wire n_11603;
wire n_13798;
wire n_1477;
wire n_7277;
wire n_6455;
wire n_15277;
wire n_15092;
wire n_13804;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_14778;
wire n_15714;
wire n_13099;
wire n_2614;
wire n_12015;
wire n_8146;
wire n_4492;
wire n_13690;
wire n_14822;
wire n_2833;
wire n_2758;
wire n_8813;
wire n_5607;
wire n_11562;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_10194;
wire n_14566;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_12157;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_13386;
wire n_13846;
wire n_8910;
wire n_12311;
wire n_4376;
wire n_6203;
wire n_1001;
wire n_6408;
wire n_14374;
wire n_2241;
wire n_9448;
wire n_13064;
wire n_7683;
wire n_10739;
wire n_14815;
wire n_6555;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_4708;
wire n_13619;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_12031;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_8643;
wire n_1076;
wire n_15660;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_15357;
wire n_1378;
wire n_855;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_1377;
wire n_11718;
wire n_10821;
wire n_8565;
wire n_13648;
wire n_14831;
wire n_14996;
wire n_11170;
wire n_695;
wire n_11758;
wire n_12126;
wire n_14383;
wire n_8550;
wire n_14543;
wire n_4081;
wire n_1542;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_14450;
wire n_14747;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_15722;
wire n_14683;
wire n_10599;
wire n_9667;
wire n_14192;
wire n_14181;
wire n_6401;
wire n_7322;
wire n_1716;
wire n_278;
wire n_15278;
wire n_9053;
wire n_11658;
wire n_15504;
wire n_11893;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_13492;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_14001;
wire n_14213;
wire n_5562;
wire n_15397;
wire n_3303;
wire n_978;
wire n_4324;
wire n_7051;
wire n_10850;
wire n_384;
wire n_9185;
wire n_8477;
wire n_1976;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_4382;
wire n_12195;
wire n_13376;
wire n_14842;
wire n_2905;
wire n_13115;
wire n_1291;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_749;
wire n_13864;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_11601;
wire n_13289;
wire n_15279;
wire n_11971;
wire n_13182;
wire n_2122;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_9919;
wire n_3160;
wire n_12135;
wire n_1065;
wire n_6574;
wire n_11116;
wire n_13324;
wire n_12604;
wire n_6571;
wire n_13305;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_1255;
wire n_568;
wire n_8876;
wire n_15215;
wire n_5124;
wire n_143;
wire n_9151;
wire n_3951;
wire n_8829;
wire n_823;
wire n_7824;
wire n_9359;
wire n_13381;
wire n_1074;
wire n_698;
wire n_13236;
wire n_3569;
wire n_14189;
wire n_739;
wire n_14299;
wire n_7094;
wire n_3874;
wire n_15761;
wire n_2528;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8971;
wire n_8140;
wire n_15111;
wire n_8060;
wire n_1338;
wire n_1097;
wire n_10558;
wire n_3027;
wire n_781;
wire n_4083;
wire n_7036;
wire n_9579;
wire n_11124;
wire n_9475;
wire n_15273;
wire n_6392;
wire n_1810;
wire n_182;
wire n_5915;
wire n_8527;
wire n_573;
wire n_12899;
wire n_13777;
wire n_15301;
wire n_9049;
wire n_7351;
wire n_1583;
wire n_13718;
wire n_4480;
wire n_1730;
wire n_9352;
wire n_2295;
wire n_2746;
wire n_389;
wire n_814;
wire n_14775;
wire n_7608;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_6260;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_13202;
wire n_7909;
wire n_15350;
wire n_7413;
wire n_13638;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_14392;
wire n_222;
wire n_11340;
wire n_15759;
wire n_10734;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_15383;
wire n_11903;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_13279;
wire n_13644;
wire n_6912;
wire n_11560;
wire n_721;
wire n_10395;
wire n_1461;
wire n_742;
wire n_7175;
wire n_691;
wire n_3617;
wire n_8276;
wire n_10330;
wire n_2076;
wire n_13291;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_14966;
wire n_3567;
wire n_11465;
wire n_377;
wire n_1598;
wire n_7524;
wire n_15255;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_11564;
wire n_14015;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_11265;
wire n_9370;
wire n_11125;
wire n_918;
wire n_13136;
wire n_9670;
wire n_1114;
wire n_13513;
wire n_763;
wire n_4027;
wire n_12916;
wire n_3154;
wire n_9334;
wire n_7783;
wire n_13220;
wire n_15131;
wire n_6692;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_10276;
wire n_14322;
wire n_12331;
wire n_3520;
wire n_191;
wire n_8978;
wire n_10594;
wire n_12531;
wire n_8093;
wire n_8245;
wire n_15072;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_12521;
wire n_11302;
wire n_946;
wire n_12910;
wire n_13349;
wire n_9956;
wire n_1303;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_15509;
wire n_2881;
wire n_11745;
wire n_1116;
wire n_10098;
wire n_1570;
wire n_1702;
wire n_8891;
wire n_15240;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_11690;
wire n_9487;
wire n_1780;
wire n_3897;
wire n_11707;
wire n_1689;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_7697;
wire n_14608;
wire n_1944;
wire n_6403;
wire n_15564;
wire n_7306;
wire n_13835;
wire n_1347;
wire n_7947;
wire n_795;
wire n_10118;
wire n_1221;
wire n_14350;
wire n_7547;
wire n_7470;
wire n_6013;
wire n_13815;
wire n_7733;
wire n_13800;
wire n_1245;
wire n_7693;
wire n_9557;
wire n_3215;
wire n_6491;
wire n_448;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_14039;
wire n_14072;
wire n_15662;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_1561;
wire n_13039;
wire n_13773;
wire n_13130;
wire n_14109;
wire n_8582;
wire n_10441;
wire n_1112;
wire n_5518;
wire n_6982;
wire n_10002;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_6661;
wire n_9124;
wire n_234;
wire n_6293;
wire n_15375;
wire n_15671;
wire n_5847;
wire n_13719;
wire n_7345;
wire n_6049;
wire n_1460;
wire n_911;
wire n_8847;
wire n_9762;
wire n_11242;
wire n_8957;
wire n_14136;
wire n_10923;
wire n_7385;
wire n_14548;
wire n_5159;
wire n_2862;
wire n_472;
wire n_15793;
wire n_2615;
wire n_4068;
wire n_6558;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_2474;
wire n_3703;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_13694;
wire n_2444;
wire n_2437;
wire n_12313;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_2267;
wire n_9543;
wire n_3035;
wire n_13688;
wire n_14661;
wire n_668;
wire n_4166;
wire n_11396;
wire n_8356;
wire n_1821;
wire n_6136;
wire n_9660;
wire n_15196;
wire n_11443;
wire n_9483;
wire n_1058;
wire n_3378;
wire n_15765;
wire n_6855;
wire n_15305;
wire n_15588;
wire n_3745;
wire n_14754;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_4188;
wire n_15020;
wire n_13467;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_13093;
wire n_13062;
wire n_9328;
wire n_14252;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_14130;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_14930;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_6312;
wire n_11532;
wire n_2505;
wire n_9539;
wire n_334;
wire n_4817;
wire n_6668;
wire n_8747;
wire n_9415;
wire n_15274;
wire n_4115;
wire n_2999;
wire n_14343;
wire n_15548;
wire n_2014;
wire n_9385;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_9147;
wire n_470;
wire n_11209;
wire n_7653;
wire n_13462;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_2408;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_14276;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_13752;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_13185;
wire n_6340;
wire n_9027;
wire n_1972;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_4383;
wire n_13596;
wire n_6995;
wire n_10902;
wire n_4491;
wire n_12889;
wire n_13855;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_455;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_363;
wire n_12250;
wire n_4486;
wire n_10420;
wire n_9515;
wire n_6971;
wire n_1816;
wire n_11304;
wire n_9642;
wire n_393;
wire n_503;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_15232;
wire n_3024;
wire n_7475;
wire n_10485;
wire n_14231;
wire n_12105;
wire n_4612;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_13219;
wire n_14329;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_9079;
wire n_15544;
wire n_15721;
wire n_9382;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_307;
wire n_10444;
wire n_4529;
wire n_500;
wire n_3361;
wire n_11377;
wire n_714;
wire n_3478;
wire n_8018;
wire n_8653;
wire n_13295;
wire n_15142;
wire n_3936;
wire n_1349;
wire n_291;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_2723;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_5823;
wire n_7305;
wire n_13388;
wire n_2800;
wire n_3496;
wire n_13160;
wire n_13731;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_15249;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_14550;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_14503;
wire n_4390;
wire n_12248;
wire n_13818;
wire n_15024;
wire n_3096;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_15346;
wire n_2651;
wire n_13477;
wire n_8884;
wire n_8803;
wire n_14886;
wire n_2095;
wire n_3239;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_10978;
wire n_8222;
wire n_13808;
wire n_14644;
wire n_6822;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_11715;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_1998;
wire n_9706;
wire n_1574;
wire n_3101;
wire n_15174;
wire n_15454;
wire n_240;
wire n_10642;
wire n_15213;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_12181;
wire n_10187;
wire n_3374;
wire n_10387;
wire n_11014;
wire n_13764;
wire n_14560;
wire n_15033;
wire n_2640;
wire n_253;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_11864;
wire n_14829;
wire n_3876;
wire n_11007;
wire n_11224;
wire n_15473;
wire n_249;
wire n_11006;
wire n_15584;
wire n_9564;
wire n_15018;
wire n_3125;
wire n_7391;
wire n_8790;
wire n_15569;
wire n_9230;
wire n_6617;
wire n_4293;
wire n_10219;
wire n_941;
wire n_3552;
wire n_1031;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_15193;
wire n_849;
wire n_4684;
wire n_3116;
wire n_9591;
wire n_14067;
wire n_6407;
wire n_6429;
wire n_4091;
wire n_14108;
wire n_1753;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_14833;
wire n_10364;
wire n_15439;
wire n_2471;
wire n_10479;
wire n_11422;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_13660;
wire n_8398;
wire n_4412;
wire n_14480;
wire n_2807;
wire n_8178;
wire n_13970;
wire n_6801;
wire n_15247;
wire n_1921;
wire n_12489;
wire n_8491;
wire n_14000;
wire n_14372;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_5630;
wire n_4758;
wire n_4781;
wire n_10065;
wire n_12046;
wire n_10212;
wire n_9283;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_12030;
wire n_12738;
wire n_13408;
wire n_206;
wire n_4057;
wire n_15062;
wire n_633;
wire n_1170;
wire n_15248;
wire n_13727;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_308;
wire n_10268;
wire n_15236;
wire n_3444;
wire n_1040;
wire n_14801;
wire n_3059;
wire n_6113;
wire n_9468;
wire n_12601;
wire n_10070;
wire n_14098;
wire n_14482;
wire n_15399;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_13641;
wire n_2634;
wire n_1761;
wire n_14223;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_1890;
wire n_3017;
wire n_14947;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_14983;
wire n_14748;
wire n_10559;
wire n_2308;
wire n_2333;
wire n_13173;
wire n_8439;
wire n_3001;
wire n_9641;
wire n_1089;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_15355;
wire n_15669;
wire n_12059;
wire n_12488;
wire n_3795;
wire n_7321;
wire n_14848;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_8200;
wire n_11110;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_15001;
wire n_8304;
wire n_3896;
wire n_3815;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_3274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_13328;
wire n_7537;
wire n_10516;
wire n_4093;
wire n_1616;
wire n_8675;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_10892;
wire n_339;
wire n_434;
wire n_10493;
wire n_13542;
wire n_288;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_15037;
wire n_4794;
wire n_15130;
wire n_722;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_14604;
wire n_14735;
wire n_2223;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_629;
wire n_1621;
wire n_9016;
wire n_2547;
wire n_14426;
wire n_2415;
wire n_13101;
wire n_11887;
wire n_15456;
wire n_14349;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_11545;
wire n_9729;
wire n_5073;
wire n_12691;
wire n_827;
wire n_8846;
wire n_8315;
wire n_12471;
wire n_11033;
wire n_12451;
wire n_4834;
wire n_11040;
wire n_12665;
wire n_11850;
wire n_11754;
wire n_14916;
wire n_15740;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_14356;
wire n_4762;
wire n_192;
wire n_5581;
wire n_13748;
wire n_9029;
wire n_11672;
wire n_9411;
wire n_3113;
wire n_10353;
wire n_6837;
wire n_992;
wire n_3813;
wire n_3660;
wire n_10847;
wire n_12651;
wire n_3766;
wire n_1613;
wire n_10451;
wire n_11043;
wire n_1458;
wire n_15801;
wire n_5303;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_9414;
wire n_1027;
wire n_3266;
wire n_7023;
wire n_3574;
wire n_9615;
wire n_12003;
wire n_14205;
wire n_7496;
wire n_1189;
wire n_11277;
wire n_14564;
wire n_223;
wire n_4154;
wire n_12165;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_10866;
wire n_14190;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_365;
wire n_3844;
wire n_8777;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_11061;
wire n_11763;
wire n_15546;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_11534;
wire n_10653;
wire n_11587;
wire n_6373;
wire n_5375;
wire n_12280;
wire n_13461;
wire n_12492;
wire n_9221;
wire n_13581;
wire n_14344;
wire n_15742;
wire n_2451;
wire n_12972;
wire n_5370;
wire n_13789;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_9811;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_509;
wire n_13188;
wire n_4819;
wire n_14511;
wire n_1209;
wire n_7906;
wire n_13286;
wire n_5248;
wire n_9951;
wire n_1708;
wire n_7131;
wire n_805;
wire n_14723;
wire n_396;
wire n_6411;
wire n_350;
wire n_2051;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_14488;
wire n_11032;
wire n_2359;
wire n_5112;
wire n_13582;
wire n_480;
wire n_142;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_10507;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_11843;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_14614;
wire n_13531;
wire n_7797;
wire n_3668;
wire n_11335;
wire n_11629;
wire n_15147;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_13880;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_13988;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_7582;
wire n_15272;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_13609;
wire n_3487;
wire n_14587;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_287;
wire n_4302;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_6534;
wire n_3340;
wire n_10614;
wire n_230;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_13679;
wire n_461;
wire n_873;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_2989;
wire n_5778;
wire n_11257;
wire n_8425;
wire n_15176;
wire n_8087;
wire n_13276;
wire n_9910;
wire n_3395;
wire n_7607;
wire n_7060;
wire n_10217;
wire n_14458;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_11801;
wire n_13217;
wire n_2513;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_10743;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_250;
wire n_1711;
wire n_13424;
wire n_14658;
wire n_15066;
wire n_4884;
wire n_14830;
wire n_14397;
wire n_10853;
wire n_1579;
wire n_7867;
wire n_9651;
wire n_3275;
wire n_13565;
wire n_14281;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_836;
wire n_6135;
wire n_13802;
wire n_14594;
wire n_15474;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_10338;
wire n_9246;
wire n_15316;
wire n_522;
wire n_10270;
wire n_3678;
wire n_6814;
wire n_11115;
wire n_3440;
wire n_10557;
wire n_8669;
wire n_12978;
wire n_13784;
wire n_8001;
wire n_2094;
wire n_7525;
wire n_13468;
wire n_1511;
wire n_2356;
wire n_7257;
wire n_12363;
wire n_9372;
wire n_7553;
wire n_1422;
wire n_7529;
wire n_1772;
wire n_15668;
wire n_4692;
wire n_6791;
wire n_616;
wire n_15137;
wire n_14233;
wire n_8496;
wire n_3165;
wire n_11915;
wire n_13704;
wire n_1119;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_1433;
wire n_14976;
wire n_1902;
wire n_1842;
wire n_11788;
wire n_1620;
wire n_2739;
wire n_12544;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_13036;
wire n_3750;
wire n_14146;
wire n_1313;
wire n_3607;
wire n_7650;
wire n_12476;
wire n_13199;
wire n_3316;
wire n_8568;
wire n_516;
wire n_6903;
wire n_2418;
wire n_2864;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_4311;
wire n_12023;
wire n_1180;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_13413;
wire n_9486;
wire n_6450;
wire n_13002;
wire n_9544;
wire n_3261;
wire n_15153;
wire n_666;
wire n_12632;
wire n_12620;
wire n_9831;
wire n_7520;
wire n_13203;
wire n_13868;
wire n_4187;
wire n_6309;
wire n_940;
wire n_7903;
wire n_9697;
wire n_2058;
wire n_11303;
wire n_405;
wire n_213;
wire n_2660;
wire n_11877;
wire n_6733;
wire n_14462;
wire n_8864;
wire n_8456;
wire n_7384;
wire n_5317;
wire n_13285;
wire n_1094;
wire n_5430;
wire n_8610;
wire n_5942;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_9902;
wire n_494;
wire n_14933;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_15521;
wire n_3532;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_9039;
wire n_12598;
wire n_11854;
wire n_13374;
wire n_12416;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_2124;
wire n_8265;
wire n_4619;
wire n_381;
wire n_7639;
wire n_8704;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_11609;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_13230;
wire n_9294;
wire n_5036;
wire n_12811;
wire n_4221;
wire n_3297;
wire n_12186;
wire n_11747;
wire n_12494;
wire n_6395;
wire n_10327;
wire n_13032;
wire n_13826;
wire n_6179;
wire n_976;
wire n_7054;
wire n_7605;
wire n_3067;
wire n_11556;
wire n_15140;
wire n_2155;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_11529;
wire n_2686;
wire n_5327;
wire n_10021;
wire n_13684;
wire n_14199;
wire n_9146;
wire n_2364;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_14027;
wire n_2996;
wire n_15108;
wire n_15753;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_3803;
wire n_2085;
wire n_8941;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_10075;
wire n_9073;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_13750;
wire n_6171;
wire n_8775;
wire n_14104;
wire n_808;
wire n_12272;
wire n_9302;
wire n_5519;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_14684;
wire n_11895;
wire n_13458;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_15713;
wire n_1193;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_3412;
wire n_8279;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_12191;
wire n_9580;
wire n_8019;
wire n_14572;
wire n_13963;
wire n_9972;
wire n_3791;
wire n_13003;
wire n_6083;
wire n_13091;
wire n_12909;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_551;
wire n_699;
wire n_4320;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_3884;
wire n_9465;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_451;
wire n_11137;
wire n_8390;
wire n_8898;
wire n_13811;
wire n_14316;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_13839;
wire n_757;
wire n_594;
wire n_6120;
wire n_2190;
wire n_5231;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_14011;
wire n_8521;
wire n_3438;
wire n_166;
wire n_4141;
wire n_13954;
wire n_10436;
wire n_8464;
wire n_15701;
wire n_6547;
wire n_12794;
wire n_8799;
wire n_5193;
wire n_6423;
wire n_15496;
wire n_9442;
wire n_2850;
wire n_572;
wire n_6342;
wire n_6641;
wire n_1481;
wire n_15260;
wire n_6984;
wire n_1441;
wire n_15612;
wire n_3373;
wire n_5789;
wire n_15104;
wire n_10763;
wire n_2104;
wire n_7441;
wire n_9957;
wire n_513;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_12112;
wire n_13060;
wire n_14689;
wire n_3883;
wire n_10245;
wire n_14132;
wire n_10905;
wire n_5961;
wire n_261;
wire n_11235;
wire n_9449;
wire n_14817;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_6687;
wire n_9313;
wire n_5822;
wire n_9173;
wire n_433;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_15055;
wire n_3949;
wire n_5726;
wire n_9563;
wire n_11015;
wire n_14087;
wire n_2792;
wire n_9160;
wire n_15705;
wire n_219;
wire n_5364;
wire n_9974;
wire n_12129;
wire n_14753;
wire n_11166;
wire n_3315;
wire n_7031;
wire n_9285;
wire n_13658;
wire n_263;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_788;
wire n_9631;
wire n_14671;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_15172;
wire n_14751;
wire n_329;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_14438;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_4720;
wire n_10784;
wire n_12202;
wire n_4893;
wire n_14674;
wire n_3857;
wire n_13836;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_243;
wire n_12815;
wire n_1873;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_1866;
wire n_9945;
wire n_8661;
wire n_12431;
wire n_2130;
wire n_7424;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_7523;
wire n_2228;
wire n_8654;
wire n_5039;
wire n_11855;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_14229;
wire n_15060;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_15115;
wire n_15520;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_3099;
wire n_11156;
wire n_8531;
wire n_14188;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_4468;
wire n_13799;
wire n_5718;
wire n_4161;
wire n_6459;
wire n_1663;
wire n_6505;
wire n_12333;
wire n_12636;
wire n_8609;
wire n_13854;
wire n_8379;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_7626;
wire n_13576;
wire n_15380;
wire n_13100;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_1107;
wire n_12334;
wire n_2457;
wire n_3294;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_9209;
wire n_7311;
wire n_3686;
wire n_7669;
wire n_11218;
wire n_4502;
wire n_12119;
wire n_11787;
wire n_12618;
wire n_5958;
wire n_8793;
wire n_12355;
wire n_8103;
wire n_15052;
wire n_318;
wire n_9838;
wire n_2971;
wire n_1713;
wire n_9767;
wire n_10195;
wire n_715;
wire n_13722;
wire n_4277;
wire n_4526;
wire n_9300;
wire n_1265;
wire n_11500;
wire n_3490;
wire n_4849;
wire n_12943;
wire n_530;
wire n_15129;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_14306;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_11891;
wire n_8367;
wire n_618;
wire n_7367;
wire n_199;
wire n_14752;
wire n_5792;
wire n_11021;
wire n_3581;
wire n_12401;
wire n_8543;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_14897;
wire n_15447;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_6905;
wire n_10243;
wire n_612;
wire n_9700;
wire n_10564;
wire n_13829;
wire n_3725;
wire n_8682;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_3933;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_1175;
wire n_7244;
wire n_10745;
wire n_7368;
wire n_2311;
wire n_429;
wire n_1012;
wire n_3691;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_903;
wire n_7633;
wire n_13937;
wire n_4146;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_1802;
wire n_1504;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_286;
wire n_11509;
wire n_8640;
wire n_254;
wire n_14359;
wire n_8063;
wire n_15141;
wire n_3961;
wire n_11960;
wire n_4855;
wire n_12599;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_7878;
wire n_9514;
wire n_6803;
wire n_12411;
wire n_6186;
wire n_816;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_1188;
wire n_12465;
wire n_10605;
wire n_7427;
wire n_2206;
wire n_4004;
wire n_11029;
wire n_13532;
wire n_2967;
wire n_14013;
wire n_13250;
wire n_13118;
wire n_14419;
wire n_5404;
wire n_9933;
wire n_11449;
wire n_2916;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_4292;
wire n_9892;
wire n_15251;
wire n_8570;
wire n_6163;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_2467;
wire n_5549;
wire n_9408;
wire n_267;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_10163;
wire n_10454;
wire n_3983;
wire n_15401;
wire n_13339;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_12568;
wire n_3280;
wire n_13478;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_12970;
wire n_1515;
wire n_8916;
wire n_8902;
wire n_961;
wire n_14295;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_593;
wire n_8843;
wire n_9891;
wire n_10146;
wire n_12959;
wire n_9946;
wire n_7128;
wire n_14367;
wire n_637;
wire n_2377;
wire n_701;
wire n_6849;
wire n_9885;
wire n_7594;
wire n_950;
wire n_12330;
wire n_13915;
wire n_8129;
wire n_8162;
wire n_14890;
wire n_14819;
wire n_15057;
wire n_13906;
wire n_7457;
wire n_10643;
wire n_8744;
wire n_3009;
wire n_10504;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_13783;
wire n_6760;
wire n_10701;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_13664;
wire n_13987;
wire n_14265;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_3889;
wire n_13566;
wire n_15626;
wire n_2687;
wire n_12591;
wire n_12466;
wire n_1630;
wire n_2887;
wire n_15775;
wire n_9509;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_13416;
wire n_2194;
wire n_12798;
wire n_14885;
wire n_2619;
wire n_5329;
wire n_9015;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_9925;
wire n_10874;
wire n_6825;
wire n_1987;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_11831;
wire n_13726;
wire n_507;
wire n_9628;
wire n_968;
wire n_14399;
wire n_7767;
wire n_14412;
wire n_8294;
wire n_2271;
wire n_1008;
wire n_12279;
wire n_12243;
wire n_9419;
wire n_6611;
wire n_8562;
wire n_2583;
wire n_4560;
wire n_13705;
wire n_12614;
wire n_11378;
wire n_2606;
wire n_4899;
wire n_10250;
wire n_14631;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_10032;
wire n_10592;
wire n_11433;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_2391;
wire n_14063;
wire n_304;
wire n_2431;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_13425;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_7744;
wire n_2078;
wire n_7021;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_10595;
wire n_13591;
wire n_7748;
wire n_8537;
wire n_3450;
wire n_6827;
wire n_10126;
wire n_14421;
wire n_12041;
wire n_449;
wire n_4663;
wire n_11713;
wire n_2893;
wire n_11073;
wire n_13653;
wire n_1208;
wire n_15586;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_12566;
wire n_12931;
wire n_2728;
wire n_15525;
wire n_1072;
wire n_815;
wire n_13680;
wire n_6227;
wire n_7215;
wire n_15157;
wire n_7485;
wire n_3421;
wire n_13074;
wire n_9066;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_14332;
wire n_10302;
wire n_11974;
wire n_1067;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_3405;
wire n_14920;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_14716;
wire n_255;
wire n_10645;
wire n_13058;
wire n_15313;
wire n_284;
wire n_1952;
wire n_5074;
wire n_10604;
wire n_11096;
wire n_12036;
wire n_12876;
wire n_15286;
wire n_4044;
wire n_6564;
wire n_3436;
wire n_11161;
wire n_9671;
wire n_8782;
wire n_8709;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_14698;
wire n_2631;
wire n_12911;
wire n_289;
wire n_15715;
wire n_12491;
wire n_14994;
wire n_3937;
wire n_6468;
wire n_10080;
wire n_11216;
wire n_14368;
wire n_12228;
wire n_10570;
wire n_1293;
wire n_9857;
wire n_3159;
wire n_4701;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_14323;
wire n_794;
wire n_12929;
wire n_10882;
wire n_727;
wire n_894;
wire n_685;
wire n_9338;
wire n_13071;
wire n_353;
wire n_6857;
wire n_3240;
wire n_8144;
wire n_15075;
wire n_12261;
wire n_3576;
wire n_10435;
wire n_1863;
wire n_9542;
wire n_12536;
wire n_3385;
wire n_10921;
wire n_10795;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_12106;
wire n_12061;
wire n_3293;
wire n_872;
wire n_3922;
wire n_15116;
wire n_14585;
wire n_11085;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_7925;
wire n_7068;
wire n_7186;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_10609;
wire n_11157;
wire n_13649;
wire n_13739;
wire n_4991;
wire n_14804;
wire n_5594;
wire n_15126;
wire n_2554;
wire n_12291;
wire n_14510;
wire n_9097;
wire n_5422;
wire n_12124;
wire n_6871;
wire n_11755;
wire n_1513;
wire n_9783;
wire n_13806;
wire n_14364;
wire n_9510;
wire n_15472;
wire n_9389;
wire n_1913;
wire n_12074;
wire n_4934;
wire n_13497;
wire n_9404;
wire n_15406;
wire n_837;
wire n_8357;
wire n_10912;
wire n_6904;
wire n_5087;
wire n_14396;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_13234;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_9314;
wire n_11918;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_14466;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_14473;
wire n_12887;
wire n_2590;
wire n_5551;
wire n_7652;
wire n_3150;
wire n_10220;
wire n_8701;
wire n_10341;
wire n_11347;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_10550;
wire n_6499;
wire n_7830;
wire n_14673;
wire n_4011;
wire n_5131;
wire n_12217;
wire n_12365;
wire n_1959;
wire n_3133;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_13738;
wire n_13851;
wire n_9679;
wire n_14972;
wire n_765;
wire n_1492;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_14138;
wire n_13272;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_8712;
wire n_10232;
wire n_4058;
wire n_14113;
wire n_10461;
wire n_631;
wire n_14586;
wire n_8289;
wire n_11178;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_8591;
wire n_7966;
wire n_5059;
wire n_156;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_843;
wire n_8824;
wire n_11673;
wire n_2604;
wire n_2407;
wire n_14938;
wire n_1277;
wire n_14784;
wire n_2816;
wire n_11432;
wire n_14641;
wire n_14179;
wire n_14031;
wire n_7191;
wire n_14979;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_10412;
wire n_5242;
wire n_15433;
wire n_10326;
wire n_12650;
wire n_5219;
wire n_8417;
wire n_2675;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_3537;
wire n_10499;
wire n_8340;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_12487;
wire n_12658;
wire n_14324;
wire n_614;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_2119;
wire n_13613;
wire n_14740;
wire n_947;
wire n_9210;
wire n_12185;
wire n_1117;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_6893;
wire n_7406;
wire n_8681;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_3223;
wire n_10617;
wire n_12704;
wire n_12271;
wire n_3140;
wire n_7807;
wire n_3185;
wire n_4749;
wire n_9592;
wire n_2605;
wire n_5155;
wire n_14198;
wire n_7680;
wire n_9180;
wire n_14846;
wire n_15190;
wire n_10922;
wire n_10544;
wire n_12958;
wire n_926;
wire n_13030;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_12056;
wire n_14539;
wire n_1698;
wire n_15094;
wire n_8106;
wire n_9502;
wire n_4100;
wire n_13821;
wire n_6447;
wire n_13712;
wire n_4264;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_3788;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_777;
wire n_6422;
wire n_1299;
wire n_13896;
wire n_14761;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_3837;
wire n_2718;
wire n_15243;
wire n_1436;
wire n_14420;
wire n_1384;
wire n_11087;
wire n_15041;
wire n_11477;
wire n_3325;
wire n_2238;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_4085;
wire n_13299;
wire n_15393;
wire n_13243;
wire n_4464;
wire n_14314;
wire n_8612;
wire n_13042;
wire n_14144;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_15658;
wire n_10095;
wire n_14227;
wire n_4659;
wire n_13725;
wire n_10309;
wire n_3600;
wire n_6741;
wire n_11773;
wire n_12608;
wire n_8459;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_14164;
wire n_8268;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_10050;
wire n_6650;
wire n_8221;
wire n_9871;
wire n_11682;
wire n_7066;
wire n_15595;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_796;
wire n_1195;
wire n_7789;
wire n_13197;
wire n_10306;
wire n_15081;
wire n_184;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_1811;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_7193;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_11919;
wire n_14860;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_10450;
wire n_623;
wire n_1048;
wire n_5721;
wire n_11414;
wire n_11472;
wire n_3638;
wire n_9114;
wire n_11978;
wire n_4816;
wire n_12520;
wire n_10529;
wire n_8515;
wire n_2110;
wire n_13632;
wire n_5719;
wire n_1502;
wire n_14685;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_8812;
wire n_14505;
wire n_14892;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_3451;
wire n_9392;
wire n_13148;
wire n_1418;
wire n_10429;
wire n_1250;
wire n_292;
wire n_4937;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_14531;
wire n_3615;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_11538;
wire n_3072;
wire n_3087;
wire n_10037;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_12808;
wire n_13871;
wire n_4222;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_13435;
wire n_4401;
wire n_889;
wire n_15408;
wire n_12744;
wire n_2710;
wire n_6064;
wire n_15173;
wire n_11136;
wire n_9903;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_13801;
wire n_5793;
wire n_477;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_15480;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_10179;
wire n_11539;
wire n_4976;
wire n_12143;
wire n_9228;
wire n_2389;
wire n_9499;
wire n_7710;
wire n_11899;
wire n_7892;
wire n_2132;
wire n_2892;
wire n_13168;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_13879;
wire n_14038;
wire n_14771;
wire n_9522;
wire n_1564;
wire n_5578;
wire n_15617;
wire n_15463;
wire n_11215;
wire n_4658;
wire n_231;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_11076;
wire n_1457;
wire n_11890;
wire n_505;
wire n_9366;
wire n_14339;
wire n_14253;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_1787;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_537;
wire n_1993;
wire n_11806;
wire n_2281;
wire n_11054;
wire n_9148;
wire n_8406;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_10754;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_11050;
wire n_3705;
wire n_3211;
wire n_12443;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_11683;
wire n_8554;
wire n_546;
wire n_10920;
wire n_9275;
wire n_386;
wire n_10223;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_8896;
wire n_14398;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_11484;
wire n_7206;
wire n_4223;
wire n_11126;
wire n_7538;
wire n_2387;
wire n_5674;
wire n_12934;
wire n_15758;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_2846;
wire n_13598;
wire n_5282;
wire n_970;
wire n_10295;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_9409;
wire n_6799;
wire n_2237;
wire n_1060;
wire n_10336;
wire n_1951;
wire n_10228;
wire n_444;
wire n_12555;
wire n_4362;
wire n_1252;
wire n_3913;
wire n_3311;
wire n_1223;
wire n_7716;
wire n_6487;
wire n_11646;
wire n_511;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_8818;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_4348;
wire n_12980;
wire n_13966;
wire n_9881;
wire n_12530;
wire n_5013;
wire n_1597;
wire n_6807;
wire n_9463;
wire n_8954;
wire n_12212;
wire n_4489;
wire n_4839;
wire n_7251;
wire n_7254;
wire n_10466;
wire n_2596;
wire n_12973;
wire n_3163;
wire n_7540;
wire n_775;
wire n_11953;
wire n_4404;
wire n_13123;
wire n_14669;
wire n_1153;
wire n_5589;
wire n_439;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_13231;
wire n_12624;
wire n_1531;
wire n_7882;
wire n_2828;
wire n_453;
wire n_8552;
wire n_10425;
wire n_7554;
wire n_2384;
wire n_8069;
wire n_13165;
wire n_4261;
wire n_4204;
wire n_10848;
wire n_7558;
wire n_8373;
wire n_759;
wire n_2724;
wire n_426;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_11482;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_12151;
wire n_4006;
wire n_15201;
wire n_2226;
wire n_11089;
wire n_2801;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_13422;
wire n_15204;
wire n_6384;
wire n_1901;
wire n_3869;
wire n_7421;
wire n_15579;
wire n_2556;
wire n_13828;
wire n_10166;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_1647;
wire n_14702;
wire n_13179;
wire n_14562;
wire n_15585;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_12033;
wire n_1892;
wire n_1614;
wire n_11839;
wire n_3742;
wire n_9844;
wire n_3683;
wire n_12826;
wire n_4801;
wire n_8318;
wire n_14376;
wire n_13834;
wire n_401;
wire n_3260;
wire n_10366;
wire n_2550;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_11365;
wire n_3175;
wire n_9595;
wire n_7188;
wire n_15015;
wire n_3736;
wire n_5475;
wire n_11217;
wire n_15651;
wire n_15555;
wire n_15341;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_13923;
wire n_1096;
wire n_9287;
wire n_7991;
wire n_15477;
wire n_13051;
wire n_6233;
wire n_2227;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_14991;
wire n_14686;
wire n_3284;
wire n_12214;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_427;
wire n_13330;
wire n_8926;
wire n_6257;
wire n_2159;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_4386;
wire n_10361;
wire n_11228;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_13924;
wire n_4955;
wire n_8965;
wire n_11290;
wire n_4149;
wire n_5936;
wire n_12518;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_501;
wire n_2276;
wire n_3234;
wire n_9052;
wire n_13476;
wire n_14047;
wire n_856;
wire n_2803;
wire n_8817;
wire n_379;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_11488;
wire n_13671;
wire n_12162;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_6587;
wire n_14627;
wire n_1129;
wire n_14876;
wire n_6987;
wire n_7781;
wire n_602;
wire n_7360;
wire n_11037;
wire n_2181;
wire n_14568;
wire n_11702;
wire n_6069;
wire n_13699;
wire n_171;
wire n_2911;
wire n_14319;
wire n_7497;
wire n_169;
wire n_4655;
wire n_11372;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_7665;
wire n_9354;
wire n_3429;
wire n_10501;
wire n_10817;
wire n_11829;
wire n_14026;
wire n_15324;
wire n_2379;
wire n_11517;
wire n_326;
wire n_7793;
wire n_587;
wire n_8355;
wire n_3554;
wire n_1593;
wire n_6991;
wire n_10556;
wire n_15287;
wire n_1202;
wire n_12741;
wire n_7671;
wire n_7101;
wire n_9436;
wire n_1635;
wire n_7530;
wire n_13150;
wire n_8489;
wire n_15006;
wire n_13776;
wire n_5431;
wire n_15103;
wire n_15619;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_11551;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_14818;
wire n_3462;
wire n_13343;
wire n_7654;
wire n_2851;
wire n_13152;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_9022;
wire n_9238;
wire n_8369;
wire n_358;
wire n_13809;
wire n_160;
wire n_8059;
wire n_10230;
wire n_6633;
wire n_12675;
wire n_2420;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_6579;
wire n_11665;
wire n_13590;
wire n_13907;
wire n_3722;
wire n_186;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_2984;
wire n_11138;
wire n_575;
wire n_11731;
wire n_5187;
wire n_5875;
wire n_9839;
wire n_12821;
wire n_14782;
wire n_4024;
wire n_8831;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_15704;
wire n_732;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_10807;
wire n_12837;
wire n_2240;
wire n_392;
wire n_12478;
wire n_7120;
wire n_12233;
wire n_2538;
wire n_724;
wire n_3250;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_8853;
wire n_1042;
wire n_14070;
wire n_4582;
wire n_14330;
wire n_15327;
wire n_13491;
wire n_1728;
wire n_6252;
wire n_13545;
wire n_557;
wire n_13471;
wire n_1871;
wire n_13760;
wire n_13883;
wire n_4860;
wire n_6211;
wire n_15716;
wire n_845;
wire n_10511;
wire n_140;
wire n_5844;
wire n_8862;
wire n_15748;
wire n_3414;
wire n_10580;
wire n_1549;
wire n_14235;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_768;
wire n_8081;
wire n_7576;
wire n_9675;
wire n_14851;
wire n_6173;
wire n_7786;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_10058;
wire n_2102;
wire n_2563;
wire n_10873;
wire n_14484;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_11454;
wire n_3449;
wire n_13442;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_8900;
wire n_597;
wire n_12523;
wire n_280;
wire n_14444;
wire n_6630;
wire n_6934;
wire n_10484;
wire n_1187;
wire n_9017;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_6737;
wire n_11744;
wire n_4488;
wire n_15726;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_14307;
wire n_8478;
wire n_13450;
wire n_6606;
wire n_2544;
wire n_6695;
wire n_3550;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_15302;
wire n_4211;
wire n_7779;
wire n_10388;
wire n_8999;
wire n_14178;
wire n_6189;
wire n_1206;
wire n_11626;
wire n_12148;
wire n_4016;
wire n_11072;
wire n_15299;
wire n_5867;
wire n_621;
wire n_750;
wire n_5508;
wire n_4656;
wire n_10791;
wire n_6479;
wire n_10506;
wire n_12907;
wire n_15500;
wire n_3839;
wire n_8497;
wire n_2823;
wire n_10770;
wire n_8820;
wire n_6410;
wire n_14891;
wire n_11917;
wire n_9318;
wire n_6158;
wire n_5597;
wire n_9028;
wire n_13944;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_15592;
wire n_8020;
wire n_6090;
wire n_6413;
wire n_1057;
wire n_9374;
wire n_7419;
wire n_15319;
wire n_6506;
wire n_2785;
wire n_235;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_13634;
wire n_12132;
wire n_710;
wire n_1818;
wire n_3730;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_1298;
wire n_10593;
wire n_13019;
wire n_14452;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_13464;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_12182;
wire n_1611;
wire n_12670;
wire n_5050;
wire n_10636;
wire n_12043;
wire n_2740;
wire n_746;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_10203;
wire n_3498;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_15369;
wire n_2401;
wire n_8992;
wire n_15134;
wire n_1589;
wire n_12708;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_9983;
wire n_1497;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_3672;
wire n_7182;
wire n_15453;
wire n_5318;
wire n_13573;
wire n_7365;
wire n_6608;
wire n_10467;
wire n_3533;
wire n_9849;
wire n_1622;
wire n_9109;
wire n_13622;
wire n_6105;
wire n_4725;
wire n_11207;
wire n_6022;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_12493;
wire n_3138;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_14794;
wire n_9237;
wire n_13931;
wire n_11668;
wire n_7885;
wire n_15208;
wire n_15684;
wire n_6860;
wire n_6557;
wire n_14404;
wire n_8466;
wire n_6753;
wire n_12137;
wire n_2171;
wire n_6527;
wire n_7341;
wire n_11328;
wire n_2988;
wire n_9349;
wire n_12306;
wire n_15275;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_11200;
wire n_12088;
wire n_14442;
wire n_15210;
wire n_15423;
wire n_11091;
wire n_8094;
wire n_4109;
wire n_4192;
wire n_10940;
wire n_14377;
wire n_12508;
wire n_4824;
wire n_2808;
wire n_2037;
wire n_4567;
wire n_12096;
wire n_6430;
wire n_6639;
wire n_5150;
wire n_782;
wire n_13418;
wire n_809;
wire n_8832;
wire n_10987;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_1797;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_12891;
wire n_402;
wire n_1870;
wire n_11098;
wire n_11615;
wire n_10533;
wire n_1171;
wire n_11059;
wire n_460;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_1827;
wire n_14616;
wire n_11965;
wire n_4904;
wire n_10938;
wire n_2187;
wire n_10176;
wire n_7517;
wire n_1152;
wire n_6627;
wire n_8080;
wire n_14696;
wire n_450;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_711;
wire n_7745;
wire n_12941;
wire n_3105;
wire n_13551;
wire n_14006;
wire n_2872;
wire n_6666;
wire n_3692;
wire n_10927;
wire n_14258;
wire n_12200;
wire n_4616;
wire n_8321;
wire n_14024;
wire n_9954;
wire n_8735;
wire n_8772;
wire n_4982;
wire n_370;
wire n_1695;
wire n_11722;
wire n_2046;
wire n_2272;
wire n_8786;
wire n_8592;
wire n_15597;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_13682;
wire n_6249;
wire n_2738;
wire n_972;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_1332;
wire n_10155;
wire n_5480;
wire n_9805;
wire n_4323;
wire n_624;
wire n_13593;
wire n_8157;
wire n_2346;
wire n_4831;
wire n_7095;
wire n_936;
wire n_3821;
wire n_3045;
wire n_11461;
wire n_13902;
wire n_10714;
wire n_11701;
wire n_6969;
wire n_885;
wire n_7459;
wire n_6161;
wire n_6615;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_7294;
wire n_3676;
wire n_4896;
wire n_8206;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_11811;
wire n_9110;
wire n_10569;
wire n_2541;
wire n_13745;
wire n_8622;
wire n_2940;
wire n_5904;
wire n_13917;
wire n_4739;
wire n_15367;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_599;
wire n_9335;
wire n_13546;
wire n_14595;
wire n_14468;
wire n_7908;
wire n_12550;
wire n_6062;
wire n_1974;
wire n_4122;
wire n_9452;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_13350;
wire n_13861;
wire n_10051;
wire n_934;
wire n_4209;
wire n_8104;
wire n_10414;
wire n_11255;
wire n_8344;
wire n_2768;
wire n_13592;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_11720;
wire n_4298;
wire n_12673;
wire n_14694;
wire n_2314;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_13874;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_4128;
wire n_10746;
wire n_12225;
wire n_9188;
wire n_6294;
wire n_543;
wire n_5147;
wire n_9611;
wire n_15506;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_1355;
wire n_8779;
wire n_9810;
wire n_14469;
wire n_2258;
wire n_8621;
wire n_5503;
wire n_325;
wire n_5845;
wire n_9250;
wire n_5945;
wire n_804;
wire n_9550;
wire n_11212;
wire n_12884;
wire n_13145;
wire n_10697;
wire n_11714;
wire n_11263;
wire n_10641;
wire n_2390;
wire n_6246;
wire n_8868;
wire n_959;
wire n_2562;
wire n_15070;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_12207;
wire n_1343;
wire n_1522;
wire n_9975;
wire n_2734;
wire n_7250;
wire n_1782;
wire n_5755;
wire n_5600;
wire n_8762;
wire n_12011;
wire n_13195;
wire n_8043;
wire n_8694;
wire n_14492;
wire n_707;
wire n_13965;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_11994;
wire n_7252;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_13419;
wire n_9207;
wire n_13358;
wire n_14134;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_11860;
wire n_11990;
wire n_8728;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_10926;
wire n_14519;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_10626;
wire n_15457;
wire n_6901;
wire n_14345;
wire n_4935;
wire n_13273;
wire n_4694;
wire n_11503;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_2962;
wire n_8171;
wire n_8376;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_1672;
wire n_6774;
wire n_12854;
wire n_15640;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_14816;
wire n_8710;
wire n_737;
wire n_15683;
wire n_12806;
wire n_4045;
wire n_3517;
wire n_3893;
wire n_4598;
wire n_2945;
wire n_3061;
wire n_3932;
wire n_14302;
wire n_3469;
wire n_8599;
wire n_2960;
wire n_8549;
wire n_13460;
wire n_15451;
wire n_10172;
wire n_8054;
wire n_5993;
wire n_11273;
wire n_13904;
wire n_10400;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_138;
wire n_3258;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_14035;
wire n_14496;
wire n_14467;
wire n_13218;
wire n_9096;
wire n_9081;
wire n_13952;
wire n_11697;
wire n_333;
wire n_14789;
wire n_15784;
wire n_13076;
wire n_15526;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_11762;
wire n_11969;
wire n_9236;
wire n_12950;
wire n_7914;
wire n_8628;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_13028;
wire n_14413;
wire n_15150;
wire n_8857;
wire n_8517;
wire n_459;
wire n_4850;
wire n_14243;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_10433;
wire n_2840;
wire n_6779;
wire n_8010;
wire n_285;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_9116;
wire n_1375;
wire n_14096;
wire n_10774;
wire n_3972;
wire n_12332;
wire n_4153;
wire n_10901;
wire n_11034;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_7216;
wire n_12762;
wire n_11499;
wire n_13574;
wire n_1928;
wire n_15364;
wire n_10825;
wire n_14583;
wire n_3091;
wire n_4317;
wire n_14893;
wire n_8275;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_10761;
wire n_14777;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_14057;
wire n_5459;
wire n_9035;
wire n_11579;
wire n_1019;
wire n_10398;
wire n_15303;
wire n_8291;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_11535;
wire n_3642;
wire n_15661;
wire n_12558;
wire n_2845;
wire n_14915;
wire n_4650;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_438;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_1860;
wire n_5016;
wire n_15654;
wire n_1904;
wire n_12975;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_11402;
wire n_479;
wire n_6458;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_9678;
wire n_11401;
wire n_7642;
wire n_8247;
wire n_6577;
wire n_12506;
wire n_13850;
wire n_6740;
wire n_3308;
wire n_12718;
wire n_1113;
wire n_1600;
wire n_12956;
wire n_2253;
wire n_11510;
wire n_12638;
wire n_2366;
wire n_10581;
wire n_14116;
wire n_14856;
wire n_14949;
wire n_15235;
wire n_4912;
wire n_6315;
wire n_4799;
wire n_2261;
wire n_9284;
wire n_12736;
wire n_5086;
wire n_4423;
wire n_5283;
wire n_9111;
wire n_2210;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_3602;
wire n_187;
wire n_3300;
wire n_2978;
wire n_15461;
wire n_12086;
wire n_2516;
wire n_15711;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_6910;
wire n_6262;
wire n_7604;
wire n_14800;
wire n_2827;
wire n_1177;
wire n_7703;
wire n_3515;
wire n_1150;
wire n_9606;
wire n_6319;
wire n_13459;
wire n_566;
wire n_1023;
wire n_2951;
wire n_10470;
wire n_1118;
wire n_14268;
wire n_11589;
wire n_194;
wire n_2949;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_14888;
wire n_1807;
wire n_15034;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_5028;
wire n_5839;
wire n_14240;
wire n_14504;
wire n_1814;
wire n_1631;
wire n_13449;
wire n_14127;
wire n_1879;
wire n_6536;
wire n_12747;
wire n_256;
wire n_440;
wire n_6175;
wire n_3806;
wire n_8827;
wire n_10625;
wire n_7040;
wire n_8280;
wire n_12561;
wire n_12390;
wire n_14460;
wire n_5514;
wire n_13216;
wire n_2931;
wire n_209;
wire n_367;
wire n_8388;
wire n_12849;
wire n_14730;
wire n_2569;
wire n_10235;
wire n_11312;
wire n_3866;
wire n_6978;
wire n_13786;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_671;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_4543;
wire n_10445;
wire n_15110;
wire n_740;
wire n_10738;
wire n_703;
wire n_7378;
wire n_14894;
wire n_12866;
wire n_4157;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_15491;
wire n_15025;
wire n_9190;
wire n_14925;
wire n_6947;
wire n_11612;
wire n_4229;
wire n_9482;
wire n_14918;
wire n_5293;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_12900;
wire n_13414;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_8569;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_14598;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_8877;
wire n_15489;
wire n_9412;
wire n_1401;
wire n_7498;
wire n_10679;
wire n_1516;
wire n_11323;
wire n_10799;
wire n_3846;
wire n_15561;
wire n_6321;
wire n_12914;
wire n_11916;
wire n_180;
wire n_3512;
wire n_7501;
wire n_5201;
wire n_2029;
wire n_10136;
wire n_9506;
wire n_6819;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_1394;
wire n_10585;
wire n_12764;
wire n_13696;
wire n_15148;
wire n_15325;
wire n_1326;
wire n_4783;
wire n_11356;
wire n_1379;
wire n_214;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_13322;
wire n_15158;
wire n_14238;
wire n_9092;
wire n_10034;
wire n_935;
wire n_11148;
wire n_4910;
wire n_9451;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_13934;
wire n_1130;
wire n_3083;
wire n_6899;
wire n_15389;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_676;
wire n_14826;
wire n_15331;
wire n_15776;
wire n_832;
wire n_6592;
wire n_11280;
wire n_12337;
wire n_13254;
wire n_3049;
wire n_14987;
wire n_13466;
wire n_15082;
wire n_15191;
wire n_8686;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_15676;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_14042;
wire n_7613;
wire n_3541;
wire n_11493;
wire n_6101;
wire n_9220;
wire n_14440;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_10528;
wire n_10860;
wire n_12763;
wire n_4930;
wire n_372;
wire n_8588;
wire n_314;
wire n_15229;
wire n_378;
wire n_11339;
wire n_5623;
wire n_15209;
wire n_15269;
wire n_12273;
wire n_13875;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_338;
wire n_15310;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_12712;
wire n_14076;
wire n_506;
wire n_11220;
wire n_360;
wire n_2149;
wire n_9012;
wire n_2396;
wire n_15078;
wire n_4557;
wire n_13012;
wire n_4917;
wire n_8698;
wire n_895;
wire n_8924;
wire n_12584;
wire n_14435;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_14638;
wire n_14946;
wire n_10376;
wire n_15510;
wire n_12752;
wire n_15674;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_15511;
wire n_4593;
wire n_7238;
wire n_344;
wire n_9994;
wire n_2769;
wire n_4465;
wire n_14226;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_14936;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_11596;
wire n_1392;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_14278;
wire n_11885;
wire n_5117;
wire n_1924;
wire n_15618;
wire n_5663;
wire n_525;
wire n_2463;
wire n_3363;
wire n_10224;
wire n_11955;
wire n_12777;
wire n_7572;
wire n_8214;
wire n_1677;
wire n_14706;
wire n_5990;
wire n_611;
wire n_7043;
wire n_10777;
wire n_3721;
wire n_11462;
wire n_3062;
wire n_11732;
wire n_2679;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_14159;
wire n_9134;
wire n_9753;
wire n_13306;
wire n_12819;
wire n_14515;
wire n_8514;
wire n_8722;
wire n_11654;
wire n_12268;
wire n_10214;
wire n_8241;
wire n_8589;
wire n_838;
wire n_12077;
wire n_3969;
wire n_12982;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_15321;
wire n_4231;
wire n_6281;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_13133;
wire n_14757;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_10469;
wire n_445;
wire n_11194;
wire n_9229;
wire n_11480;
wire n_15282;
wire n_6311;
wire n_930;
wire n_7590;
wire n_9342;
wire n_12237;
wire n_13271;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_1945;
wire n_5426;
wire n_10175;
wire n_1656;
wire n_5803;
wire n_11481;
wire n_2112;
wire n_13372;
wire n_1464;
wire n_2430;
wire n_653;
wire n_9868;
wire n_11375;
wire n_1414;
wire n_5285;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_2721;
wire n_944;
wire n_4335;
wire n_9311;
wire n_12275;
wire n_2034;
wire n_576;
wire n_6593;
wire n_13742;
wire n_8630;
wire n_270;
wire n_15177;
wire n_2683;
wire n_12376;
wire n_563;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_8145;
wire n_8405;
wire n_10447;
wire n_9260;
wire n_15063;
wire n_7176;
wire n_14534;
wire n_8928;
wire n_13630;
wire n_7682;
wire n_15223;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_626;
wire n_990;
wire n_11925;
wire n_13700;
wire n_12509;
wire n_8948;
wire n_10406;
wire n_6231;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_14902;
wire n_8672;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_11985;
wire n_6746;
wire n_13527;
wire n_498;
wire n_8447;
wire n_7901;
wire n_870;
wire n_5395;
wire n_1253;
wire n_10522;
wire n_366;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_13793;
wire n_11782;
wire n_1693;
wire n_6446;
wire n_10278;
wire n_14290;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_3802;
wire n_348;
wire n_3256;
wire n_6996;
wire n_7218;
wire n_9430;
wire n_8828;
wire n_376;
wire n_15384;
wire n_11407;
wire n_2118;
wire n_2111;
wire n_13882;
wire n_390;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_2915;
wire n_12710;
wire n_15686;
wire n_1148;
wire n_6749;
wire n_2188;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_1989;
wire n_7005;
wire n_10408;
wire n_2802;
wire n_8572;
wire n_10798;
wire n_10965;
wire n_7732;
wire n_13325;
wire n_14850;
wire n_15135;
wire n_3643;
wire n_6181;
wire n_6337;
wire n_7447;
wire n_2425;
wire n_9776;
wire n_11911;
wire n_6777;
wire n_4265;
wire n_11987;
wire n_11442;
wire n_12936;
wire n_8227;
wire n_12721;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_8475;
wire n_3060;
wire n_11730;
wire n_10482;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_4105;
wire n_1851;
wire n_14064;
wire n_14524;
wire n_1090;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_12039;
wire n_4926;
wire n_1518;
wire n_11651;
wire n_1362;
wire n_11388;
wire n_14151;
wire n_3123;
wire n_9386;
wire n_3380;
wire n_8314;
wire n_10154;
wire n_5617;
wire n_1829;
wire n_15120;
wire n_7922;
wire n_13089;
wire n_15459;
wire n_15192;
wire n_10377;
wire n_5580;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_10033;
wire n_9926;
wire n_3038;
wire n_570;
wire n_11121;
wire n_13167;
wire n_11270;
wire n_1789;
wire n_12329;
wire n_6310;
wire n_15161;
wire n_11689;
wire n_620;
wire n_10003;
wire n_15601;
wire n_519;
wire n_8311;
wire n_2523;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_12253;
wire n_1482;
wire n_11147;
wire n_12928;
wire n_15005;
wire n_5310;
wire n_9661;
wire n_9843;
wire n_15013;
wire n_9877;
wire n_8764;
wire n_14284;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_14945;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_13001;
wire n_5390;
wire n_13232;
wire n_9901;
wire n_1710;
wire n_2161;
wire n_13320;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_12990;
wire n_14246;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_2047;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_11817;
wire n_13278;
wire n_8567;
wire n_15455;
wire n_1609;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_13597;
wire n_14957;
wire n_5133;
wire n_409;
wire n_13488;
wire n_11042;
wire n_1763;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_13447;
wire n_3989;
wire n_7089;
wire n_2490;
wire n_7144;
wire n_7286;
wire n_11479;
wire n_11737;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_14681;
wire n_635;
wire n_12028;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_13016;
wire n_11272;
wire n_13668;
wire n_13095;
wire n_14230;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_1996;
wire n_14708;
wire n_6332;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_12048;
wire n_5853;
wire n_15032;
wire n_8283;
wire n_5982;
wire n_1158;
wire n_10930;
wire n_2248;
wire n_11600;
wire n_15085;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_14546;
wire n_7129;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_13938;
wire n_12057;
wire n_6696;
wire n_15440;
wire n_753;
wire n_3925;
wire n_13251;
wire n_9882;
wire n_9527;
wire n_3180;
wire n_8566;
wire n_7343;
wire n_2795;
wire n_12766;
wire n_14875;
wire n_3472;
wire n_8516;
wire n_10637;
wire n_8302;
wire n_15056;
wire n_8317;
wire n_5376;
wire n_15610;
wire n_12229;
wire n_14003;
wire n_5106;
wire n_269;
wire n_6116;
wire n_9205;
wire n_359;
wire n_9511;
wire n_8167;
wire n_15329;
wire n_7859;
wire n_14315;
wire n_6730;
wire n_7872;
wire n_7492;
wire n_13670;
wire n_7972;
wire n_11254;
wire n_13319;
wire n_15023;
wire n_1479;
wire n_4768;
wire n_11617;
wire n_1675;
wire n_13858;
wire n_13512;
wire n_9071;
wire n_7916;
wire n_3717;
wire n_9368;
wire n_10415;
wire n_7694;
wire n_5561;
wire n_13069;
wire n_7480;
wire n_11711;
wire n_5410;
wire n_571;
wire n_2215;
wire n_12362;
wire n_404;
wire n_8944;
wire n_6167;
wire n_15666;
wire n_158;
wire n_1884;
wire n_13233;
wire n_11931;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_665;
wire n_8109;
wire n_13297;
wire n_9459;
wire n_14185;
wire n_2055;
wire n_5156;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_2553;
wire n_6307;
wire n_149;
wire n_10410;
wire n_632;
wire n_6094;
wire n_9098;
wire n_2038;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_14953;
wire n_9133;
wire n_12664;
wire n_14942;
wire n_14873;
wire n_15604;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_373;
wire n_9504;
wire n_15359;
wire n_14840;
wire n_8975;
wire n_6267;
wire n_9063;
wire n_7787;
wire n_1833;
wire n_3903;
wire n_12360;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_9268;
wire n_1850;
wire n_15431;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_15035;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_1417;
wire n_10456;
wire n_15631;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_14083;
wire n_13186;
wire n_5916;
wire n_681;
wire n_11907;
wire n_15655;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_3094;
wire n_10025;
wire n_412;
wire n_10627;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_14755;
wire n_6299;
wire n_6813;
wire n_965;
wire n_8825;
wire n_1428;
wire n_12969;
wire n_1576;
wire n_15430;
wire n_1856;
wire n_11753;
wire n_2077;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_15732;
wire n_8266;
wire n_5691;
wire n_1059;
wire n_12457;
wire n_4951;
wire n_8981;
wire n_422;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_3079;
wire n_165;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_13519;
wire n_15750;
wire n_540;
wire n_14170;
wire n_4039;
wire n_457;
wire n_3800;
wire n_3070;
wire n_13496;
wire n_15641;
wire n_4566;
wire n_3263;
wire n_12939;
wire n_6316;
wire n_15038;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_1748;
wire n_13884;
wire n_10404;
wire n_8639;
wire n_8138;
wire n_8058;
wire n_9308;
wire n_3504;
wire n_6638;
wire n_12779;
wire n_11838;
wire n_10508;
wire n_531;
wire n_7719;
wire n_4272;
wire n_10811;
wire n_14049;
wire n_8333;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_7562;
wire n_6220;
wire n_3111;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_336;
wire n_6985;
wire n_7619;
wire n_12783;
wire n_7170;
wire n_13853;
wire n_9211;
wire n_12019;
wire n_1885;
wire n_8176;
wire n_8124;
wire n_14529;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_10891;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_3054;
wire n_10803;
wire n_15284;
wire n_1538;
wire n_8147;
wire n_1240;
wire n_13190;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_1234;
wire n_14014;
wire n_14195;
wire n_5262;
wire n_10700;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_11695;
wire n_4620;
wire n_3152;
wire n_8458;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_7935;
wire n_14247;
wire n_6772;
wire n_8113;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_11453;
wire n_4127;
wire n_14300;
wire n_15443;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_168;
wire n_6318;
wire n_15418;
wire n_2353;
wire n_11970;
wire n_4099;
wire n_14678;
wire n_7918;
wire n_13599;
wire n_4517;
wire n_4168;
wire n_14690;
wire n_15008;
wire n_5188;
wire n_13647;
wire n_6916;
wire n_1738;
wire n_15524;
wire n_4490;
wire n_13683;
wire n_1575;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_1923;
wire n_10783;
wire n_2260;
wire n_10147;
wire n_12163;
wire n_11862;
wire n_14839;
wire n_10725;
wire n_3952;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_12944;
wire n_3911;
wire n_8290;
wire n_15409;
wire n_7536;
wire n_7472;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_11660;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_10812;
wire n_14709;
wire n_1743;
wire n_12297;
wire n_13848;
wire n_14249;
wire n_6366;
wire n_6230;
wire n_14241;
wire n_2997;
wire n_6604;
wire n_1991;
wire n_14497;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_10001;
wire n_3708;
wire n_11107;
wire n_14280;
wire n_4078;
wire n_13724;
wire n_13280;
wire n_9301;
wire n_12145;
wire n_3046;
wire n_11088;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_10284;
wire n_12757;
wire n_8160;
wire n_12054;
wire n_14379;
wire n_5659;
wire n_8099;
wire n_14446;
wire n_11595;
wire n_8840;
wire n_3619;
wire n_11405;
wire n_14719;
wire n_15575;
wire n_13768;
wire n_1415;
wire n_13189;
wire n_5881;
wire n_8522;
wire n_12971;
wire n_1370;
wire n_7222;
wire n_1786;
wire n_7942;
wire n_6473;
wire n_13103;
wire n_13838;
wire n_8578;
wire n_15630;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_10046;
wire n_12328;
wire n_14558;
wire n_15696;
wire n_2291;
wire n_415;
wire n_11318;
wire n_9083;
wire n_1371;
wire n_7725;
wire n_383;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_10977;
wire n_200;
wire n_11299;
wire n_2184;
wire n_10397;
wire n_2982;
wire n_6483;
wire n_1803;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_4065;
wire n_14004;
wire n_5863;
wire n_229;
wire n_7647;
wire n_10936;
wire n_8626;
wire n_2645;
wire n_12442;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_2630;
wire n_15123;
wire n_1444;
wire n_9835;
wire n_15068;
wire n_15442;
wire n_1603;
wire n_7300;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_2470;
wire n_4446;
wire n_14666;
wire n_1263;
wire n_13605;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_13995;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_4733;
wire n_13441;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_14237;
wire n_1261;
wire n_15095;
wire n_3879;
wire n_11240;
wire n_2286;
wire n_4743;
wire n_10207;
wire n_13857;
wire n_13841;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_13556;
wire n_1143;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_13367;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_658;
wire n_1874;
wire n_13816;
wire n_11487;
wire n_2865;
wire n_2825;
wire n_8441;
wire n_11441;
wire n_2013;
wire n_14203;
wire n_6076;
wire n_8933;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_7778;
wire n_15231;
wire n_758;
wire n_12844;
wire n_5851;
wire n_14736;
wire n_11287;
wire n_2256;
wire n_9755;
wire n_7073;
wire n_943;
wire n_4060;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_4879;
wire n_10139;
wire n_13246;
wire n_13409;
wire n_14061;
wire n_6390;
wire n_5796;
wire n_10104;
wire n_772;
wire n_8726;
wire n_12986;
wire n_11381;
wire n_2806;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_770;
wire n_15789;
wire n_9117;
wire n_9720;
wire n_3028;
wire n_9381;
wire n_3662;
wire n_10169;
wire n_2981;
wire n_6958;
wire n_3076;
wire n_7746;
wire n_15727;
wire n_12049;
wire n_12690;
wire n_14498;
wire n_15417;
wire n_886;
wire n_7563;
wire n_343;
wire n_12475;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_539;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_14667;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_14713;
wire n_15512;
wire n_4117;
wire n_7853;
wire n_12526;
wire n_4687;
wire n_14414;
wire n_15565;
wire n_2836;
wire n_7531;
wire n_12377;
wire n_638;
wire n_1404;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_13214;
wire n_8615;
wire n_11062;
wire n_13650;
wire n_2378;
wire n_7721;
wire n_887;
wire n_7192;
wire n_14202;
wire n_15636;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_14554;
wire n_9887;
wire n_9149;
wire n_2655;
wire n_4600;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_13211;
wire n_1467;
wire n_8316;
wire n_4250;
wire n_9990;
wire n_5829;
wire n_3906;
wire n_10005;
wire n_224;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_14874;
wire n_2599;
wire n_15311;
wire n_8505;
wire n_15113;
wire n_9273;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_15498;
wire n_2370;
wire n_2612;
wire n_8970;
wire n_7527;
wire n_13061;
wire n_7417;
wire n_9682;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_12513;
wire n_2214;
wire n_4253;
wire n_10640;
wire n_407;
wire n_913;
wire n_6582;
wire n_5734;
wire n_15098;
wire n_2593;
wire n_13395;
wire n_4255;
wire n_867;
wire n_4071;
wire n_10729;
wire n_12545;
wire n_14656;
wire n_7388;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_11657;
wire n_9924;
wire n_14745;
wire n_8717;
wire n_14744;
wire n_13336;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_13176;
wire n_4605;
wire n_15091;
wire n_9064;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_13102;
wire n_163;
wire n_1644;
wire n_11268;
wire n_12753;
wire n_14760;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_14135;
wire n_9254;
wire n_1558;
wire n_12894;
wire n_7090;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_4305;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_13375;
wire n_13390;
wire n_13691;
wire n_824;
wire n_15769;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_4297;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_13264;
wire n_8378;
wire n_2907;
wire n_577;
wire n_8687;
wire n_5374;
wire n_14194;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_12010;
wire n_1843;
wire n_619;
wire n_5675;
wire n_9738;
wire n_12026;
wire n_9570;
wire n_4227;
wire n_521;
wire n_2778;
wire n_12356;
wire n_11857;
wire n_13825;
wire n_395;
wire n_1909;
wire n_6240;
wire n_11077;
wire n_8243;
wire n_8633;
wire n_6347;
wire n_5020;
wire n_9593;
wire n_9846;
wire n_13262;
wire n_13482;
wire n_7689;
wire n_6511;
wire n_606;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_1123;
wire n_1309;
wire n_9469;
wire n_10764;
wire n_13398;
wire n_9677;
wire n_2961;
wire n_15598;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_483;
wire n_6804;
wire n_1970;
wire n_14676;
wire n_8449;
wire n_6358;
wire n_630;
wire n_2059;
wire n_13204;
wire n_2669;
wire n_4094;
wire n_14331;
wire n_6603;
wire n_4765;
wire n_2546;
wire n_13873;
wire n_3193;
wire n_2522;
wire n_476;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_1957;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_8801;
wire n_4732;
wire n_3912;
wire n_6986;
wire n_10438;
wire n_3118;
wire n_9322;
wire n_15017;
wire n_11201;
wire n_5959;
wire n_3720;
wire n_10531;
wire n_1907;
wire n_14964;
wire n_2529;
wire n_8031;
wire n_8918;
wire n_264;
wire n_12878;
wire n_15591;
wire n_9348;
wire n_14262;
wire n_12188;
wire n_860;
wire n_8219;
wire n_1530;
wire n_15373;
wire n_8696;
wire n_4745;
wire n_938;
wire n_1302;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_15167;
wire n_12630;
wire n_4581;
wire n_6890;
wire n_549;
wire n_11028;
wire n_12171;
wire n_4377;
wire n_12299;
wire n_15706;
wire n_12022;
wire n_9249;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_2143;
wire n_8180;
wire n_905;
wire n_10741;
wire n_15211;
wire n_6109;
wire n_14727;
wire n_10760;
wire n_4792;
wire n_15580;
wire n_12425;
wire n_14762;
wire n_9444;
wire n_15334;
wire n_7731;
wire n_1680;
wire n_3842;
wire n_10772;
wire n_322;
wire n_993;
wire n_11527;
wire n_689;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_1605;
wire n_13507;
wire n_3514;
wire n_11327;
wire n_10915;
wire n_4979;
wire n_1988;
wire n_9535;
wire n_558;
wire n_6770;
wire n_2654;
wire n_3036;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_5302;
wire n_12000;
wire n_966;
wire n_15410;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_12490;
wire n_15151;
wire n_3357;
wire n_13594;
wire n_692;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_14182;
wire n_3895;
wire n_487;
wire n_8943;
wire n_8486;
wire n_241;
wire n_14767;
wire n_10279;
wire n_4520;
wire n_5299;
wire n_12829;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_14352;
wire n_13889;
wire n_14773;
wire n_10680;
wire n_2459;
wire n_10127;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_13654;
wire n_5361;
wire n_11610;
wire n_7132;
wire n_2711;
wire n_11814;
wire n_12255;
wire n_12739;
wire n_7081;
wire n_13015;
wire n_4199;
wire n_6663;
wire n_5885;
wire n_14228;
wire n_1912;
wire n_9723;
wire n_5356;
wire n_12609;
wire n_4441;
wire n_7319;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_1312;
wire n_11176;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_11360;
wire n_8155;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5038;
wire n_268;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_10039;
wire n_11726;
wire n_10854;
wire n_11358;
wire n_5463;
wire n_3022;
wire n_13366;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_247;
wire n_12904;
wire n_8833;
wire n_9191;
wire n_10142;
wire n_1165;
wire n_5892;
wire n_7828;
wire n_14623;
wire n_4773;
wire n_5489;
wire n_7940;
wire n_9918;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_9034;
wire n_328;
wire n_1386;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_9390;
wire n_5113;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_8074;
wire n_15381;
wire n_8485;
wire n_13639;
wire n_14852;
wire n_8860;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_6621;
wire n_11958;
wire n_15624;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_1214;
wire n_13070;
wire n_690;
wire n_850;
wire n_8271;
wire n_15514;
wire n_5692;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_4800;
wire n_9266;
wire n_1157;
wire n_3453;
wire n_14491;
wire n_12728;
wire n_5555;
wire n_3410;
wire n_15011;
wire n_10027;
wire n_12784;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_825;
wire n_13678;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_14582;
wire n_8699;
wire n_3785;
wire n_14261;
wire n_14677;
wire n_6897;
wire n_13523;
wire n_2963;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_5366;
wire n_14928;
wire n_2602;
wire n_15550;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_9078;
wire n_8225;
wire n_9536;
wire n_2980;
wire n_13778;
wire n_696;
wire n_14250;
wire n_4886;
wire n_9931;
wire n_13198;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_13741;
wire n_13819;
wire n_4055;
wire n_15777;
wire n_12610;
wire n_14634;
wire n_2178;
wire n_11671;
wire n_10328;
wire n_14416;
wire n_5968;
wire n_11251;
wire n_14424;
wire n_14523;
wire n_12293;
wire n_11063;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_10753;
wire n_6497;
wire n_9989;
wire n_8319;
wire n_13174;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_7108;
wire n_14455;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_1796;
wire n_8368;
wire n_15691;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_11879;
wire n_2082;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_15376;
wire n_8546;
wire n_10963;
wire n_8300;
wire n_15336;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_15050;
wire n_678;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_14161;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_283;
wire n_8148;
wire n_11400;
wire n_13290;
wire n_8150;
wire n_13500;
wire n_3578;
wire n_909;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_15398;
wire n_10483;
wire n_15593;
wire n_12160;
wire n_4737;
wire n_590;
wire n_11563;
wire n_4925;
wire n_9620;
wire n_4116;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_362;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_5419;
wire n_11243;
wire n_1990;
wire n_3805;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_14513;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_11939;
wire n_6409;
wire n_1634;
wire n_3252;
wire n_627;
wire n_3253;
wire n_7954;
wire n_9824;
wire n_1465;
wire n_11119;
wire n_342;
wire n_14347;
wire n_2622;
wire n_15089;
wire n_7951;
wire n_2658;
wire n_7552;
wire n_8096;
wire n_2665;
wire n_11468;
wire n_14602;
wire n_13901;
wire n_12166;
wire n_2133;
wire n_1712;
wire n_8233;
wire n_4603;
wire n_6130;
wire n_7273;
wire n_9683;
wire n_1523;
wire n_10646;
wire n_14750;
wire n_7231;
wire n_15725;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_11704;
wire n_3128;
wire n_14074;
wire n_15252;
wire n_15132;
wire n_1527;
wire n_495;
wire n_5732;
wire n_5372;
wire n_14050;
wire n_11878;
wire n_15763;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_15749;
wire n_15317;
wire n_7449;
wire n_12800;
wire n_2230;
wire n_8763;
wire n_7772;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_14197;
wire n_8679;
wire n_15638;
wire n_1565;
wire n_7239;
wire n_14289;
wire n_1493;
wire n_15582;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_15145;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_2573;
wire n_2646;
wire n_15297;
wire n_2535;
wire n_9561;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_13979;
wire n_6623;
wire n_12070;
wire n_9714;
wire n_1364;
wire n_9740;
wire n_3078;
wire n_9773;
wire n_13316;
wire n_2436;
wire n_10313;
wire n_14898;
wire n_15672;
wire n_615;
wire n_3838;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_13689;
wire n_3941;
wire n_15413;
wire n_3793;
wire n_10216;
wire n_15628;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_15160;
wire n_3789;
wire n_605;
wire n_1514;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_12354;
wire n_12666;
wire n_14297;
wire n_14395;
wire n_13528;
wire n_12581;
wire n_6047;
wire n_8292;
wire n_12631;
wire n_3037;
wire n_1646;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_3729;
wire n_10773;
wire n_8601;
wire n_4994;
wire n_6652;
wire n_9377;
wire n_2537;
wire n_11932;
wire n_10971;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_6970;
wire n_6921;
wire n_5168;
wire n_14836;
wire n_4661;
wire n_1308;
wire n_13027;
wire n_12867;
wire n_4988;
wire n_7674;
wire n_14675;
wire n_9826;
wire n_3171;
wire n_12607;
wire n_14516;
wire n_7568;
wire n_15343;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_15782;
wire n_12075;
wire n_4540;
wire n_11942;
wire n_6344;
wire n_2097;
wire n_12305;
wire n_13489;
wire n_12123;
wire n_3459;
wire n_9772;
wire n_12170;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_15370;
wire n_9630;
wire n_3499;
wire n_7724;
wire n_6624;
wire n_6956;
wire n_4284;
wire n_13313;
wire n_13927;
wire n_12966;
wire n_13877;
wire n_15308;
wire n_6305;
wire n_9255;
wire n_1005;
wire n_1947;
wire n_6209;
wire n_10231;
wire n_12547;
wire n_8310;
wire n_9758;
wire n_15577;
wire n_3426;
wire n_11922;
wire n_4971;
wire n_14020;
wire n_15175;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_12358;
wire n_14502;
wire n_7329;
wire n_15206;
wire n_8646;
wire n_7408;
wire n_13415;
wire n_9691;
wire n_12997;
wire n_14533;
wire n_10259;
wire n_14005;
wire n_2650;
wire n_7107;
wire n_14293;
wire n_5652;
wire n_6457;
wire n_10488;
wire n_8597;
wire n_14334;
wire n_987;
wire n_7690;
wire n_8969;
wire n_14187;
wire n_15245;
wire n_7123;
wire n_10752;
wire n_11577;
wire n_15225;
wire n_5499;
wire n_720;
wire n_8117;
wire n_10067;
wire n_153;
wire n_15169;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_13562;
wire n_14537;
wire n_12498;
wire n_13888;
wire n_656;
wire n_11475;
wire n_6950;
wire n_8208;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_797;
wire n_11010;
wire n_2933;
wire n_10274;
wire n_15614;
wire n_9590;
wire n_2717;
wire n_1723;
wire n_11588;
wire n_1878;
wire n_189;
wire n_738;
wire n_2012;
wire n_6694;
wire n_3497;
wire n_13956;
wire n_15318;
wire n_9168;
wire n_5066;
wire n_6880;
wire n_7418;
wire n_2842;
wire n_3580;
wire n_14220;
wire n_11221;
wire n_13837;
wire n_12387;
wire n_2335;
wire n_9497;
wire n_15772;
wire n_8536;
wire n_13255;
wire n_9435;
wire n_7229;
wire n_14245;
wire n_8350;
wire n_529;
wire n_2307;
wire n_3704;
wire n_11448;
wire n_684;
wire n_9219;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_15502;
wire n_8914;
wire n_15076;
wire n_1181;
wire n_12576;
wire n_15559;
wire n_7258;
wire n_15276;
wire n_5190;
wire n_13892;
wire n_8391;
wire n_14221;
wire n_10579;
wire n_10832;
wire n_13345;
wire n_3173;
wire n_13964;
wire n_13749;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_1049;
wire n_14559;
wire n_6466;
wire n_7864;
wire n_15552;
wire n_6727;
wire n_4097;
wire n_14360;
wire n_1666;
wire n_10584;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_12862;
wire n_2449;
wire n_11445;
wire n_13151;
wire n_3880;
wire n_13621;
wire n_13601;
wire n_14052;
wire n_14311;
wire n_3685;
wire n_8216;
wire n_11552;
wire n_13765;
wire n_2868;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_15102;
wire n_14733;
wire n_11874;
wire n_13926;
wire n_2231;
wire n_3609;
wire n_9982;
wire n_10171;
wire n_15184;
wire n_14157;
wire n_1228;
wire n_5455;
wire n_417;
wire n_5442;
wire n_6386;
wire n_14317;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_12656;
wire n_9852;
wire n_272;
wire n_6820;
wire n_2896;
wire n_11623;
wire n_8313;
wire n_3019;
wire n_2639;
wire n_14828;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_15779;
wire n_2368;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_458;
wire n_4175;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_10540;
wire n_11936;
wire n_15366;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_3200;
wire n_4771;
wire n_10200;
wire n_13392;
wire n_12734;
wire n_7332;
wire n_3259;
wire n_2524;
wire n_10382;
wire n_13164;
wire n_3167;
wire n_2460;
wire n_7185;
wire n_5836;
wire n_6291;
wire n_11489;
wire n_13662;
wire n_3867;
wire n_10269;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_12262;
wire n_13223;
wire n_1073;
wire n_13340;
wire n_9169;
wire n_252;
wire n_14910;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_13728;
wire n_7512;
wire n_14385;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_11018;
wire n_10981;
wire n_14499;
wire n_8738;
wire n_7766;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_15368;
wire n_12797;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_11376;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_9481;
wire n_13379;
wire n_8798;
wire n_9600;
wire n_13781;
wire n_2877;
wire n_9122;
wire n_14731;
wire n_8085;
wire n_11274;
wire n_5098;
wire n_1021;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_811;
wire n_683;
wire n_1207;
wire n_12012;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_9927;
wire n_14613;
wire n_5497;
wire n_10076;
wire n_11515;
wire n_8721;
wire n_880;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_3505;
wire n_13558;
wire n_3540;
wire n_3577;
wire n_11554;
wire n_15657;
wire n_7637;
wire n_2432;
wire n_10148;
wire n_150;
wire n_1478;
wire n_10318;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_3641;
wire n_4203;
wire n_7127;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_9635;
wire n_13890;
wire n_5481;
wire n_12890;
wire n_3590;
wire n_8666;
wire n_2435;
wire n_15513;
wire n_5344;
wire n_954;
wire n_9264;
wire n_13994;
wire n_14483;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_15724;
wire n_14308;
wire n_1382;
wire n_5408;
wire n_7801;
wire n_1736;
wire n_13484;
wire n_9155;
wire n_4053;
wire n_10234;
wire n_8460;
wire n_1483;
wire n_3848;
wire n_10416;
wire n_1372;
wire n_3327;
wire n_14370;
wire n_14593;
wire n_1719;
wire n_8836;
wire n_7959;
wire n_13430;
wire n_319;
wire n_7019;
wire n_8181;
wire n_2701;
wire n_2511;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_8254;
wire n_13452;
wire n_13521;
wire n_4167;
wire n_8071;
wire n_1427;
wire n_2745;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_1080;
wire n_6667;
wire n_14926;
wire n_7409;
wire n_5271;
wire n_10735;
wire n_10583;
wire n_10731;
wire n_9878;
wire n_562;
wire n_6004;
wire n_13807;
wire n_10806;
wire n_14591;
wire n_5964;
wire n_2323;
wire n_14363;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_11628;
wire n_7444;
wire n_14576;
wire n_162;
wire n_5234;
wire n_4431;
wire n_7546;
wire n_6357;
wire n_2421;
wire n_1136;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_14274;
wire n_6588;
wire n_3265;
wire n_11549;
wire n_2464;
wire n_1125;
wire n_4042;
wire n_3755;
wire n_5128;
wire n_14033;
wire n_12286;
wire n_9001;
wire n_2224;
wire n_10393;
wire n_15403;
wire n_11498;
wire n_13081;
wire n_2329;
wire n_1092;
wire n_15221;
wire n_15602;
wire n_10513;
wire n_12252;
wire n_441;
wire n_5467;
wire n_10439;
wire n_14545;
wire n_8013;
wire n_4299;
wire n_7296;
wire n_12627;
wire n_4890;
wire n_146;
wire n_1784;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_193;
wire n_1775;
wire n_12281;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_2410;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_1093;
wire n_9373;
wire n_15012;
wire n_14337;
wire n_1783;
wire n_6268;
wire n_2929;
wire n_4176;
wire n_12347;
wire n_5199;
wire n_14551;
wire n_5827;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_296;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_9967;
wire n_13553;
wire n_7521;
wire n_651;
wire n_14088;
wire n_3407;
wire n_5992;
wire n_217;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_13817;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_7187;
wire n_9971;
wire n_3425;
wire n_215;
wire n_15517;
wire n_10894;
wire n_3894;
wire n_14118;
wire n_13974;
wire n_9524;
wire n_12277;
wire n_14917;
wire n_3127;
wire n_1831;
wire n_12698;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_9243;
wire n_9182;
wire n_6467;
wire n_9282;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_1453;
wire n_15680;
wire n_10083;
wire n_6336;
wire n_6796;
wire n_2502;
wire n_3646;
wire n_10347;
wire n_9224;
wire n_5513;
wire n_5614;
wire n_497;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_12410;
wire n_4830;
wire n_4706;
wire n_13225;
wire n_14855;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_14707;
wire n_15326;
wire n_1224;
wire n_2783;
wire n_10208;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_14726;
wire n_1470;
wire n_8141;
wire n_14612;
wire n_12294;
wire n_14180;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_14058;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_13355;
wire n_12957;
wire n_2732;
wire n_4693;
wire n_13141;
wire n_4206;
wire n_11616;
wire n_14065;
wire n_8791;
wire n_11920;
wire n_2249;
wire n_8288;
wire n_10793;
wire n_1091;
wire n_2000;
wire n_14672;
wire n_3862;
wire n_14366;
wire n_4267;
wire n_15127;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_2270;
wire n_1425;
wire n_12786;
wire n_5049;
wire n_13382;
wire n_12711;
wire n_11675;
wire n_983;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_15543;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_10440;
wire n_1733;
wire n_8006;
wire n_10391;
wire n_8323;
wire n_7636;
wire n_9799;
wire n_9695;
wire n_8296;
wire n_2955;
wire n_11083;
wire n_5592;
wire n_6954;
wire n_2158;
wire n_6938;
wire n_4609;
wire n_7866;
wire n_1855;
wire n_3051;
wire n_11306;
wire n_7190;
wire n_15143;
wire n_9784;
wire n_11198;
wire n_3367;
wire n_7205;
wire n_385;
wire n_1687;
wire n_8757;
wire n_1439;
wire n_2328;
wire n_7990;
wire n_7020;
wire n_2859;
wire n_10036;
wire n_2202;
wire n_13035;
wire n_13021;
wire n_1331;
wire n_613;
wire n_736;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_14905;
wire n_8596;
wire n_15128;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_11840;
wire n_2993;
wire n_4754;
wire n_3016;
wire n_4647;
wire n_11698;
wire n_1134;
wire n_3688;
wire n_11292;
wire n_9556;
wire n_10261;
wire n_13157;
wire n_8590;
wire n_8720;
wire n_4003;
wire n_5708;
wire n_554;
wire n_1995;
wire n_3751;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_4894;
wire n_5474;
wire n_14084;
wire n_15798;
wire n_12289;
wire n_4113;
wire n_10813;
wire n_1889;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_11326;
wire n_13046;
wire n_6421;
wire n_435;
wire n_1905;
wire n_13935;
wire n_11870;
wire n_7407;
wire n_9827;
wire n_14009;
wire n_3466;
wire n_13334;
wire n_10907;
wire n_762;
wire n_5704;
wire n_15787;
wire n_11431;
wire n_4983;
wire n_1778;
wire n_7148;
wire n_14002;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_13646;
wire n_11834;
wire n_9417;
wire n_6236;
wire n_1079;
wire n_13361;
wire n_2139;
wire n_12020;
wire n_419;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_15061;
wire n_6007;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_3338;
wire n_144;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_2219;
wire n_6835;
wire n_1203;
wire n_8834;
wire n_3636;
wire n_11624;
wire n_13399;
wire n_2327;
wire n_14010;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_15262;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_11234;
wire n_10822;
wire n_14697;
wire n_15030;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_13967;
wire n_12099;
wire n_12858;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_2304;
wire n_14609;
wire n_15351;
wire n_7799;
wire n_8364;
wire n_2487;
wire n_5698;
wire n_11092;
wire n_3276;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_14310;
wire n_15228;
wire n_13380;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_13053;
wire n_9792;
wire n_10720;
wire n_7513;
wire n_9336;
wire n_10535;
wire n_3572;
wire n_11836;
wire n_349;
wire n_6602;
wire n_10924;
wire n_3886;
wire n_15281;
wire n_15792;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_15675;
wire n_9647;
wire n_15515;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_10885;
wire n_15106;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_443;
wire n_892;
wire n_13201;
wire n_3637;
wire n_6242;
wire n_12527;
wire n_4574;
wire n_14759;
wire n_13274;
wire n_12379;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_9312;
wire n_2156;
wire n_9019;
wire n_1718;
wire n_13891;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_4234;
wire n_12477;
wire n_7469;
wire n_5538;
wire n_14325;
wire n_15503;
wire n_14078;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_1768;
wire n_14309;
wire n_10895;
wire n_3974;
wire n_198;
wire n_1847;
wire n_3634;
wire n_10875;
wire n_11736;
wire n_11977;
wire n_7560;
wire n_14729;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_15576;
wire n_1397;
wire n_14222;
wire n_3236;
wire n_11696;
wire n_12400;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_11734;
wire n_1841;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_12114;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_1623;
wire n_11507;
wire n_14430;
wire n_9145;
wire n_15337;
wire n_1015;
wire n_13996;
wire n_7082;
wire n_12092;
wire n_14749;
wire n_3112;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_4270;
wire n_11837;
wire n_5428;
wire n_4151;
wire n_13709;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_3417;
wire n_13898;
wire n_9000;
wire n_5677;
wire n_9454;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_14704;
wire n_785;
wire n_8307;
wire n_5153;
wire n_11967;
wire n_9383;
wire n_9253;
wire n_15084;
wire n_609;
wire n_13559;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_15258;
wire n_5927;
wire n_15071;
wire n_7495;
wire n_7392;
wire n_11996;
wire n_11338;
wire n_9566;
wire n_5435;
wire n_2337;
wire n_13426;
wire n_12174;
wire n_9765;
wire n_1356;
wire n_3213;
wire n_9807;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_8706;
wire n_9057;
wire n_15220;
wire n_6400;
wire n_2607;
wire n_7945;
wire n_7666;
wire n_8894;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_6941;
wire n_12053;
wire n_1943;
wire n_5566;
wire n_11250;
wire n_7829;
wire n_12619;
wire n_3249;
wire n_1320;
wire n_7543;
wire n_13504;
wire n_15328;
wire n_8680;
wire n_11289;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_13169;
wire n_7877;
wire n_7963;
wire n_13555;
wire n_9672;
wire n_2499;
wire n_12582;
wire n_4152;
wire n_5487;
wire n_15291;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_302;
wire n_5486;
wire n_9503;
wire n_15345;
wire n_12423;
wire n_137;
wire n_11391;
wire n_15426;
wire n_15462;
wire n_1596;
wire n_5244;
wire n_5092;
wire n_14721;
wire n_14137;
wire n_1734;
wire n_3172;
wire n_13265;
wire n_12714;
wire n_4832;
wire n_8270;
wire n_2902;
wire n_5889;
wire n_11738;
wire n_3217;
wire n_7284;
wire n_12153;
wire n_1983;
wire n_7264;
wire n_5391;
wire n_11522;
wire n_1938;
wire n_9763;
wire n_14163;
wire n_7737;
wire n_13666;
wire n_15523;
wire n_6537;
wire n_8614;
wire n_2472;
wire n_7328;
wire n_11070;
wire n_10702;
wire n_13337;
wire n_10958;
wire n_15682;
wire n_15112;
wire n_9479;
wire n_3394;
wire n_15556;
wire n_9162;
wire n_9568;
wire n_1715;
wire n_13730;
wire n_14849;
wire n_15621;
wire n_3536;
wire n_12405;
wire n_8816;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_14041;
wire n_3710;
wire n_9119;
wire n_4195;
wire n_10319;
wire n_5849;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_13529;
wire n_6578;
wire n_6224;
wire n_3040;
wire n_8802;
wire n_9859;
wire n_3279;
wire n_14763;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_10879;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_1692;
wire n_1084;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_10639;
wire n_3475;
wire n_3501;
wire n_374;
wire n_1705;
wire n_12554;
wire n_3905;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_13351;
wire n_8121;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_15549;
wire n_10491;
wire n_921;
wire n_12037;
wire n_15371;
wire n_13453;
wire n_579;
wire n_2789;
wire n_5152;
wire n_15080;
wire n_5265;
wire n_12792;
wire n_2257;
wire n_11717;
wire n_9943;
wire n_4927;
wire n_5574;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_7152;
wire n_11723;
wire n_15246;
wire n_2200;
wire n_9575;
wire n_650;
wire n_14940;
wire n_6165;
wire n_9796;
wire n_8320;
wire n_10409;
wire n_1940;
wire n_4548;
wire n_11822;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_1405;
wire n_2376;
wire n_11830;
wire n_12438;
wire n_15395;
wire n_5469;
wire n_14393;
wire n_8766;
wire n_456;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_12838;
wire n_6567;
wire n_9165;
wire n_2670;
wire n_313;
wire n_2700;
wire n_13505;
wire n_14016;
wire n_12323;
wire n_5910;
wire n_15566;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_565;
wire n_3134;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_1569;
wire n_13703;
wire n_3115;
wire n_14369;
wire n_1062;
wire n_7240;
wire n_7570;
wire n_896;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_15354;
wire n_2084;
wire n_4875;
wire n_10476;
wire n_9966;
wire n_13156;
wire n_7817;
wire n_5682;
wire n_15529;
wire n_10710;
wire n_5387;
wire n_654;
wire n_5557;
wire n_411;
wire n_11394;
wire n_2458;
wire n_8850;
wire n_1222;
wire n_11906;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_14647;
wire n_2673;
wire n_2456;
wire n_14298;
wire n_8002;
wire n_9741;
wire n_13897;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_11486;
wire n_1407;
wire n_1795;
wire n_14792;
wire n_15280;
wire n_2871;
wire n_12677;
wire n_420;
wire n_4321;
wire n_10180;
wire n_4183;
wire n_14248;
wire n_14112;
wire n_8370;
wire n_7237;
wire n_164;
wire n_13300;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_9090;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_1271;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_4901;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_12901;
wire n_1640;
wire n_4040;
wire n_10518;
wire n_8301;
wire n_2406;
wire n_12895;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_15170;
wire n_806;
wire n_9771;
wire n_13401;
wire n_584;
wire n_2141;
wire n_15774;
wire n_5316;
wire n_7718;
wire n_244;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_13844;
wire n_14122;
wire n_548;
wire n_7396;
wire n_282;
wire n_10942;
wire n_12668;
wire n_12726;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_833;
wire n_15437;
wire n_13010;
wire n_523;
wire n_6320;
wire n_8126;
wire n_345;
wire n_11239;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4943;
wire n_799;
wire n_10953;
wire n_12432;
wire n_3044;
wire n_4757;
wire n_7561;
wire n_15603;
wire n_7842;
wire n_6810;
wire n_2196;
wire n_2629;
wire n_12352;
wire n_2809;
wire n_787;
wire n_2172;
wire n_6202;
wire n_10099;
wire n_9969;
wire n_11437;
wire n_4682;
wire n_9961;
wire n_12898;
wire n_14068;
wire n_12879;
wire n_14853;
wire n_5564;
wire n_11869;
wire n_13746;
wire n_14895;
wire n_12559;
wire n_13508;
wire n_5620;
wire n_14660;
wire n_15540;
wire n_7163;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_10343;
wire n_2021;
wire n_10836;
wire n_4942;
wire n_15270;
wire n_9899;
wire n_9258;
wire n_159;
wire n_1086;
wire n_13004;
wire n_10181;
wire n_15670;
wire n_10286;
wire n_5406;
wire n_2125;
wire n_8072;
wire n_10371;
wire n_13479;
wire n_14990;
wire n_2561;
wire n_8277;
wire n_7236;
wire n_652;
wire n_4604;
wire n_13117;
wire n_10257;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_7130;
wire n_1241;
wire n_7201;
wire n_11219;
wire n_3157;
wire n_4841;
wire n_14437;
wire n_10047;
wire n_14541;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_13759;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_10949;
wire n_3457;
wire n_4338;
wire n_13766;
wire n_10486;
wire n_11226;
wire n_11282;
wire n_306;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_3005;
wire n_11413;
wire n_3151;
wire n_14700;
wire n_3411;
wire n_15146;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_7491;
wire n_13969;
wire n_5353;
wire n_9995;
wire n_1706;
wire n_13710;
wire n_5186;
wire n_5710;
wire n_9076;
wire n_11232;
wire n_1498;
wire n_12351;
wire n_12693;
wire n_2417;
wire n_9105;
wire n_6792;
wire n_1210;
wire n_12080;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_9316;
wire n_9636;
wire n_5979;
wire n_13359;
wire n_9668;
wire n_3558;
wire n_10372;
wire n_14867;
wire n_7559;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_8867;
wire n_13259;
wire n_9491;
wire n_13335;
wire n_4326;
wire n_6044;
wire n_14022;
wire n_12702;
wire n_1269;
wire n_2083;
wire n_15188;
wire n_2834;
wire n_5517;
wire n_13175;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_2441;
wire n_14954;
wire n_3401;
wire n_10744;
wire n_12648;
wire n_3242;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_655;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_1045;
wire n_5907;
wire n_11334;
wire n_786;
wire n_15757;
wire n_1559;
wire n_13075;
wire n_13736;
wire n_13129;
wire n_6045;
wire n_1872;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_14186;
wire n_7526;
wire n_5040;
wire n_14023;
wire n_6063;
wire n_10736;
wire n_10917;
wire n_1325;
wire n_6504;
wire n_3761;
wire n_11575;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_7004;
wire n_7821;
wire n_14418;
wire n_1727;
wire n_12407;
wire n_13586;
wire n_8308;
wire n_6154;
wire n_11284;
wire n_6943;
wire n_4301;
wire n_10597;
wire n_14668;
wire n_11827;
wire n_151;
wire n_13049;
wire n_3744;
wire n_8165;
wire n_13961;
wire n_14283;
wire n_12038;
wire n_14776;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_15745;
wire n_2041;
wire n_11656;
wire n_8210;
wire n_12644;
wire n_1360;
wire n_10446;
wire n_13134;
wire n_5977;
wire n_11826;
wire n_7879;
wire n_10271;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_15415;
wire n_14808;
wire n_2126;
wire n_7696;
wire n_11570;
wire n_6003;
wire n_12952;
wire n_6684;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_2045;
wire n_14795;
wire n_817;
wire n_9323;
wire n_5451;
wire n_14140;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_9331;
wire n_3621;
wire n_6031;
wire n_9922;
wire n_10170;
wire n_13252;
wire n_11909;
wire n_12024;
wire n_13084;
wire n_8331;
wire n_14479;
wire n_10603;
wire n_12004;
wire n_8217;
wire n_2903;
wire n_6962;
wire n_3216;
wire n_15374;
wire n_332;
wire n_12830;
wire n_12637;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_398;
wire n_4365;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_1882;
wire n_7929;
wire n_10255;
wire n_10572;
wire n_14172;
wire n_3726;
wire n_12009;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_13612;
wire n_1592;
wire n_2719;
wire n_7270;
wire n_591;
wire n_13985;
wire n_11490;
wire n_3758;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_14124;
wire n_2587;
wire n_10113;
wire n_7550;
wire n_15086;
wire n_15077;
wire n_3199;
wire n_12414;
wire n_680;
wire n_9760;
wire n_10690;
wire n_3339;
wire n_6853;
wire n_6742;
wire n_10188;
wire n_13525;
wire n_4923;
wire n_2400;
wire n_10686;
wire n_5864;
wire n_15733;
wire n_9841;
wire n_14997;
wire n_13552;
wire n_6691;
wire n_8743;
wire n_12681;
wire n_7087;
wire n_14207;
wire n_8753;
wire n_1953;
wire n_14799;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_3343;
wire n_12634;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_13863;
wire n_2752;
wire n_8627;
wire n_14305;
wire n_9513;
wire n_14774;
wire n_9863;
wire n_12680;
wire n_15330;
wire n_11613;
wire n_4885;
wire n_13659;
wire n_10233;
wire n_12034;
wire n_751;
wire n_10500;
wire n_15446;
wire n_10555;
wire n_5432;
wire n_15261;
wire n_15492;
wire n_1399;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_11929;
wire n_11075;
wire n_10810;
wire n_7851;
wire n_6894;
wire n_13303;
wire n_13346;
wire n_12176;
wire n_9791;
wire n_13702;
wire n_10311;
wire n_9179;
wire n_2358;
wire n_5453;
wire n_13656;
wire n_3658;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_11177;
wire n_13667;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_10937;
wire n_6817;
wire n_5842;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_400;
wire n_12449;
wire n_337;
wire n_5814;
wire n_2814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_15470;
wire n_11310;
wire n_13275;
wire n_12094;
wire n_6215;
wire n_789;
wire n_3231;
wire n_11165;
wire n_4212;
wire n_9736;
wire n_2979;
wire n_5699;
wire n_181;
wire n_5531;
wire n_14411;
wire n_5765;
wire n_12823;
wire n_2953;
wire n_15412;
wire n_12517;
wire n_6517;
wire n_15754;
wire n_327;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_15441;
wire n_10167;
wire n_7862;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_2946;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_8808;
wire n_10061;
wire n_15257;
wire n_12963;
wire n_10428;
wire n_13087;
wire n_300;
wire n_13972;
wire n_15599;
wire n_11865;
wire n_15436;
wire n_12366;
wire n_15633;
wire n_8528;
wire n_747;
wire n_13024;
wire n_8204;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_14951;
wire n_2565;
wire n_5495;
wire n_10694;
wire n_15646;
wire n_1389;
wire n_12339;
wire n_10602;
wire n_535;
wire n_7100;
wire n_12729;
wire n_3583;
wire n_13292;
wire n_12198;
wire n_3860;
wire n_11041;
wire n_14632;
wire n_9420;
wire n_3851;
wire n_14490;
wire n_5655;
wire n_6393;
wire n_9708;
wire n_14336;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_14738;
wire n_15479;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_8154;
wire n_6966;
wire n_8889;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_13986;
wire n_9790;
wire n_13849;
wire n_13796;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_15522;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_13258;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_7874;
wire n_957;
wire n_1994;
wire n_6035;
wire n_13329;
wire n_7622;
wire n_8490;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_13166;
wire n_15435;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_13946;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_2566;
wire n_14464;
wire n_6364;
wire n_387;
wire n_15028;
wire n_744;
wire n_971;
wire n_8635;
wire n_2702;
wire n_3241;
wire n_7102;
wire n_7420;
wire n_15482;
wire n_2906;
wire n_4342;
wire n_12605;
wire n_13618;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_1258;
wire n_15535;
wire n_2438;
wire n_6253;
wire n_7831;
wire n_2914;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_8532;
wire n_14993;
wire n_14327;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_14097;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_3100;
wire n_2180;
wire n_11140;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_1016;
wire n_8796;
wire n_12218;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_12343;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_12597;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_197;
wire n_4711;
wire n_13744;
wire n_11478;
wire n_12834;
wire n_3068;
wire n_15650;
wire n_10066;
wire n_13017;
wire n_12236;
wire n_14335;
wire n_12902;
wire n_2685;
wire n_6419;
wire n_1083;
wire n_7784;
wire n_9272;
wire n_8372;
wire n_5768;
wire n_3553;
wire n_10088;
wire n_14887;
wire n_13038;
wire n_2275;
wire n_2465;
wire n_7225;
wire n_15199;
wire n_15087;
wire n_8077;
wire n_2568;
wire n_12892;
wire n_2022;
wire n_3811;
wire n_11294;
wire n_910;
wire n_15667;
wire n_3494;
wire n_1721;
wire n_6244;
wire n_6900;
wire n_9812;
wire n_1737;
wire n_9337;
wire n_3486;
wire n_15419;
wire n_4086;
wire n_15219;
wire n_752;
wire n_908;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_9949;
wire n_10289;
wire n_9432;
wire n_1028;
wire n_6942;
wire n_7705;
wire n_11819;
wire n_14889;
wire n_2106;
wire n_2265;
wire n_7228;
wire n_13762;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_7932;
wire n_4409;
wire n_11573;
wire n_9576;
wire n_7509;
wire n_10145;
wire n_13420;
wire n_5872;
wire n_6862;
wire n_14225;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_15053;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_708;
wire n_1973;
wire n_6840;
wire n_13005;
wire n_3181;
wire n_6338;
wire n_14805;
wire n_15267;
wire n_15009;
wire n_8262;
wire n_8423;
wire n_7981;
wire n_1500;
wire n_6037;
wire n_9874;
wire n_9577;
wire n_5700;
wire n_3699;
wire n_12588;
wire n_15648;
wire n_854;
wire n_4913;
wire n_12589;
wire n_2312;
wire n_5874;
wire n_6266;
wire n_14796;
wire n_14143;
wire n_6488;
wire n_904;
wire n_11844;
wire n_709;
wire n_1266;
wire n_2242;
wire n_7164;
wire n_9231;
wire n_8337;
wire n_15390;
wire n_14044;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_185;
wire n_11364;
wire n_3868;
wire n_9569;
wire n_1276;
wire n_13184;
wire n_14823;
wire n_15634;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_14691;
wire n_13535;
wire n_2530;
wire n_14982;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_10009;
wire n_8358;
wire n_14770;
wire n_1085;
wire n_12927;
wire n_9552;
wire n_11100;
wire n_2042;
wire n_9279;
wire n_13822;
wire n_14948;
wire n_11902;
wire n_771;
wire n_6317;
wire n_475;
wire n_924;
wire n_8199;
wire n_298;
wire n_1582;
wire n_492;
wire n_5588;
wire n_11993;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_10443;
wire n_8656;
wire n_10756;
wire n_265;
wire n_7167;
wire n_12813;
wire n_14909;
wire n_6480;
wire n_15105;
wire n_3645;
wire n_14387;
wire n_10918;
wire n_13122;
wire n_13534;
wire n_5075;
wire n_11797;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_12765;
wire n_14106;
wire n_7865;
wire n_15553;
wire n_13616;
wire n_2666;
wire n_1585;
wire n_15690;
wire n_12663;
wire n_10384;
wire n_1799;
wire n_9289;
wire n_2564;
wire n_5085;
wire n_11315;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_2035;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_7134;
wire n_9633;
wire n_15468;
wire n_11153;
wire n_12312;
wire n_3422;
wire n_10074;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_406;
wire n_4845;
wire n_4104;
wire n_9547;
wire n_13097;
wire n_6875;
wire n_13627;
wire n_10934;
wire n_1770;
wire n_10197;
wire n_15786;
wire n_878;
wire n_8346;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_13112;
wire n_8761;
wire n_15458;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_13734;
wire n_8226;
wire n_11949;
wire n_10478;
wire n_8402;
wire n_7079;
wire n_9690;
wire n_9084;
wire n_981;
wire n_5928;
wire n_12256;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_2071;
wire n_11746;
wire n_11812;
wire n_3219;
wire n_9371;
wire n_14051;
wire n_13163;
wire n_3702;
wire n_9711;
wire n_9431;
wire n_8754;
wire n_9847;
wire n_2233;
wire n_4779;
wire n_14650;
wire n_7267;
wire n_481;
wire n_10367;
wire n_14610;
wire n_3233;
wire n_4599;
wire n_12315;
wire n_997;
wire n_11505;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_14100;
wire n_12375;
wire n_12556;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_12998;
wire n_7812;
wire n_1198;
wire n_7103;
wire n_13723;
wire n_13143;
wire n_9080;
wire n_4061;
wire n_14601;
wire n_14549;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_2174;
wire n_436;
wire n_9519;
wire n_14717;
wire n_14814;
wire n_6367;
wire n_3881;
wire n_11363;
wire n_12156;
wire n_13564;
wire n_15794;
wire n_14459;
wire n_13128;
wire n_4508;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_11530;
wire n_12671;
wire n_2426;
wire n_10621;
wire n_14913;
wire n_13411;
wire n_2478;
wire n_7056;
wire n_14645;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_1133;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_13260;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_7813;
wire n_10085;
wire n_15382;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_6080;
wire n_4865;
wire n_12525;
wire n_8182;
wire n_8387;
wire n_1039;
wire n_12076;
wire n_10613;
wire n_10716;
wire n_14090;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_13758;
wire n_7200;
wire n_11359;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_7688;
wire n_4562;
wire n_553;
wire n_3383;
wire n_8707;
wire n_12357;
wire n_15424;
wire n_4903;
wire n_3709;
wire n_10561;
wire n_11434;
wire n_3738;
wire n_9208;
wire n_11791;
wire n_14695;
wire n_15554;
wire n_7611;
wire n_6873;
wire n_15309;
wire n_4186;
wire n_13212;
wire n_14463;
wire n_8494;
wire n_15166;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_15216;
wire n_8544;
wire n_11848;
wire n_13503;
wire n_3610;
wire n_11152;
wire n_4998;
wire n_10749;
wire n_15138;
wire n_3330;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_14166;
wire n_12180;
wire n_2065;
wire n_2879;
wire n_8788;
wire n_15608;
wire n_14405;
wire n_967;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_14081;
wire n_2001;
wire n_7723;
wire n_4341;
wire n_11621;
wire n_679;
wire n_1629;
wire n_10160;
wire n_9327;
wire n_10560;
wire n_7404;
wire n_12857;
wire n_13171;
wire n_5368;
wire n_4263;
wire n_225;
wire n_1260;
wire n_1819;
wire n_309;
wire n_8177;
wire n_3555;
wire n_9854;
wire n_14271;
wire n_12025;
wire n_11667;
wire n_7450;
wire n_7059;
wire n_14854;
wire n_8962;
wire n_915;
wire n_9538;
wire n_14254;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_812;
wire n_12208;
wire n_6145;
wire n_1131;
wire n_11964;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_15266;
wire n_1006;
wire n_13421;
wire n_3110;
wire n_7271;
wire n_1632;
wire n_7826;
wire n_9713;
wire n_14565;
wire n_11298;
wire n_15796;
wire n_13495;
wire n_5933;
wire n_257;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_1311;
wire n_7076;
wire n_13474;
wire n_4780;
wire n_10300;
wire n_13949;
wire n_13314;
wire n_670;
wire n_9588;
wire n_11403;
wire n_14903;
wire n_14218;
wire n_2697;
wire n_11741;
wire n_15107;
wire n_12383;
wire n_11912;
wire n_3908;
wire n_4973;
wire n_15537;
wire n_6842;
wire n_3467;
wire n_12773;
wire n_6866;
wire n_13876;
wire n_14967;
wire n_1887;
wire n_9044;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_9423;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_14487;
wire n_4750;
wire n_14883;
wire n_12962;
wire n_6451;
wire n_9813;
wire n_3039;
wire n_9127;
wire n_14596;
wire n_1226;
wire n_6514;
wire n_3740;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_9244;
wire n_9869;
wire n_11142;
wire n_1958;
wire n_15304;
wire n_315;
wire n_7049;
wire n_5903;
wire n_14449;
wire n_15271;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_12885;
wire n_14865;
wire n_11644;
wire n_2579;
wire n_6345;
wire n_15539;
wire n_2105;
wire n_9715;
wire n_1423;
wire n_8618;
wire n_3387;
wire n_12108;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_364;
wire n_5782;
wire n_7535;
wire n_3420;
wire n_5041;
wire n_13170;
wire n_1915;
wire n_4275;
wire n_10862;
wire n_11531;
wire n_4283;
wire n_4959;
wire n_900;
wire n_8248;
wire n_9056;
wire n_8911;
wire n_11357;
wire n_14471;
wire n_4426;
wire n_9407;
wire n_2912;
wire n_11476;
wire n_14476;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_13633;
wire n_9985;
wire n_15244;
wire n_4449;
wire n_2116;
wire n_12089;
wire n_12496;
wire n_14538;
wire n_2320;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_1013;
wire n_1259;
wire n_11959;
wire n_11367;
wire n_15478;
wire n_2183;
wire n_3002;
wire n_6957;
wire n_9361;
wire n_649;
wire n_1612;
wire n_11921;
wire n_4809;
wire n_8495;
wire n_14532;
wire n_12676;
wire n_13976;
wire n_8783;
wire n_12987;
wire n_13579;
wire n_14557;
wire n_11566;
wire n_1199;
wire n_3392;
wire n_13913;
wire n_8529;
wire n_8733;
wire n_14639;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_625;
wire n_7976;
wire n_6444;
wire n_15392;
wire n_10254;
wire n_14340;
wire n_226;
wire n_14032;
wire n_14715;
wire n_7944;
wire n_13080;
wire n_11208;
wire n_15702;
wire n_7262;
wire n_212;
wire n_3773;
wire n_11374;
wire n_12967;
wire n_13403;
wire n_12452;
wire n_8647;
wire n_2003;
wire n_14899;
wire n_8574;
wire n_1038;
wire n_1581;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_13557;
wire n_12232;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_14952;
wire n_1853;
wire n_11859;
wire n_12818;
wire n_15616;
wire n_15773;
wire n_10386;
wire n_12128;
wire n_6379;
wire n_14060;
wire n_15589;
wire n_798;
wire n_2324;
wire n_14018;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_5563;
wire n_15307;
wire n_245;
wire n_1348;
wire n_13583;
wire n_11026;
wire n_14111;
wire n_8044;
wire n_2977;
wire n_1739;
wire n_13309;
wire n_5840;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9439;
wire n_1380;
wire n_9553;
wire n_11633;
wire n_15292;
wire n_11467;
wire n_2847;
wire n_15239;
wire n_12672;
wire n_2557;
wire n_7506;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_14361;
wire n_8330;
wire n_12760;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_15444;
wire n_13455;
wire n_15560;
wire n_1160;
wire n_883;
wire n_2647;
wire n_15065;
wire n_6232;
wire n_15289;
wire n_9132;
wire n_1032;
wire n_13172;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_9696;
wire n_14943;
wire n_10861;
wire n_2521;
wire n_9120;
wire n_8879;
wire n_15771;
wire n_15508;
wire n_1099;
wire n_11203;
wire n_471;
wire n_11159;
wire n_424;
wire n_8052;
wire n_12168;
wire n_4578;
wire n_2211;
wire n_6362;
wire n_4777;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_14148;
wire n_369;
wire n_8903;
wire n_11030;
wire n_2672;
wire n_4702;
wire n_12590;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_12924;
wire n_5871;
wire n_15605;
wire n_7142;
wire n_141;
wire n_1285;
wire n_12577;
wire n_10182;
wire n_12732;
wire n_1985;
wire n_13928;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_1172;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_10073;
wire n_4531;
wire n_3282;
wire n_11655;
wire n_14619;
wire n_15781;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_11017;
wire n_12843;
wire n_7247;
wire n_14279;
wire n_14448;
wire n_12069;
wire n_10419;
wire n_7241;
wire n_7172;
wire n_15656;
wire n_3106;
wire n_1140;
wire n_15427;
wire n_1670;
wire n_14622;
wire n_10333;
wire n_2344;
wire n_12430;
wire n_10317;
wire n_2365;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_14739;
wire n_15687;
wire n_375;
wire n_7235;
wire n_11248;
wire n_2447;
wire n_8540;
wire n_12613;
wire n_12270;
wire n_14365;
wire n_6239;
wire n_9915;
wire n_4617;
wire n_2340;
wire n_9325;
wire n_9196;
wire n_13407;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_13676;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_13788;
wire n_14555;
wire n_11141;
wire n_5105;
wire n_12695;
wire n_15467;
wire n_10893;
wire n_1572;
wire n_4308;
wire n_11093;
wire n_5021;
wire n_14219;
wire n_9251;
wire n_3463;
wire n_11576;
wire n_8939;
wire n_13584;
wire n_428;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_15471;
wire n_2510;
wire n_1954;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_8468;
wire n_822;
wire n_7657;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_13181;
wire n_5134;
wire n_7096;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_12210;
wire n_13327;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_8778;
wire n_11197;
wire n_491;
wire n_3998;
wire n_7442;
wire n_15047;
wire n_1591;
wire n_3632;
wire n_10093;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_1344;
wire n_15014;
wire n_6174;
wire n_15428;
wire n_12006;
wire n_2730;
wire n_2495;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_14168;
wire n_6087;
wire n_371;
wire n_7593;
wire n_12246;
wire n_5249;
wire n_14085;
wire n_2603;
wire n_2090;
wire n_8068;
wire n_15342;
wire n_9955;
wire n_15534;
wire n_538;
wire n_3829;
wire n_10539;
wire n_14080;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_10107;
wire n_13975;
wire n_5969;
wire n_3655;
wire n_10196;
wire n_10121;
wire n_8198;
wire n_493;
wire n_14573;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_13085;
wire n_2108;
wire n_15536;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_1211;
wire n_13224;
wire n_11469;
wire n_6454;
wire n_5022;
wire n_12625;
wire n_9270;
wire n_14046;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_14142;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_14512;
wire n_8557;
wire n_1280;
wire n_6918;
wire n_6041;
wire n_9099;
wire n_12389;
wire n_13761;
wire n_9309;
wire n_3296;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_15097;
wire n_10814;
wire n_5276;
wire n_9627;
wire n_13971;
wire n_11252;
wire n_8012;
wire n_14456;
wire n_13364;
wire n_1445;
wire n_7672;
wire n_11494;
wire n_2551;
wire n_6664;
wire n_1526;
wire n_5047;
wire n_14743;
wire n_196;
wire n_7318;
wire n_2985;
wire n_1978;
wire n_6472;
wire n_10218;
wire n_574;
wire n_8114;
wire n_13131;
wire n_14941;
wire n_3792;
wire n_4202;
wire n_12995;
wire n_14406;
wire n_1446;
wire n_3938;
wire n_13209;
wire n_4791;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_14859;
wire n_5879;
wire n_14563;
wire n_8062;
wire n_4403;
wire n_11883;
wire n_5238;
wire n_11256;
wire n_11832;
wire n_14959;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_12370;
wire n_3531;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_15387;
wire n_473;
wire n_10975;
wire n_11901;
wire n_6352;
wire n_12974;
wire n_1054;
wire n_9460;
wire n_559;
wire n_8542;
wire n_12136;
wire n_10859;
wire n_13078;
wire n_7063;
wire n_1956;
wire n_7047;
wire n_11652;
wire n_14768;
wire n_4139;
wire n_14320;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_14807;
wire n_13885;
wire n_6238;
wire n_15795;
wire n_1986;
wire n_10542;
wire n_8038;
wire n_13631;
wire n_13932;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_10681;
wire n_15162;
wire n_15606;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_11572;
wire n_13370;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_11894;
wire n_3603;
wire n_14493;
wire n_10222;
wire n_6724;
wire n_13113;
wire n_13387;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_813;
wire n_11583;
wire n_11336;
wire n_8716;
wire n_6705;
wire n_3822;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_4163;
wire n_818;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_14764;
wire n_645;
wire n_8734;
wire n_3812;
wire n_3910;
wire n_9204;
wire n_9476;
wire n_7074;
wire n_11849;
wire n_12142;
wire n_9689;
wire n_15237;
wire n_2633;
wire n_10659;
wire n_6591;
wire n_2207;
wire n_7585;
wire n_4948;
wire n_12564;
wire n_5268;
wire n_13643;
wire n_9780;
wire n_6946;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_13433;
wire n_2198;
wire n_3319;
wire n_15505;
wire n_541;
wire n_10403;
wire n_13607;
wire n_12983;
wire n_15538;
wire n_2073;
wire n_2273;
wire n_6289;
wire n_7037;
wire n_3748;
wire n_13697;
wire n_3272;
wire n_11784;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_3396;
wire n_14244;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_15541;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_12886;
wire n_1162;
wire n_14114;
wire n_13980;
wire n_6532;
wire n_4372;
wire n_821;
wire n_1068;
wire n_7293;
wire n_13000;
wire n_982;
wire n_12035;
wire n_14362;
wire n_13006;
wire n_5640;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_14742;
wire n_408;
wire n_932;
wire n_4318;
wire n_2831;
wire n_6778;
wire n_4158;
wire n_14904;
wire n_3978;
wire n_3317;
wire n_6721;
wire n_5560;
wire n_13205;
wire n_6644;
wire n_2123;
wire n_1697;
wire n_6512;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_12810;
wire n_6108;
wire n_10370;
wire n_8258;
wire n_4918;
wire n_3824;
wire n_9597;
wire n_5067;
wire n_13820;
wire n_13947;
wire n_11322;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_11892;
wire n_12122;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_15283;
wire n_13428;
wire n_354;
wire n_5841;
wire n_12241;
wire n_12396;
wire n_15407;
wire n_9343;
wire n_7614;
wire n_15731;
wire n_2941;
wire n_1278;
wire n_547;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_9837;
wire n_1396;
wire n_11421;
wire n_11057;
wire n_634;
wire n_2355;
wire n_4147;
wire n_10969;
wire n_10896;
wire n_136;
wire n_4477;
wire n_11966;
wire n_14474;
wire n_12748;
wire n_3168;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_10562;
wire n_5941;
wire n_2009;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_1793;
wire n_14417;
wire n_3601;
wire n_5611;
wire n_10355;
wire n_10054;
wire n_3092;
wire n_1289;
wire n_6219;
wire n_3055;
wire n_6706;
wire n_7479;
wire n_3966;
wire n_12571;
wire n_11853;
wire n_9692;
wire n_2866;
wire n_7395;
wire n_10598;
wire n_13034;
wire n_13402;
wire n_8947;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_9609;
wire n_11118;
wire n_10717;
wire n_10029;
wire n_15494;
wire n_1703;
wire n_7078;
wire n_2580;
wire n_13831;
wire n_8188;
wire n_6761;
wire n_882;
wire n_8972;
wire n_10007;
wire n_3649;
wire n_11751;
wire n_2821;
wire n_11423;
wire n_1875;
wire n_11725;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_13635;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_12674;
wire n_8510;
wire n_11410;
wire n_3384;
wire n_12230;
wire n_15698;
wire n_9567;
wire n_14637;
wire n_1950;
wire n_6811;
wire n_9061;
wire n_1563;
wire n_11495;
wire n_3419;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_7372;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_12220;
wire n_674;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_922;
wire n_10704;
wire n_1335;
wire n_11520;
wire n_11622;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_12169;
wire n_12283;
wire n_12336;
wire n_7174;
wire n_14783;
wire n_13268;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_13383;
wire n_10457;
wire n_12543;
wire n_15088;
wire n_702;
wire n_4965;
wire n_347;
wire n_8021;
wire n_3346;
wire n_9705;
wire n_7803;
wire n_15124;
wire n_1896;
wire n_11012;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_14158;
wire n_12595;
wire n_9624;
wire n_3861;
wire n_9701;
wire n_675;
wire n_11502;
wire n_14236;
wire n_15348;
wire n_11429;
wire n_1540;
wire n_15802;
wire n_1977;
wire n_15163;
wire n_10389;
wire n_11631;
wire n_13588;
wire n_13510;
wire n_13570;
wire n_14640;
wire n_3891;
wire n_2193;
wire n_6659;
wire n_15688;
wire n_4523;
wire n_1655;
wire n_9709;
wire n_13677;
wire n_13983;
wire n_242;
wire n_6011;
wire n_9416;
wire n_1886;
wire n_9295;
wire n_13757;
wire n_14036;
wire n_4371;
wire n_6225;
wire n_11842;
wire n_14710;
wire n_12463;
wire n_10990;
wire n_2994;
wire n_11640;
wire n_5502;
wire n_12263;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_877;
wire n_9929;
wire n_12920;
wire n_10264;
wire n_5850;
wire n_13317;
wire n_4673;
wire n_13910;
wire n_15029;
wire n_2519;
wire n_9953;
wire n_13737;
wire n_7086;
wire n_728;
wire n_3415;
wire n_1063;
wire n_6648;
wire n_4607;
wire n_14286;
wire n_15578;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_12717;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_598;
wire n_12141;
wire n_8584;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_13196;
wire n_13520;
wire n_15363;
wire n_437;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_697;
wire n_10301;
wire n_3271;
wire n_295;
wire n_5088;
wire n_14955;
wire n_4248;
wire n_8034;
wire n_388;
wire n_13018;
wire n_484;
wire n_7025;
wire n_9364;
wire n_8228;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_15139;
wire n_8076;
wire n_6826;
wire n_1825;
wire n_1757;
wire n_170;
wire n_1792;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_15642;
wire n_9836;
wire n_1412;
wire n_2497;
wire n_10929;
wire n_14357;
wire n_9107;
wire n_3809;
wire n_11279;
wire n_11724;
wire n_13044;
wire n_11789;
wire n_14152;
wire n_3139;
wire n_13228;
wire n_11525;
wire n_13518;
wire n_13862;
wire n_11999;
wire n_4070;
wire n_13446;
wire n_8100;
wire n_13086;
wire n_10837;
wire n_3545;
wire n_14869;
wire n_3885;
wire n_1369;
wire n_14008;
wire n_881;
wire n_10554;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_12746;
wire n_4031;
wire n_5837;
wire n_148;
wire n_4675;
wire n_10149;
wire n_10970;
wire n_7768;
wire n_2663;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_14651;
wire n_5491;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_7982;
wire n_15791;
wire n_12190;
wire n_14927;
wire n_12787;
wire n_8804;
wire n_13881;
wire n_15484;
wire n_297;
wire n_3337;
wire n_11383;
wire n_12799;
wire n_15152;
wire n_4002;
wire n_11847;
wire n_11976;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_12657;
wire n_9317;
wire n_2165;
wire n_9769;
wire n_5547;
wire n_15205;
wire n_13747;
wire n_1391;
wire n_8158;
wire n_12511;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_6879;
wire n_12532;
wire n_1295;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_10102;
wire n_3477;
wire n_8433;
wire n_8765;
wire n_2349;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_8213;
wire n_5983;
wire n_3146;
wire n_1495;
wire n_14472;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_10534;
wire n_11825;
wire n_585;
wire n_4653;
wire n_4435;
wire n_10932;
wire n_10619;
wire n_7684;
wire n_11049;
wire n_14354;
wire n_14974;
wire n_15532;
wire n_5604;
wire n_1756;
wire n_8451;
wire n_1128;
wire n_5411;
wire n_673;
wire n_12743;
wire n_8334;
wire n_4019;
wire n_1071;
wire n_8731;
wire n_10589;
wire n_11681;
wire n_11611;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_11202;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_15587;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_865;
wire n_3616;
wire n_9748;
wire n_7370;
wire n_5815;
wire n_13365;
wire n_15254;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_8539;
wire n_10205;
wire n_2151;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_14618;
wire n_1839;
wire n_2341;
wire n_15747;
wire n_9226;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_10110;
wire n_2707;
wire n_13899;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_11688;
wire n_6888;
wire n_826;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_12715;
wire n_1714;
wire n_11709;
wire n_12434;
wire n_14328;
wire n_12628;
wire n_8122;
wire n_718;
wire n_6095;
wire n_13444;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_14209;
wire n_542;
wire n_11331;
wire n_14429;
wire n_5311;
wire n_305;
wire n_12979;
wire n_9528;
wire n_6590;
wire n_14348;
wire n_2089;
wire n_10638;
wire n_7583;
wire n_12201;
wire n_14086;
wire n_3522;
wire n_6559;
wire n_12499;
wire n_2747;
wire n_3924;
wire n_9112;
wire n_15799;
wire n_12448;
wire n_791;
wire n_4621;
wire n_4216;
wire n_11876;
wire n_5797;
wire n_510;
wire n_9235;
wire n_10610;
wire n_11187;
wire n_4240;
wire n_12761;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_13852;
wire n_9333;
wire n_704;
wire n_2148;
wire n_7151;
wire n_15004;
wire n_4162;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_8950;
wire n_2339;
wire n_14089;
wire n_10758;
wire n_2861;
wire n_13431;
wire n_10190;
wire n_1999;
wire n_2731;
wire n_622;
wire n_5520;
wire n_147;
wire n_3353;
wire n_11804;
wire n_14234;
wire n_3975;
wire n_3018;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_1838;
wire n_6287;
wire n_2638;
wire n_12809;
wire n_13614;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_14552;
wire n_7353;
wire n_2002;
wire n_12538;
wire n_9330;
wire n_14208;
wire n_2138;
wire n_14025;
wire n_7758;
wire n_4021;
wire n_2414;
wire n_13779;
wire n_12446;
wire n_9490;
wire n_3014;
wire n_15693;
wire n_1771;
wire n_2316;
wire n_12029;
wire n_4103;
wire n_11052;
wire n_9355;
wire n_5060;
wire n_9523;
wire n_14584;
wire n_3148;
wire n_15386;
wire n_4022;
wire n_4986;
wire n_14620;
wire n_5888;
wire n_5669;
wire n_14575;
wire n_9574;
wire n_9024;
wire n_11694;
wire n_5772;
wire n_15349;
wire n_7571;
wire n_9582;
wire n_145;
wire n_2208;
wire n_4775;
wire n_10060;
wire n_5884;
wire n_6671;
wire n_13470;
wire n_11009;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_9288;
wire n_9686;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_13068;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_11446;
wire n_10910;
wire n_1304;
wire n_10162;
wire n_294;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_15002;
wire n_2134;
wire n_1176;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_13248;
wire n_7792;
wire n_13842;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_15338;
wire n_15378;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_425;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_1431;
wire n_14501;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_2958;
wire n_10014;
wire n_8703;
wire n_15723;
wire n_7109;
wire n_12642;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_8822;
wire n_14790;
wire n_14999;
wire n_10677;
wire n_12187;
wire n_657;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_12321;
wire n_5924;
wire n_1505;
wire n_9992;
wire n_290;
wire n_11247;
wire n_15180;
wire n_15692;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_12669;
wire n_13106;
wire n_3129;
wire n_8476;
wire n_14296;
wire n_14294;
wire n_6702;
wire n_11927;
wire n_3620;
wire n_13720;
wire n_11179;
wire n_478;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_14862;
wire n_2520;
wire n_13706;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_13903;
wire n_3693;
wire n_446;
wire n_9051;
wire n_10385;
wire n_11514;
wire n_4497;
wire n_7749;
wire n_10078;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_10105;
wire n_12470;
wire n_12994;
wire n_15785;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_8705;
wire n_14574;
wire n_10215;
wire n_526;
wire n_14451;
wire n_11779;
wire n_2251;
wire n_14059;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_14211;
wire n_15234;
wire n_10834;
wire n_293;
wire n_7574;
wire n_1070;
wire n_2403;
wire n_14092;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_14509;
wire n_1665;
wire n_4306;
wire n_14394;
wire n_11882;
wire n_13516;
wire n_11647;
wire n_154;
wire n_4224;
wire n_12064;
wire n_15027;
wire n_14273;
wire n_15404;
wire n_10706;
wire n_2127;
wire n_12462;
wire n_3341;
wire n_6005;
wire n_8872;
wire n_12696;
wire n_4453;
wire n_9555;
wire n_15735;
wire n_11133;
wire n_3559;
wire n_5449;
wire n_14845;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_15230;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_12735;
wire n_7713;
wire n_15465;
wire n_4564;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_11222;
wire n_9200;
wire n_5146;
wire n_10709;
wire n_3056;
wire n_745;
wire n_2424;
wire n_12646;
wire n_3201;
wire n_10871;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_10304;
wire n_6936;
wire n_2589;
wire n_4535;
wire n_14624;
wire n_10244;
wire n_15036;
wire n_14765;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_14120;
wire n_14995;
wire n_755;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_527;
wire n_2442;
wire n_7641;
wire n_13794;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_7203;
wire n_12999;
wire n_13537;
wire n_14260;
wire n_14407;
wire n_9397;
wire n_1137;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_12682;
wire n_3612;
wire n_9673;
wire n_14434;
wire n_14175;
wire n_14802;
wire n_4695;
wire n_6848;
wire n_2545;
wire n_8642;
wire n_3509;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11875;
wire n_11941;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_14834;
wire n_12111;
wire n_15780;
wire n_8912;
wire n_14346;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_13463;
wire n_7439;
wire n_1314;
wire n_600;
wire n_9496;
wire n_3196;
wire n_15189;
wire n_8110;
wire n_864;
wire n_14275;
wire n_5319;
wire n_2504;
wire n_10796;
wire n_14506;
wire n_2623;
wire n_10016;
wire n_9008;
wire n_12903;
wire n_12079;
wire n_15335;
wire n_399;
wire n_6343;
wire n_12593;
wire n_1440;
wire n_14615;
wire n_5270;
wire n_2063;
wire n_10030;
wire n_15227;
wire n_15222;
wire n_8805;
wire n_1534;
wire n_6850;
wire n_12864;
wire n_15285;
wire n_5005;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_13294;
wire n_15689;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_7209;
wire n_6014;
wire n_7112;
wire n_15026;
wire n_13895;
wire n_1339;
wire n_2475;
wire n_11307;
wire n_5181;
wire n_13936;
wire n_13933;
wire n_6979;
wire n_7815;
wire n_13222;
wire n_403;
wire n_7934;
wire n_9545;
wire n_723;
wire n_3144;
wire n_13813;
wire n_8111;
wire n_3244;
wire n_596;
wire n_9629;
wire n_9603;
wire n_11578;
wire n_6865;
wire n_10432;
wire n_1141;
wire n_1268;
wire n_12719;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_15361;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_8739;
wire n_6747;
wire n_9674;
wire n_13714;
wire n_2357;
wire n_2025;
wire n_5583;
wire n_4654;
wire n_13438;
wire n_6433;
wire n_10462;
wire n_12725;
wire n_3640;
wire n_642;
wire n_1159;
wire n_995;
wire n_3481;
wire n_6640;
wire n_15469;
wire n_11769;
wire n_8856;
wire n_2250;
wire n_3033;
wire n_303;
wire n_6142;
wire n_9930;
wire n_11908;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_14901;
wire n_6462;
wire n_7769;
wire n_14988;
wire n_2374;
wire n_416;
wire n_1681;
wire n_6034;
wire n_520;
wire n_9781;
wire n_418;
wire n_10291;
wire n_13159;
wire n_4597;
wire n_9659;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_14333;
wire n_7233;
wire n_13636;
wire n_8732;
wire n_13506;
wire n_13287;
wire n_11913;
wire n_14788;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_14590;
wire n_11341;
wire n_1618;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_13389;
wire n_10669;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_14603;
wire n_8231;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_5061;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_13905;
wire n_1653;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_4063;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_4237;
wire n_2601;
wire n_13717;
wire n_5029;
wire n_5127;
wire n_12317;
wire n_13302;
wire n_6071;
wire n_2920;
wire n_773;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_15119;
wire n_920;
wire n_1374;
wire n_10185;
wire n_8908;
wire n_11182;
wire n_2648;
wire n_3212;
wire n_10092;
wire n_15768;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_1169;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_1617;
wire n_12782;
wire n_3370;
wire n_3386;
wire n_335;
wire n_4721;
wire n_15256;
wire n_11231;
wire n_14145;
wire n_463;
wire n_3093;
wire n_8090;
wire n_13740;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_848;
wire n_12875;
wire n_274;
wire n_15064;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_13918;
wire n_8137;
wire n_7045;
wire n_13775;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_3169;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_9987;
wire n_1806;
wire n_10983;
wire n_15218;
wire n_15452;
wire n_7984;
wire n_11727;
wire n_13615;
wire n_15625;
wire n_6788;
wire n_2023;
wire n_7014;
wire n_12192;
wire n_12633;
wire n_2720;
wire n_2204;
wire n_496;
wire n_10430;
wire n_14779;
wire n_15114;
wire n_8305;
wire n_4614;
wire n_177;
wire n_3360;
wire n_2087;
wire n_10277;
wire n_1636;
wire n_14973;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_1323;
wire n_6709;
wire n_14465;
wire n_13412;
wire n_2627;
wire n_4422;
wire n_960;
wire n_10948;
wire n_11749;
wire n_6550;
wire n_6712;
wire n_10525;
wire n_9507;
wire n_14287;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_15296;
wire n_778;
wire n_3004;
wire n_8841;
wire n_14553;
wire n_3870;
wire n_13457;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_15136;
wire n_1764;
wire n_6743;
wire n_12497;
wire n_4632;
wire n_15043;
wire n_10354;
wire n_1610;
wire n_12412;
wire n_3084;
wire n_11880;
wire n_5785;
wire n_2343;
wire n_793;
wire n_7465;
wire n_14528;
wire n_13177;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_12724;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_14958;
wire n_15551;
wire n_6672;
wire n_9457;
wire n_2942;
wire n_4966;
wire n_9485;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_13940;
wire n_2515;
wire n_7936;
wire n_8966;
wire n_316;
wire n_6084;
wire n_11249;
wire n_1551;
wire n_15449;
wire n_4847;
wire n_10287;
wire n_4054;
wire n_11039;
wire n_8538;
wire n_7738;
wire n_14342;
wire n_2555;
wire n_12101;
wire n_10119;
wire n_13693;
wire n_11145;
wire n_3586;
wire n_12606;
wire n_11986;
wire n_3653;
wire n_8395;
wire n_10900;
wire n_14798;
wire n_5966;
wire n_2201;
wire n_725;
wire n_10349;
wire n_6634;
wire n_14107;
wire n_14758;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_8961;
wire n_14781;
wire n_10849;
wire n_7462;
wire n_13333;
wire n_4635;
wire n_368;
wire n_13229;
wire n_994;
wire n_12118;
wire n_5735;
wire n_13311;
wire n_14409;
wire n_14724;
wire n_7490;
wire n_11380;
wire n_2278;
wire n_15737;
wire n_14291;
wire n_7545;
wire n_1020;
wire n_10792;
wire n_15573;
wire n_11513;
wire n_13296;
wire n_8625;
wire n_1273;
wire n_9809;
wire n_7160;
wire n_8937;
wire n_4214;
wire n_7464;
wire n_6919;
wire n_14611;
wire n_10750;
wire n_13756;
wire n_3448;
wire n_7805;
wire n_10995;
wire n_617;
wire n_13092;
wire n_7295;
wire n_7115;
wire n_2924;
wire n_12087;
wire n_9192;
wire n_13675;
wire n_1036;
wire n_15022;
wire n_3595;
wire n_14338;
wire n_7348;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_10537;
wire n_421;
wire n_11861;
wire n_3991;
wire n_15051;
wire n_6548;
wire n_15394;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_8511;
wire n_1095;
wire n_6993;
wire n_6973;
wire n_12081;
wire n_1270;
wire n_10426;
wire n_4405;
wire n_610;
wire n_4413;
wire n_9558;
wire n_11594;
wire n_1852;
wire n_7453;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_15639;
wire n_4036;
wire n_10684;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_3670;
wire n_2381;
wire n_11436;
wire n_12346;
wire n_2052;
wire n_179;
wire n_4667;
wire n_5081;
wire n_517;
wire n_11729;
wire n_4182;
wire n_15039;
wire n_667;
wire n_3230;
wire n_8371;
wire n_8702;
wire n_13916;
wire n_15195;
wire n_8116;
wire n_1279;
wire n_1115;
wire n_7946;
wire n_8195;
wire n_1499;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_14069;
wire n_12244;
wire n_504;
wire n_1409;
wire n_5877;
wire n_9991;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_11366;
wire n_11872;
wire n_8845;
wire n_7681;
wire n_15198;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_13620;
wire n_5189;
wire n_1503;
wire n_13930;
wire n_7702;
wire n_6676;
wire n_13981;
wire n_2819;
wire n_8149;
wire n_10823;
wire n_3041;
wire n_4637;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_11516;
wire n_14766;
wire n_603;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_8392;
wire n_9560;
wire n_14592;
wire n_8095;
wire n_7210;
wire n_14659;
wire n_5869;
wire n_10830;
wire n_15109;
wire n_2439;
wire n_11132;
wire n_2404;
wire n_1182;
wire n_6718;
wire n_15007;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_4155;
wire n_6854;
wire n_4238;
wire n_3011;
wire n_15400;
wire n_2061;
wire n_15197;
wire n_2757;
wire n_15485;
wire n_4977;
wire n_167;
wire n_14841;
wire n_13624;
wire n_5632;
wire n_8519;
wire n_14277;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_1216;
wire n_13493;
wire n_2716;
wire n_6032;
wire n_9047;
wire n_13805;
wire n_12953;
wire n_2452;
wire n_12842;
wire n_15224;
wire n_3650;
wire n_8968;
wire n_12481;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_5446;
wire n_11316;
wire n_3010;
wire n_7855;
wire n_14029;
wire n_3043;
wire n_11047;
wire n_14963;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_4590;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_14648;
wire n_3137;
wire n_11767;
wire n_9599;
wire n_14056;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_13866;
wire n_3177;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_13695;
wire n_12435;
wire n_10340;
wire n_10946;
wire n_9428;
wire n_11586;
wire n_6981;
wire n_15344;
wire n_13288;
wire n_2220;
wire n_7065;
wire n_2577;
wire n_12149;
wire n_13669;
wire n_9216;
wire n_1262;
wire n_3238;
wire n_218;
wire n_3529;
wire n_12002;
wire n_12836;
wire n_4835;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_13840;
wire n_11229;
wire n_13548;
wire n_15710;
wire n_2232;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_14251;
wire n_4038;
wire n_6122;
wire n_11397;
wire n_11225;
wire n_2790;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_4565;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_4159;
wire n_12840;
wire n_3784;
wire n_7330;
wire n_14605;
wire n_5437;
wire n_8883;
wire n_220;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_1608;
wire n_7336;
wire n_11471;
wire n_2373;
wire n_1472;
wire n_14705;
wire n_7446;
wire n_13543;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_10577;
wire n_13772;
wire n_800;
wire n_14679;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_15487;
wire n_7357;
wire n_1491;
wire n_8756;
wire n_11324;
wire n_8737;
wire n_1840;
wire n_13925;
wire n_10334;
wire n_4434;
wire n_12945;
wire n_13406;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_2244;
wire n_10151;
wire n_14040;
wire n_11614;
wire n_4290;
wire n_6439;
wire n_8602;
wire n_14054;
wire n_2586;
wire n_1684;
wire n_13368;
wire n_2446;
wire n_1346;
wire n_12850;
wire n_14507;
wire n_13469;
wire n_8240;
wire n_7714;
wire n_1352;
wire n_5407;
wire n_10411;
wire n_15242;
wire n_13249;
wire n_9484;
wire n_12984;
wire n_10989;
wire n_2017;
wire n_8422;
wire n_3029;
wire n_10939;
wire n_13587;
wire n_12224;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_1046;
wire n_2560;
wire n_9394;
wire n_9305;
wire n_9999;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_8878;
wire n_11144;
wire n_10090;
wire n_7440;
wire n_11361;
wire n_14857;
wire n_1102;
wire n_1963;
wire n_6406;
wire n_6945;
wire n_14872;
wire n_8112;
wire n_258;
wire n_14034;
wire n_11567;
wire n_3790;
wire n_10962;
wire n_7029;
wire n_2766;
wire n_260;
wire n_14797;
wire n_11128;
wire n_9622;
wire n_9292;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_356;
wire n_12197;
wire n_14177;
wire n_14093;
wire n_10186;
wire n_3318;
wire n_14607;
wire n_4833;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_6618;
wire n_13326;
wire n_6474;
wire n_13082;
wire n_14453;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_4888;
wire n_13094;
wire n_10856;
wire n_12403;
wire n_7317;
wire n_776;
wire n_321;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_6000;
wire n_2782;
wire n_12679;
wire n_13481;
wire n_9584;
wire n_3977;
wire n_227;
wire n_9461;
wire n_11168;
wire n_8055;
wire n_13692;
wire n_8194;
wire n_14921;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_12018;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_8360;
wire n_6425;
wire n_1456;
wire n_14457;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_9845;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_14382;
wire n_14389;
wire n_11937;
wire n_12872;
wire n_13396;
wire n_7522;
wire n_6492;
wire n_2229;
wire n_10071;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_11460;
wire n_14517;
wire n_2099;
wire n_13713;
wire n_8251;
wire n_5323;
wire n_11565;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_14621;
wire n_3184;
wire n_12372;
wire n_9618;
wire n_14911;
wire n_6118;
wire n_13608;
wire n_5810;
wire n_4561;
wire n_15405;
wire n_4461;
wire n_464;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_11192;
wire n_11808;
wire n_4007;
wire n_15643;
wire n_13257;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_15420;
wire n_2642;
wire n_4239;
wire n_8677;
wire n_13052;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_14934;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_13914;
wire n_1319;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_14663;
wire n_2986;
wire n_5702;
wire n_10035;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_2536;
wire n_3915;
wire n_139;
wire n_14962;
wire n_1633;
wire n_15652;
wire n_13922;
wire n_9699;
wire n_13423;
wire n_12340;
wire n_3489;
wire n_13277;
wire n_8108;
wire n_2835;
wire n_14578;
wire n_8736;
wire n_15653;
wire n_5914;
wire n_1416;
wire n_5243;
wire n_2820;
wire n_2293;
wire n_12955;
wire n_12068;
wire n_10252;
wire n_5250;
wire n_11555;
wire n_3074;
wire n_13494;
wire n_6869;
wire n_3102;
wire n_10041;
wire n_9321;
wire n_15499;
wire n_14625;
wire n_5590;
wire n_10345;
wire n_14514;
wire n_2026;
wire n_1282;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_550;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_14256;
wire n_15016;
wire n_10543;
wire n_275;
wire n_2727;
wire n_3377;
wire n_7924;
wire n_560;
wire n_4782;
wire n_12394;
wire n_13578;
wire n_1321;
wire n_7659;
wire n_2533;
wire n_569;
wire n_3530;
wire n_9161;
wire n_9005;
wire n_14204;
wire n_2869;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_1235;
wire n_2759;
wire n_12954;
wire n_7836;
wire n_2361;
wire n_10737;
wire n_1292;
wire n_12662;
wire n_15697;
wire n_2266;
wire n_4876;
wire n_14082;
wire n_10464;
wire n_6146;
wire n_346;
wire n_14688;
wire n_7280;
wire n_10644;
wire n_12801;
wire n_13448;
wire n_8504;
wire n_5813;
wire n_9293;
wire n_12503;
wire n_13708;
wire n_10365;
wire n_13767;
wire n_790;
wire n_5833;
wire n_11781;
wire n_2611;
wire n_2901;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_15728;
wire n_14832;
wire n_15202;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_2653;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_299;
wire n_1248;
wire n_12965;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_14571;
wire n_902;
wire n_2189;
wire n_2246;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_15707;
wire n_431;
wire n_5816;
wire n_3156;
wire n_10809;
wire n_15396;
wire n_8927;
wire n_10899;
wire n_15347;
wire n_672;
wire n_9639;
wire n_15155;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_15250;
wire n_6228;
wire n_6711;
wire n_1941;
wire n_3483;
wire n_11884;
wire n_5416;
wire n_8946;
wire n_11997;
wire n_14881;
wire n_13090;
wire n_14527;
wire n_12822;
wire n_706;
wire n_1794;
wire n_1236;
wire n_13541;
wire n_13307;
wire n_13371;
wire n_11863;
wire n_4493;
wire n_4924;
wire n_7971;
wire n_7279;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_743;
wire n_766;
wire n_12264;
wire n_13312;
wire n_11761;
wire n_430;
wire n_1746;
wire n_9984;
wire n_8474;
wire n_3524;
wire n_7275;
wire n_8232;
wire n_489;
wire n_2885;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_636;
wire n_9649;
wire n_14703;
wire n_8904;
wire n_11199;
wire n_13533;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_10629;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_660;
wire n_2062;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_8382;
wire n_4421;
wire n_13023;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_2839;
wire n_9501;
wire n_11896;
wire n_2856;
wire n_4793;
wire n_13856;
wire n_15607;
wire n_4498;
wire n_10006;
wire n_2070;
wire n_7259;
wire n_11757;
wire n_12320;
wire n_1607;
wire n_12274;
wire n_14588;
wire n_1454;
wire n_15315;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_12622;
wire n_11185;
wire n_12659;
wire n_2348;
wire n_2944;
wire n_13440;
wire n_8128;
wire n_6818;
wire n_6992;
wire n_3831;
wire n_15226;
wire n_15746;
wire n_869;
wire n_1154;
wire n_13436;
wire n_646;
wire n_528;
wire n_391;
wire n_10206;
wire n_1329;
wire n_6322;
wire n_5167;
wire n_15425;
wire n_5661;
wire n_5932;
wire n_5830;
wire n_3589;
wire n_262;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_897;
wire n_846;
wire n_2066;
wire n_7539;
wire n_841;
wire n_1476;
wire n_12586;
wire n_3391;
wire n_12629;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_508;
wire n_1800;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_1463;
wire n_10275;
wire n_11081;
wire n_13011;
wire n_3458;
wire n_7775;
wire n_8481;
wire n_4505;
wire n_11392;
wire n_9981;
wire n_3190;
wire n_1562;
wire n_14858;
wire n_7930;
wire n_5558;
wire n_1826;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_13911;
wire n_5383;
wire n_14495;
wire n_5126;
wire n_1759;
wire n_14165;
wire n_8205;
wire n_5051;
wire n_9907;
wire n_13088;
wire n_5587;
wire n_12269;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_13538;
wire n_6976;
wire n_853;
wire n_7640;
wire n_14617;
wire n_13701;
wire n_9816;
wire n_13787;
wire n_10498;
wire n_875;
wire n_11424;
wire n_13486;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_1678;
wire n_13674;
wire n_14263;
wire n_11463;
wire n_13912;
wire n_14303;
wire n_10292;
wire n_661;
wire n_7969;
wire n_6864;
wire n_11278;
wire n_14445;
wire n_8605;
wire n_10358;
wire n_3787;
wire n_1256;
wire n_7548;
wire n_3585;
wire n_10635;
wire n_13626;
wire n_3565;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_12913;
wire n_12832;
wire n_5025;
wire n_933;
wire n_8067;
wire n_6998;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_12301;
wire n_3135;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_14427;
wire n_1217;
wire n_7197;
wire n_5645;
wire n_9676;
wire n_3990;
wire n_11881;
wire n_7393;
wire n_11332;
wire n_6917;
wire n_13629;
wire n_6937;
wire n_7591;
wire n_13207;
wire n_310;
wire n_1628;
wire n_14980;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_2109;
wire n_7727;
wire n_7358;
wire n_988;
wire n_2796;
wire n_7324;
wire n_2507;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_11935;
wire n_13589;
wire n_15730;
wire n_4534;
wire n_15685;
wire n_1536;
wire n_6301;
wire n_9788;
wire n_1204;
wire n_1132;
wire n_6929;
wire n_15570;
wire n_233;
wire n_15562;
wire n_11309;
wire n_1327;
wire n_8719;
wire n_955;
wire n_8045;
wire n_10785;
wire n_7729;
wire n_13872;
wire n_246;
wire n_2787;
wire n_2969;
wire n_15493;
wire n_2395;
wire n_12341;
wire n_12615;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_14475;
wire n_8209;
wire n_13357;
wire n_10802;
wire n_14477;
wire n_769;
wire n_2380;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_1120;
wire n_6699;
wire n_12926;
wire n_14809;
wire n_9213;
wire n_555;
wire n_4579;
wire n_7291;
wire n_14725;
wire n_7631;
wire n_14522;
wire n_669;
wire n_8784;
wire n_2290;
wire n_7382;
wire n_4811;
wire n_13869;
wire n_2048;
wire n_13955;
wire n_176;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_2005;
wire n_13561;
wire n_12167;
wire n_14720;
wire n_9473;
wire n_14400;
wire n_4857;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_15019;
wire n_6677;
wire n_12161;
wire n_13499;
wire n_3432;
wire n_12085;
wire n_14843;
wire n_2736;
wire n_2883;
wire n_11735;
wire n_1408;
wire n_7618;
wire n_4282;
wire n_1196;
wire n_10647;
wire n_3493;
wire n_10523;
wire n_9320;
wire n_8769;
wire n_6764;
wire n_13554;
wire n_8575;
wire n_12298;
wire n_10081;
wire n_863;
wire n_3774;
wire n_5733;
wire n_10324;
wire n_6780;
wire n_11189;
wire n_8815;
wire n_11582;
wire n_12569;
wire n_2910;
wire n_14929;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_748;
wire n_3268;
wire n_1785;
wire n_9303;
wire n_1147;
wire n_11105;
wire n_1754;
wire n_3057;
wire n_11705;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_2584;
wire n_7673;
wire n_13698;
wire n_1812;
wire n_6830;
wire n_866;
wire n_13894;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_7282;
wire n_2287;
wire n_452;
wire n_6586;
wire n_9968;
wire n_10808;
wire n_11474;
wire n_10474;
wire n_6333;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_761;
wire n_15466;
wire n_13595;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_13943;
wire n_2492;
wire n_7953;
wire n_13540;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_14642;
wire n_9722;
wire n_13283;
wire n_12042;
wire n_12155;
wire n_14827;
wire n_5657;
wire n_15481;
wire n_174;
wire n_1173;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_13465;
wire n_8695;
wire n_4974;
wire n_12373;
wire n_15615;
wire n_5975;
wire n_15664;
wire n_4911;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_4436;
wire n_14579;
wire n_8363;
wire n_15388;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_1174;
wire n_13733;
wire n_13098;
wire n_8665;
wire n_6510;
wire n_8282;
wire n_3334;
wire n_9388;
wire n_5938;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_12654;
wire n_14141;
wire n_5602;
wire n_647;
wire n_11992;
wire n_9379;
wire n_5097;
wire n_15790;
wire n_844;
wire n_4985;
wire n_7751;
wire n_2117;
wire n_2234;
wire n_10869;
wire n_3823;
wire n_14880;
wire n_14718;
wire n_4384;
wire n_14975;
wire n_2741;
wire n_3114;
wire n_13142;
wire n_7581;
wire n_13180;
wire n_888;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_15217;
wire n_2203;
wire n_14589;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_10453;
wire n_236;
wire n_12386;
wire n_14257;
wire n_4858;
wire n_4678;
wire n_13308;
wire n_9952;
wire n_2649;
wire n_3556;
wire n_15323;
wire n_9911;
wire n_12183;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_414;
wire n_1922;
wire n_15187;
wire n_10668;
wire n_9256;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_13785;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_1215;
wire n_12964;
wire n_839;
wire n_10473;
wire n_15712;
wire n_14007;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_15099;
wire n_8493;
wire n_10331;
wire n_7346;
wire n_11439;
wire n_14655;
wire n_779;
wire n_1537;
wire n_10957;
wire n_13373;
wire n_2205;
wire n_4243;
wire n_13517;
wire n_7579;
wire n_12863;
wire n_10352;
wire n_4025;
wire n_11188;
wire n_7428;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_12221;
wire n_4059;
wire n_9195;
wire n_10442;
wire n_1509;
wire n_11687;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_8870;
wire n_13973;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_11774;
wire n_4313;
wire n_4142;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_7015;
wire n_6475;
wire n_3982;
wire n_8507;
wire n_7283;
wire n_7699;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_13206;
wire n_9623;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_7249;
wire n_10713;
wire n_5546;
wire n_3796;
wire n_232;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_14102;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_10954;
wire n_13637;
wire n_4246;
wire n_12267;
wire n_15803;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_13941;
wire n_13978;
wire n_4532;
wire n_15339;
wire n_13439;
wire n_228;
wire n_13780;
wire n_8893;
wire n_1525;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_14133;
wire n_2594;
wire n_14433;
wire n_11329;
wire n_6495;
wire n_7194;
wire n_5994;
wire n_9516;
wire n_4244;
wire n_2147;
wire n_13241;
wire n_592;
wire n_13187;
wire n_13162;
wire n_2503;
wire n_4049;
wire n_6752;
wire n_1156;
wire n_12768;
wire n_8976;
wire n_6426;
wire n_2600;
wire n_984;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_15059;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_11661;
wire n_8156;
wire n_7494;
wire n_868;
wire n_4353;
wire n_11120;
wire n_14923;
wire n_9222;
wire n_735;
wire n_13031;
wire n_8882;
wire n_6350;
wire n_8435;
wire n_4787;
wire n_7736;
wire n_10622;
wire n_5633;
wire n_13661;
wire n_13155;
wire n_9546;
wire n_469;
wire n_1218;
wire n_5664;
wire n_7589;
wire n_14259;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_15673;
wire n_13410;
wire n_4537;
wire n_14012;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_357;
wire n_13066;
wire n_8660;
wire n_2429;
wire n_13360;
wire n_11296;
wire n_13665;
wire n_8479;
wire n_985;
wire n_14214;
wire n_15558;
wire n_13770;
wire n_12993;
wire n_2440;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_3521;
wire n_11314;
wire n_8723;
wire n_13511;
wire n_802;
wire n_11019;
wire n_561;
wire n_8606;
wire n_9663;
wire n_980;
wire n_2681;
wire n_6235;
wire n_7843;
wire n_15678;
wire n_8235;
wire n_13083;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_12647;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_15340;
wire n_9820;
wire n_14569;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_14071;
wire n_1244;
wire n_1685;
wire n_9743;
wire n_6496;
wire n_3066;
wire n_15744;
wire n_7756;
wire n_2844;
wire n_12749;
wire n_15557;
wire n_8940;
wire n_8342;
wire n_2303;
wire n_1619;
wire n_13048;
wire n_11584;
wire n_2285;
wire n_5280;
wire n_8448;
wire n_13563;
wire n_14154;
wire n_7700;
wire n_4451;
wire n_14169;
wire n_8472;
wire n_4332;
wire n_810;
wire n_7555;
wire n_10000;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_2742;
wire n_10582;
wire n_12066;
wire n_12812;
wire n_3695;
wire n_10427;
wire n_12060;
wire n_11816;
wire n_3976;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_14174;
wire n_3563;
wire n_6513;
wire n_10246;
wire n_2367;
wire n_7500;
wire n_11910;
wire n_15377;
wire n_201;
wire n_3198;
wire n_11693;
wire n_3495;
wire n_15583;
wire n_1034;
wire n_15429;
wire n_13347;
wire n_14269;
wire n_5925;
wire n_2909;
wire n_9248;
wire n_754;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_9822;
wire n_10835;
wire n_975;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_13991;
wire n_13823;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_14821;
wire n_13323;
wire n_3359;
wire n_12164;
wire n_15096;
wire n_5272;
wire n_11368;
wire n_14992;
wire n_10125;
wire n_12824;
wire n_13111;
wire n_13434;
wire n_6330;
wire n_15563;
wire n_10117;
wire n_9065;
wire n_467;
wire n_3187;
wire n_12716;
wire n_10844;
wire n_14153;
wire n_3218;
wire n_8457;
wire n_6802;
wire n_13456;
wire n_10654;
wire n_9153;
wire n_9086;
wire n_10505;
wire n_9339;
wire n_582;
wire n_10198;
wire n_861;
wire n_7157;
wire n_6909;
wire n_11064;
wire n_13237;
wire n_6908;
wire n_857;
wire n_14312;
wire n_8237;
wire n_13445;
wire n_15448;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_15045;
wire n_11409;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_7266;
wire n_15760;
wire n_2221;
wire n_8046;
wire n_588;
wire n_14746;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_13284;
wire n_12437;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_10840;
wire n_12052;
wire n_6477;
wire n_9746;
wire n_14606;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_1166;
wire n_15501;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_15751;
wire n_15298;
wire n_11533;
wire n_11605;
wire n_2709;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_534;
wire n_7198;
wire n_1578;
wire n_8335;
wire n_1861;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_10144;
wire n_9440;
wire n_3955;
wire n_9684;
wire n_15741;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_14793;
wire n_730;
wire n_6184;
wire n_5817;
wire n_5214;
wire n_15486;
wire n_203;
wire n_10973;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_13472;
wire n_2162;
wire n_15596;
wire n_1868;
wire n_207;
wire n_2079;
wire n_9493;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_15475;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_3433;
wire n_11330;
wire n_12720;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_205;
wire n_2185;
wire n_6038;
wire n_10551;
wire n_13318;
wire n_15379;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_10553;
wire n_2774;
wire n_13127;
wire n_14884;
wire n_3162;
wire n_1274;
wire n_8309;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_15121;
wire n_12687;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_14075;
wire n_1899;
wire n_9032;
wire n_9814;
wire n_6313;
wire n_784;
wire n_4804;
wire n_6112;
wire n_5619;
wire n_13208;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_13867;
wire n_15594;
wire n_5859;
wire n_12325;
wire n_14423;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_13443;
wire n_862;
wire n_5776;
wire n_8166;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_2813;
wire n_14626;
wire n_1935;
wire n_5826;
wire n_15766;
wire n_2027;
wire n_10108;
wire n_2091;
wire n_8960;
wire n_13865;
wire n_12789;
wire n_5920;
wire n_2991;
wire n_10307;
wire n_5030;
wire n_14530;
wire n_15402;
wire n_4194;
wire n_7994;
wire n_1449;
wire n_14206;
wire n_4703;
wire n_8443;
wire n_361;
wire n_7349;
wire n_8657;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_2419;
wire n_6180;
wire n_14481;
wire n_8683;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_2677;
wire n_15044;
wire n_12127;
wire n_12504;
wire n_12382;
wire n_3182;
wire n_5756;
wire n_15306;
wire n_12602;
wire n_3283;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_13673;
wire n_12062;
wire n_14119;
wire n_1742;
wire n_4030;
wire n_12573;

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_39),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_37),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_29),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_23),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_15),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_26),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_103),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_51),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_65),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_36),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_114),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_85),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_54),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_42),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_49),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_30),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_48),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_98),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_58),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_80),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_0),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_32),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_99),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_95),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_104),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_74),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_2),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_18),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_92),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_21),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_106),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_61),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_72),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_24),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_35),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_82),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_31),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_84),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_132),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_131),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_113),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_75),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_78),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_6),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_27),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_1),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_62),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_25),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_33),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_96),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_47),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_77),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_59),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_57),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_76),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_102),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_136),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_139),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_237),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_143),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_148),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_166),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_193),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_216),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_141),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_151),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_147),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_160),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_171),
.B(n_2),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_161),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_164),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_173),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_174),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_178),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_198),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_217),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_184),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_198),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_208),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_251),
.B(n_3),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_152),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_181),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_189),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_218),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_187),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_283),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_302),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_277),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_286),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_309),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_309),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_303),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_299),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_186),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_275),
.B(n_225),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_310),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_281),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_297),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_298),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_308),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_226),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_282),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_159),
.B1(n_201),
.B2(n_170),
.Y(n_362)
);

OAI22x1_ASAP7_75t_R g363 ( 
.A1(n_315),
.A2(n_260),
.B1(n_244),
.B2(n_268),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_140),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_343),
.A2(n_177),
.B1(n_137),
.B2(n_212),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_149),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_213),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_314),
.B(n_306),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_215),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_253),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_320),
.A2(n_232),
.B1(n_197),
.B2(n_222),
.Y(n_383)
);

CKINVDCx8_ASAP7_75t_R g384 ( 
.A(n_341),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_314),
.B(n_205),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_304),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_259),
.B(n_256),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_140),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_230),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_255),
.B(n_200),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_265),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_153),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_140),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_235),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_193),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_314),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_314),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_321),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_154),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_321),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_314),
.B(n_199),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_314),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_324),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_353),
.B(n_155),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_314),
.B(n_241),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_156),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_343),
.A2(n_206),
.B1(n_267),
.B2(n_266),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_343),
.B(n_157),
.Y(n_431)
);

AOI22x1_ASAP7_75t_L g432 ( 
.A1(n_351),
.A2(n_248),
.B1(n_246),
.B2(n_228),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_314),
.B(n_142),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_343),
.B(n_269),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_314),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_316),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_316),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_349),
.A2(n_162),
.B1(n_264),
.B2(n_204),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_359),
.A2(n_202),
.B(n_262),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_333),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_343),
.B(n_169),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_316),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_316),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_316),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_314),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_343),
.A2(n_183),
.B1(n_261),
.B2(n_258),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_343),
.A2(n_182),
.B1(n_257),
.B2(n_254),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_349),
.Y(n_450)
);

CKINVDCx6p67_ASAP7_75t_R g451 ( 
.A(n_319),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_314),
.B(n_196),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_314),
.B(n_191),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_343),
.B(n_176),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_316),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_314),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_314),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_314),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_314),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_316),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_333),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_343),
.B(n_203),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_333),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_343),
.B(n_175),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_314),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_324),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_314),
.B(n_263),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_343),
.B(n_207),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_343),
.B(n_169),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_353),
.B(n_172),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_353),
.B(n_211),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_324),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_316),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_324),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_314),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_316),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_343),
.A2(n_233),
.B1(n_252),
.B2(n_250),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_324),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_321),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_321),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_316),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_325),
.B(n_194),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_316),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_343),
.A2(n_190),
.B1(n_249),
.B2(n_245),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_314),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_349),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_314),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_314),
.B(n_185),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_343),
.B(n_180),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_343),
.B(n_158),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_417),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_422),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_451),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_R g497 ( 
.A(n_481),
.B(n_239),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_482),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_384),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_375),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_370),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_400),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_361),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_224),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_400),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_402),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_382),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_361),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_467),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_410),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_383),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_410),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_402),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_367),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_367),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_414),
.B(n_179),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_408),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_408),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_412),
.B(n_168),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_362),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_366),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_371),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_405),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_366),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_450),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_R g533 ( 
.A(n_484),
.B(n_167),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_454),
.B(n_214),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_411),
.B(n_165),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_381),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_450),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_377),
.B(n_380),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_488),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_459),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_440),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_488),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_419),
.A2(n_428),
.B1(n_491),
.B2(n_469),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_363),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_388),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_376),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_404),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_416),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_416),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_420),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_392),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_447),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_457),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_457),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_470),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_385),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_487),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_470),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_R g561 ( 
.A(n_407),
.B(n_220),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_413),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_424),
.B(n_238),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_489),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_231),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_444),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_462),
.B(n_243),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_385),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_489),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_R g571 ( 
.A(n_430),
.B(n_242),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_398),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_423),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_445),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_423),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_396),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_438),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_435),
.B(n_223),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_456),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_R g580 ( 
.A(n_458),
.B(n_221),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_394),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_466),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_387),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_477),
.B(n_227),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_429),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_449),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_479),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_465),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_372),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_409),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_409),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_452),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_448),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_372),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_387),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_486),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_386),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_403),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_399),
.B(n_240),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_396),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_406),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_390),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_492),
.A2(n_236),
.B1(n_234),
.B2(n_229),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

INVxp67_ASAP7_75t_R g606 ( 
.A(n_418),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_406),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_364),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_R g609 ( 
.A(n_368),
.B(n_73),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_426),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_365),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_472),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_369),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_461),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_406),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_473),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_464),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_391),
.B(n_263),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_452),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_373),
.B(n_378),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_433),
.B(n_169),
.Y(n_621)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_453),
.B(n_56),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_453),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_490),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_490),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_378),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_415),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_464),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_441),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_379),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_441),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_441),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_433),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_421),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_436),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_471),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_471),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_471),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_427),
.B(n_263),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_R g640 ( 
.A(n_395),
.B(n_55),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_437),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_427),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_395),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_442),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_395),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_443),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_446),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_455),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_460),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_463),
.B(n_3),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_475),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_483),
.B(n_8),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_393),
.A2(n_198),
.B(n_43),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_485),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_432),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_432),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_468),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_439),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_393),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_439),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_401),
.Y(n_662)
);

CKINVDCx16_ASAP7_75t_R g663 ( 
.A(n_401),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_417),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_R g665 ( 
.A(n_417),
.B(n_52),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_434),
.B(n_198),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_417),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_R g668 ( 
.A(n_417),
.B(n_105),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_417),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_414),
.B(n_108),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_451),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_R g672 ( 
.A(n_417),
.B(n_121),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_374),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_417),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_383),
.B(n_10),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_374),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_417),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_451),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_417),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_363),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_417),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_451),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_417),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_417),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_417),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_459),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_374),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_451),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_R g689 ( 
.A(n_408),
.B(n_198),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_370),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_374),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_370),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_451),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_374),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_374),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_417),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_370),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_417),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_R g699 ( 
.A(n_417),
.B(n_198),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_417),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_376),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_451),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_383),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_370),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_370),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_451),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_R g707 ( 
.A(n_417),
.B(n_422),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_451),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_416),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_374),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_R g711 ( 
.A(n_408),
.B(n_341),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_414),
.B(n_424),
.Y(n_712)
);

CKINVDCx6p67_ASAP7_75t_R g713 ( 
.A(n_451),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_417),
.B(n_422),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_434),
.B(n_454),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_417),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_409),
.B(n_407),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_417),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_451),
.Y(n_719)
);

INVxp33_ASAP7_75t_L g720 ( 
.A(n_363),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_434),
.B(n_454),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_374),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_374),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_417),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_417),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_382),
.B(n_419),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_451),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_417),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_R g729 ( 
.A(n_408),
.B(n_341),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_370),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_374),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_417),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_417),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_417),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_417),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_451),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_417),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_374),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_417),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_417),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_417),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_451),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_374),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_370),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_376),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_434),
.B(n_454),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_451),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_376),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_417),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_451),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_451),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_397),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_374),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_451),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_397),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_417),
.B(n_422),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_428),
.A2(n_462),
.B(n_431),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_417),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_451),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_417),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_417),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_374),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_374),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_374),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_376),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_370),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_417),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_417),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_414),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_414),
.B(n_424),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_R g771 ( 
.A(n_417),
.B(n_422),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_417),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_370),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_417),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_417),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_370),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_451),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_374),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_417),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_451),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_374),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_370),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_374),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_417),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_451),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_376),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_417),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_374),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_417),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_381),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_451),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_417),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_434),
.B(n_454),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_R g794 ( 
.A(n_417),
.B(n_422),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_451),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_451),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_374),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_374),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_451),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_451),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_374),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_370),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_715),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_712),
.B(n_770),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_504),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_519),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_612),
.B(n_572),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_544),
.B(n_514),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_511),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_528),
.B(n_755),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_746),
.A2(n_721),
.B1(n_757),
.B2(n_661),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_498),
.B(n_752),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_519),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_548),
.B(n_538),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_527),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_530),
.B(n_543),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_541),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_566),
.B(n_568),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_707),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_565),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_536),
.B(n_790),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_567),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_574),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_585),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_605),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_614),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

OAI22x1_ASAP7_75t_L g828 ( 
.A1(n_524),
.A2(n_529),
.B1(n_675),
.B2(n_577),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_610),
.B(n_616),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_628),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_576),
.B(n_521),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_549),
.Y(n_832)
);

AND2x6_ASAP7_75t_L g833 ( 
.A(n_662),
.B(n_660),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_596),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_606),
.B(n_726),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_599),
.B(n_594),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_597),
.B(n_600),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_502),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_690),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_525),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_596),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_590),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_596),
.B(n_633),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_692),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_586),
.B(n_587),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_697),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_595),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_506),
.B(n_757),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_550),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_496),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_501),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_505),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_704),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_633),
.B(n_646),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_769),
.B(n_507),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_705),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_512),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_588),
.B(n_510),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_647),
.B(n_649),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_552),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_518),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_625),
.B(n_549),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_554),
.B(n_555),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_712),
.B(n_770),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_526),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_730),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_531),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_493),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_545),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_689),
.Y(n_870)
);

AND2x6_ASAP7_75t_L g871 ( 
.A(n_670),
.B(n_633),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_549),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_655),
.B(n_620),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_709),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_709),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_673),
.B(n_676),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_687),
.B(n_691),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_694),
.B(n_695),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_532),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_670),
.B(n_710),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_709),
.Y(n_881)
);

INVx6_ASAP7_75t_L g882 ( 
.A(n_569),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_717),
.B(n_656),
.Y(n_883)
);

INVx4_ASAP7_75t_SL g884 ( 
.A(n_717),
.Y(n_884)
);

BUFx8_ASAP7_75t_SL g885 ( 
.A(n_509),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_711),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_591),
.B(n_592),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_703),
.A2(n_537),
.B1(n_539),
.B2(n_680),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_722),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_723),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_731),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_556),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_738),
.B(n_743),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_753),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_557),
.B(n_560),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_583),
.B(n_686),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_762),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_744),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_533),
.B(n_579),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_583),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_564),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_766),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_663),
.A2(n_622),
.B1(n_659),
.B2(n_666),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_657),
.A2(n_781),
.B1(n_801),
.B2(n_763),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_570),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_558),
.B(n_642),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_582),
.B(n_602),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_764),
.A2(n_798),
.B1(n_778),
.B2(n_797),
.Y(n_908)
);

AND2x6_ASAP7_75t_L g909 ( 
.A(n_783),
.B(n_788),
.Y(n_909)
);

INVx4_ASAP7_75t_SL g910 ( 
.A(n_717),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_773),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_714),
.Y(n_912)
);

BUFx8_ASAP7_75t_SL g913 ( 
.A(n_495),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_618),
.B(n_534),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_776),
.A2(n_802),
.B1(n_782),
.B2(n_621),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_546),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_540),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_542),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_553),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_547),
.B(n_701),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_520),
.B(n_639),
.Y(n_921)
);

NOR2x1p5_ASAP7_75t_L g922 ( 
.A(n_713),
.B(n_517),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_547),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_756),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_701),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_581),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_589),
.A2(n_717),
.B1(n_601),
.B2(n_644),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_607),
.B(n_615),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_745),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_748),
.B(n_765),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_520),
.B(n_639),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_513),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_522),
.B(n_494),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_515),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_593),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_499),
.B(n_664),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_748),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_765),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

NAND3xp33_ASAP7_75t_L g941 ( 
.A(n_667),
.B(n_792),
.C(n_725),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_608),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_771),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_786),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_669),
.B(n_674),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_630),
.B(n_598),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_699),
.B(n_603),
.Y(n_947)
);

INVx4_ASAP7_75t_SL g948 ( 
.A(n_621),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_794),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_619),
.B(n_623),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_677),
.B(n_679),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_641),
.B(n_611),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_613),
.B(n_627),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_551),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_L g955 ( 
.A(n_629),
.B(n_631),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_634),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_593),
.Y(n_957)
);

AND2x6_ASAP7_75t_L g958 ( 
.A(n_635),
.B(n_648),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_651),
.B(n_652),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_654),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_559),
.Y(n_961)
);

BUFx10_ASAP7_75t_L g962 ( 
.A(n_681),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_562),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_650),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_653),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_683),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_684),
.B(n_685),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_658),
.Y(n_968)
);

OAI22xp33_ASAP7_75t_L g969 ( 
.A1(n_624),
.A2(n_637),
.B1(n_632),
.B2(n_636),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_604),
.A2(n_638),
.B1(n_626),
.B2(n_645),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_729),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_696),
.B(n_698),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_671),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_563),
.Y(n_974)
);

INVx6_ASAP7_75t_L g975 ( 
.A(n_678),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_571),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_700),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_643),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_500),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_716),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_573),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_682),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_497),
.B(n_561),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_578),
.B(n_584),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_640),
.A2(n_609),
.B1(n_672),
.B2(n_668),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_575),
.B(n_789),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_718),
.B(n_741),
.C(n_740),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_724),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_728),
.B(n_749),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_732),
.B(n_787),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_580),
.B(n_535),
.Y(n_991)
);

NAND3xp33_ASAP7_75t_L g992 ( 
.A(n_733),
.B(n_767),
.C(n_737),
.Y(n_992)
);

AND2x6_ASAP7_75t_L g993 ( 
.A(n_665),
.B(n_784),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_523),
.B(n_779),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_734),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_735),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_688),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_739),
.B(n_758),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_760),
.B(n_775),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_761),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_768),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_772),
.B(n_774),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_503),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_693),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_720),
.B(n_516),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_508),
.B(n_702),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_706),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_708),
.B(n_719),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_727),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_736),
.B(n_742),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_747),
.B(n_750),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_800),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_751),
.Y(n_1013)
);

BUFx10_ASAP7_75t_L g1014 ( 
.A(n_754),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_759),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_777),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_780),
.B(n_785),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_791),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_795),
.B(n_796),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_799),
.B(n_793),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_528),
.B(n_399),
.Y(n_1021)
);

AND2x6_ASAP7_75t_L g1022 ( 
.A(n_793),
.B(n_662),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_SL g1023 ( 
.A(n_519),
.Y(n_1023)
);

INVx6_ASAP7_75t_L g1024 ( 
.A(n_519),
.Y(n_1024)
);

BUFx4_ASAP7_75t_L g1025 ( 
.A(n_707),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_504),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_793),
.B(n_721),
.C(n_715),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_504),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_793),
.B(n_715),
.Y(n_1029)
);

INVxp33_ASAP7_75t_L g1030 ( 
.A(n_707),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_504),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_504),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_504),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_504),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_712),
.B(n_770),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_519),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_504),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_793),
.B(n_715),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_528),
.B(n_399),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_504),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_712),
.B(n_770),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_504),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_528),
.B(n_399),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_596),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_793),
.B(n_715),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_712),
.B(n_770),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_504),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_793),
.B(n_715),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_793),
.B(n_715),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_596),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_528),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_665),
.B(n_668),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_504),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_793),
.B(n_715),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_504),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_793),
.B(n_746),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_793),
.B(n_715),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_596),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_519),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_612),
.B(n_362),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_525),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_793),
.B(n_715),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_596),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_793),
.B(n_715),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_793),
.B(n_662),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_519),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_596),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_528),
.B(n_399),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_504),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_528),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_793),
.B(n_715),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_793),
.B(n_662),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_504),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_793),
.B(n_715),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_793),
.B(n_746),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_596),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_504),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_793),
.B(n_715),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_519),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_793),
.B(n_715),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_504),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_504),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_596),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_504),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_493),
.B(n_494),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_596),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_596),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_793),
.B(n_715),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_504),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_793),
.B(n_715),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_519),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_504),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_504),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_793),
.B(n_715),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_596),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_504),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_519),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_528),
.B(n_410),
.Y(n_1100)
);

BUFx8_ASAP7_75t_SL g1101 ( 
.A(n_509),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_793),
.B(n_746),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_793),
.A2(n_721),
.B1(n_715),
.B2(n_746),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_596),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_504),
.Y(n_1105)
);

INVx4_ASAP7_75t_SL g1106 ( 
.A(n_717),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_793),
.B(n_715),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_519),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_528),
.B(n_399),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_793),
.B(n_715),
.Y(n_1110)
);

AND2x6_ASAP7_75t_L g1111 ( 
.A(n_793),
.B(n_662),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_528),
.B(n_399),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_504),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_504),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_712),
.B(n_770),
.Y(n_1115)
);

OAI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_715),
.A2(n_721),
.B1(n_793),
.B2(n_543),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_519),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_504),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_504),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_519),
.Y(n_1121)
);

AND2x6_ASAP7_75t_L g1122 ( 
.A(n_793),
.B(n_662),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_504),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_493),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_504),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_504),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_504),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_596),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_528),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_793),
.B(n_715),
.Y(n_1130)
);

CKINVDCx11_ASAP7_75t_R g1131 ( 
.A(n_509),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_793),
.B(n_715),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_504),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_504),
.Y(n_1134)
);

INVx4_ASAP7_75t_SL g1135 ( 
.A(n_717),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_504),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_519),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_793),
.B(n_715),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_612),
.B(n_362),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_793),
.B(n_715),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_519),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_793),
.B(n_746),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_528),
.B(n_399),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_528),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_504),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_519),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_793),
.B(n_715),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_793),
.B(n_715),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_519),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_596),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_519),
.Y(n_1151)
);

XNOR2xp5_ASAP7_75t_L g1152 ( 
.A(n_675),
.B(n_315),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_528),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_707),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_528),
.B(n_399),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1156)
);

AND2x6_ASAP7_75t_L g1157 ( 
.A(n_793),
.B(n_662),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_528),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_504),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_504),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_504),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_793),
.B(n_715),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_504),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_519),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_596),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_528),
.B(n_399),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_712),
.B(n_770),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_493),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_504),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_528),
.B(n_399),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_519),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_712),
.B(n_770),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_504),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_504),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_596),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_504),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_596),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_R g1179 ( 
.A(n_524),
.B(n_529),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_504),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_793),
.B(n_715),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_528),
.B(n_399),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_519),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_528),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_504),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_793),
.B(n_746),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_504),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_504),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_596),
.Y(n_1189)
);

INVx4_ASAP7_75t_SL g1190 ( 
.A(n_717),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_519),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_793),
.B(n_746),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_596),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_596),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_793),
.B(n_715),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_793),
.B(n_715),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_712),
.B(n_770),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_504),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_793),
.B(n_715),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_596),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_596),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_793),
.B(n_715),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_793),
.B(n_715),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_793),
.A2(n_715),
.B1(n_721),
.B2(n_746),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_528),
.B(n_399),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_504),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_793),
.B(n_715),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_793),
.B(n_715),
.Y(n_1209)
);

AND2x6_ASAP7_75t_L g1210 ( 
.A(n_793),
.B(n_662),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_525),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_519),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_528),
.B(n_399),
.Y(n_1213)
);

INVxp33_ASAP7_75t_L g1214 ( 
.A(n_707),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_596),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_504),
.Y(n_1216)
);

INVx6_ASAP7_75t_L g1217 ( 
.A(n_519),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_793),
.B(n_715),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_793),
.A2(n_721),
.B1(n_715),
.B2(n_746),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_793),
.B(n_715),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_793),
.B(n_715),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_596),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_612),
.B(n_362),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_519),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_793),
.B(n_715),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_504),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_504),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_504),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_504),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_793),
.A2(n_746),
.B1(n_721),
.B2(n_715),
.Y(n_1230)
);

BUFx8_ASAP7_75t_SL g1231 ( 
.A(n_509),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_504),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_715),
.A2(n_721),
.B1(n_793),
.B2(n_543),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_596),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_596),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_793),
.B(n_746),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_715),
.B(n_721),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_519),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_504),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_519),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_504),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_793),
.B(n_715),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_504),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_504),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_R g1245 ( 
.A(n_879),
.B(n_1062),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_803),
.B(n_1029),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1049),
.B(n_1072),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_805),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1075),
.B(n_1081),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_809),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_L g1252 ( 
.A(n_880),
.B(n_818),
.Y(n_1252)
);

INVx8_ASAP7_75t_L g1253 ( 
.A(n_1100),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1095),
.B(n_1130),
.Y(n_1254)
);

NOR3xp33_ASAP7_75t_L g1255 ( 
.A(n_837),
.B(n_1195),
.C(n_1148),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1256)
);

AOI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1242),
.A2(n_1205),
.B1(n_1048),
.B2(n_1054),
.C(n_1045),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1038),
.B(n_1057),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_814),
.B(n_1103),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_804),
.B(n_864),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_817),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1059),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_842),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1063),
.B(n_1065),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1027),
.A2(n_1097),
.B1(n_1120),
.B2(n_1060),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1021),
.B(n_1039),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_847),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_850),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1219),
.B(n_1156),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_851),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1079),
.B(n_1089),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1091),
.B(n_1107),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1173),
.B(n_1201),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1110),
.B(n_1132),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1044),
.Y(n_1275)
);

INVx8_ASAP7_75t_L g1276 ( 
.A(n_1100),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1086),
.B(n_967),
.Y(n_1277)
);

NOR3xp33_ASAP7_75t_L g1278 ( 
.A(n_836),
.B(n_859),
.C(n_1138),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1230),
.B(n_870),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_820),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1140),
.B(n_1147),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1162),
.B(n_1181),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1196),
.B(n_1203),
.C(n_1199),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_822),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1044),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_R g1286 ( 
.A(n_1179),
.B(n_819),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_852),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_824),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_857),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1059),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_861),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_865),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1209),
.B(n_1220),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_825),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_869),
.Y(n_1296)
);

AND2x6_ASAP7_75t_SL g1297 ( 
.A(n_972),
.B(n_989),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1225),
.B(n_1237),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_821),
.Y(n_1299)
);

BUFx5_ASAP7_75t_L g1300 ( 
.A(n_833),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_807),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1056),
.B(n_1076),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1102),
.B(n_1142),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_889),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_924),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1186),
.B(n_1192),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_873),
.B(n_816),
.Y(n_1307)
);

AND2x2_ASAP7_75t_SL g1308 ( 
.A(n_971),
.B(n_808),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1236),
.B(n_964),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_904),
.B(n_845),
.C(n_829),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_991),
.B(n_968),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_L g1312 ( 
.A(n_880),
.B(n_871),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_890),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_811),
.A2(n_985),
.B1(n_965),
.B2(n_903),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_840),
.B(n_867),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_886),
.B(n_858),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1044),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1022),
.B(n_1066),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1022),
.B(n_1066),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_984),
.B(n_835),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_908),
.B(n_1069),
.C(n_1043),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_891),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_894),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1051),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1176),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1022),
.B(n_1066),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1073),
.B(n_1111),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1073),
.B(n_1111),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_974),
.B(n_976),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_949),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_897),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_826),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1143),
.B(n_1155),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1073),
.B(n_1111),
.Y(n_1335)
);

NAND2x1_ASAP7_75t_L g1336 ( 
.A(n_871),
.B(n_833),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_876),
.A2(n_877),
.B(n_893),
.C(n_878),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_SL g1338 ( 
.A(n_983),
.B(n_1154),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1002),
.B(n_937),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_830),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1028),
.Y(n_1342)
);

XNOR2xp5_ASAP7_75t_L g1343 ( 
.A(n_1152),
.B(n_982),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1214),
.B(n_1061),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1139),
.B(n_1223),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1182),
.B(n_1206),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_918),
.B(n_1213),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1176),
.B(n_901),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1176),
.B(n_990),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_L g1351 ( 
.A(n_887),
.B(n_934),
.C(n_831),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1152),
.A2(n_828),
.B1(n_888),
.B2(n_912),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_855),
.B(n_880),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_871),
.B(n_925),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1071),
.B(n_1129),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_815),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1032),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_953),
.A2(n_1040),
.B1(n_1047),
.B2(n_1037),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_810),
.B(n_812),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_930),
.B(n_938),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_944),
.B(n_823),
.Y(n_1361)
);

OAI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_863),
.A2(n_895),
.B(n_1158),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_990),
.B(n_994),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_827),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_804),
.B(n_864),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_892),
.B(n_945),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1042),
.B(n_1053),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1055),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1093),
.B(n_1098),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1184),
.B(n_980),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1070),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_899),
.B(n_854),
.C(n_950),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1000),
.B(n_987),
.C(n_941),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_998),
.B(n_999),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1114),
.B(n_1118),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_907),
.B(n_954),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1035),
.B(n_1041),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1035),
.B(n_1041),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_977),
.B(n_1144),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1127),
.B(n_1133),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1046),
.B(n_1115),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1134),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1074),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1136),
.B(n_1145),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1024),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1078),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_913),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_841),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1160),
.B(n_1161),
.Y(n_1393)
);

NOR3xp33_ASAP7_75t_L g1394 ( 
.A(n_961),
.B(n_1062),
.C(n_879),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1082),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_980),
.B(n_996),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1163),
.B(n_1177),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1001),
.B(n_849),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_860),
.B(n_905),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1185),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1153),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1083),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1216),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1094),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1046),
.B(n_1115),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_917),
.B(n_951),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1226),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1167),
.B(n_1172),
.Y(n_1409)
);

AND2x6_ASAP7_75t_L g1410 ( 
.A(n_848),
.B(n_960),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1227),
.B(n_1229),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_916),
.A2(n_926),
.B(n_919),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1232),
.B(n_1239),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1119),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1024),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_935),
.B(n_917),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_978),
.B(n_979),
.Y(n_1417)
);

INVx4_ASAP7_75t_L g1418 ( 
.A(n_1059),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1123),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1167),
.B(n_1172),
.Y(n_1421)
);

OAI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_921),
.A2(n_932),
.B1(n_906),
.B2(n_927),
.C(n_970),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1244),
.B(n_942),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_956),
.B(n_923),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1217),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_979),
.B(n_992),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_R g1427 ( 
.A(n_1052),
.B(n_943),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1125),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1126),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1159),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_953),
.A2(n_1174),
.B1(n_1207),
.B2(n_1175),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1169),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1122),
.B(n_1157),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1217),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1210),
.B(n_914),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1180),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1210),
.B(n_1198),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_969),
.B(n_1211),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_921),
.A2(n_932),
.B1(n_952),
.B2(n_959),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1210),
.B(n_1228),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_909),
.B(n_833),
.Y(n_1443)
);

NOR3xp33_ASAP7_75t_L g1444 ( 
.A(n_961),
.B(n_1211),
.C(n_963),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_911),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_963),
.B(n_933),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1197),
.B(n_988),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_838),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_839),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_947),
.B(n_946),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_862),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_875),
.B(n_832),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_844),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_909),
.B(n_846),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1197),
.B(n_988),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_995),
.B(n_874),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_909),
.B(n_853),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_856),
.B(n_866),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_898),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_902),
.B(n_1058),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_995),
.B(n_874),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_906),
.B(n_896),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1067),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_896),
.B(n_862),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_832),
.B(n_955),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_929),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_939),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_868),
.B(n_962),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_920),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1067),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1088),
.B(n_1234),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_959),
.A2(n_993),
.B1(n_883),
.B2(n_952),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_940),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_931),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_900),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_834),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_L g1477 ( 
.A(n_993),
.B(n_958),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_915),
.B(n_958),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_993),
.A2(n_958),
.B1(n_843),
.B2(n_928),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_841),
.B(n_1064),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1050),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_874),
.B(n_1099),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1099),
.B(n_1117),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1064),
.B(n_1068),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1099),
.B(n_1117),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1117),
.B(n_1146),
.Y(n_1486)
);

NAND2xp33_ASAP7_75t_L g1487 ( 
.A(n_1146),
.B(n_1183),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_872),
.B(n_881),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1146),
.B(n_1183),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1077),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1092),
.Y(n_1492)
);

NOR3xp33_ASAP7_75t_L g1493 ( 
.A(n_981),
.B(n_1011),
.C(n_1008),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1084),
.B(n_1096),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1183),
.B(n_1240),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_868),
.B(n_962),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1087),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1104),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1128),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_872),
.B(n_881),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1096),
.B(n_1193),
.Y(n_1501)
);

AND2x2_ASAP7_75t_SL g1502 ( 
.A(n_1019),
.B(n_1007),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_885),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1150),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_L g1505 ( 
.A(n_1240),
.B(n_1137),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1165),
.B(n_1235),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1193),
.B(n_1200),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1178),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1092),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_L g1510 ( 
.A(n_1240),
.B(n_1164),
.Y(n_1510)
);

NAND2xp33_ASAP7_75t_L g1511 ( 
.A(n_1137),
.B(n_1164),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1189),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1202),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1215),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_SL g1515 ( 
.A(n_966),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1212),
.Y(n_1516)
);

INVx8_ASAP7_75t_L g1517 ( 
.A(n_1212),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_SL g1518 ( 
.A(n_966),
.Y(n_1518)
);

INVx8_ASAP7_75t_L g1519 ( 
.A(n_1023),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1194),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1194),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1200),
.B(n_1222),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1222),
.B(n_948),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_806),
.A2(n_1151),
.B(n_1149),
.C(n_1141),
.Y(n_1524)
);

NAND2xp33_ASAP7_75t_L g1525 ( 
.A(n_936),
.B(n_1121),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_948),
.B(n_1190),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_884),
.B(n_1190),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1005),
.B(n_1018),
.C(n_1017),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_813),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_884),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_957),
.B(n_910),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_957),
.B(n_910),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1106),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1106),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1124),
.B(n_1168),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1135),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_882),
.B(n_1015),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1135),
.B(n_936),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1036),
.B(n_1124),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_882),
.B(n_1238),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1080),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_986),
.A2(n_1004),
.B1(n_1009),
.B2(n_1012),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1108),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_973),
.A2(n_997),
.B(n_986),
.Y(n_1544)
);

O2A1O1Ixp5_ASAP7_75t_L g1545 ( 
.A1(n_1007),
.A2(n_1003),
.B(n_1010),
.C(n_1006),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1168),
.B(n_1171),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1191),
.B(n_1224),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1013),
.B(n_1003),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1016),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_975),
.B(n_1016),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_975),
.B(n_1016),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1014),
.B(n_1025),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_922),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1025),
.Y(n_1554)
);

BUFx5_ASAP7_75t_L g1555 ( 
.A(n_1014),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1131),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1101),
.B(n_1231),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_805),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_803),
.B(n_1029),
.Y(n_1560)
);

INVx8_ASAP7_75t_L g1561 ( 
.A(n_1100),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_803),
.A2(n_1029),
.B(n_1072),
.C(n_1049),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_803),
.B(n_1029),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_859),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_803),
.B(n_1029),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_803),
.B(n_1029),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_803),
.A2(n_1029),
.B(n_1072),
.C(n_1049),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_803),
.B(n_1029),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_805),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_803),
.B(n_1029),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_819),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_804),
.B(n_864),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_803),
.A2(n_1029),
.B(n_1072),
.C(n_1049),
.Y(n_1573)
);

NAND2xp33_ASAP7_75t_L g1574 ( 
.A(n_880),
.B(n_818),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_842),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_803),
.B(n_1029),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_842),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_859),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_859),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_803),
.B(n_1029),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_803),
.B(n_1029),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_803),
.B(n_1029),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_805),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_842),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_803),
.B(n_1029),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_803),
.B(n_1029),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_803),
.A2(n_1049),
.B1(n_1242),
.B2(n_1081),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_805),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1038),
.B(n_1045),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_803),
.B(n_1029),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_803),
.B(n_1029),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_859),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_805),
.Y(n_1597)
);

NOR2x1p5_ASAP7_75t_L g1598 ( 
.A(n_901),
.B(n_451),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_803),
.B(n_1029),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_803),
.B(n_1029),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_803),
.A2(n_1049),
.B1(n_1242),
.B2(n_1081),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_803),
.B(n_1029),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_842),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1144),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_805),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_859),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_803),
.B(n_1029),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_803),
.B(n_1029),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_803),
.B(n_1029),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_803),
.B(n_1029),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_L g1614 ( 
.A(n_880),
.B(n_818),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_803),
.B(n_1029),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_842),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1144),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1044),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_842),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_991),
.B(n_707),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_803),
.B(n_1029),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_803),
.B(n_1029),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_842),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_803),
.B(n_1029),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_803),
.B(n_1029),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_805),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_805),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_842),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_SL g1630 ( 
.A(n_990),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_803),
.B(n_1029),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_842),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1024),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_803),
.B(n_1029),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_803),
.B(n_1029),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_842),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_805),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_L g1640 ( 
.A(n_837),
.B(n_371),
.C(n_362),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_803),
.B(n_1029),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_803),
.B(n_1029),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_803),
.B(n_1029),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_803),
.B(n_1029),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_803),
.B(n_1029),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_803),
.B(n_1029),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_803),
.B(n_1029),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_803),
.B(n_1029),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_803),
.A2(n_793),
.B1(n_1049),
.B2(n_1029),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1059),
.B(n_1099),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_803),
.B(n_1029),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_803),
.B(n_1029),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_842),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1038),
.B(n_1045),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1024),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_842),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_805),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_803),
.B(n_1029),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1044),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_803),
.B(n_1029),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_803),
.B(n_1029),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_803),
.B(n_1029),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_842),
.Y(n_1667)
);

INVx8_ASAP7_75t_L g1668 ( 
.A(n_1100),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1024),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1024),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_805),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_803),
.B(n_1029),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_803),
.B(n_1029),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_803),
.B(n_1029),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_842),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_805),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_803),
.A2(n_793),
.B1(n_1049),
.B2(n_1029),
.Y(n_1677)
);

BUFx5_ASAP7_75t_L g1678 ( 
.A(n_833),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_859),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_859),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_805),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_803),
.B(n_1029),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_803),
.B(n_1029),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_803),
.A2(n_1029),
.B1(n_1072),
.B2(n_1049),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_803),
.B(n_1029),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_803),
.A2(n_1029),
.B1(n_1072),
.B2(n_1049),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_805),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_803),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_803),
.B(n_1029),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_803),
.B(n_1029),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_842),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_803),
.B(n_1029),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_803),
.B(n_1029),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_859),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_803),
.B(n_1029),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1024),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_842),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_803),
.B(n_1029),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_842),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_803),
.B(n_1029),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_805),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_803),
.B(n_1029),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_805),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_859),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_803),
.B(n_1029),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_805),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_842),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_803),
.A2(n_1029),
.B(n_1072),
.C(n_1049),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_803),
.A2(n_1029),
.B1(n_1075),
.B2(n_1072),
.C(n_1049),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_803),
.B(n_1029),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_805),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_803),
.B(n_1029),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_803),
.A2(n_1049),
.B1(n_1242),
.B2(n_1081),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_803),
.B(n_1029),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_805),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_842),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_803),
.B(n_1029),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1059),
.Y(n_1723)
);

NAND2xp33_ASAP7_75t_L g1724 ( 
.A(n_880),
.B(n_818),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_805),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1044),
.Y(n_1726)
);

A2O1A1Ixp33_ASAP7_75t_L g1727 ( 
.A1(n_803),
.A2(n_1029),
.B(n_1072),
.C(n_1049),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_819),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_805),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1086),
.B(n_493),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_803),
.B(n_1029),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_803),
.B(n_1029),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_842),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1038),
.B(n_1045),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_859),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_803),
.B(n_1029),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_803),
.B(n_1029),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1024),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1024),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_842),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_842),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_803),
.B(n_1029),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_803),
.B(n_1029),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_L g1744 ( 
.A(n_880),
.B(n_818),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_803),
.B(n_1029),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_842),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_807),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1024),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1024),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_L g1750 ( 
.A(n_880),
.B(n_818),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_805),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_803),
.B(n_1029),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_803),
.B(n_1029),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_803),
.B(n_1029),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_803),
.B(n_1029),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_803),
.B(n_1029),
.Y(n_1756)
);

BUFx5_ASAP7_75t_L g1757 ( 
.A(n_833),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_842),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_803),
.B(n_1029),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_803),
.B(n_1029),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_805),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_SL g1763 ( 
.A(n_991),
.B(n_707),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1059),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_837),
.B(n_371),
.C(n_362),
.Y(n_1765)
);

INVx8_ASAP7_75t_L g1766 ( 
.A(n_1100),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_803),
.B(n_1029),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_803),
.B(n_1029),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_L g1769 ( 
.A(n_880),
.B(n_818),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_805),
.Y(n_1770)
);

AO221x1_ASAP7_75t_L g1771 ( 
.A1(n_1116),
.A2(n_1233),
.B1(n_1205),
.B2(n_362),
.C(n_371),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_803),
.B(n_1029),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_803),
.B(n_1029),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_803),
.B(n_1029),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_803),
.B(n_1029),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_803),
.B(n_1029),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_842),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_803),
.B(n_1029),
.Y(n_1778)
);

OR2x6_ASAP7_75t_L g1779 ( 
.A(n_1024),
.B(n_1217),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_803),
.B(n_1029),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_803),
.B(n_1029),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_805),
.Y(n_1782)
);

AND2x6_ASAP7_75t_SL g1783 ( 
.A(n_967),
.B(n_972),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_SL g1784 ( 
.A(n_990),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_805),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_842),
.Y(n_1786)
);

NOR2x1p5_ASAP7_75t_L g1787 ( 
.A(n_901),
.B(n_451),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_805),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_859),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_805),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_803),
.B(n_1029),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_803),
.B(n_1029),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_803),
.B(n_1029),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_807),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1024),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_805),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_842),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_803),
.B(n_1029),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_803),
.B(n_1029),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_805),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_805),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_803),
.B(n_1029),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_803),
.B(n_1029),
.Y(n_1807)
);

BUFx3_ASAP7_75t_L g1808 ( 
.A(n_1024),
.Y(n_1808)
);

INVxp33_ASAP7_75t_L g1809 ( 
.A(n_859),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_842),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_SL g1813 ( 
.A(n_990),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_803),
.B(n_1029),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_803),
.B(n_1029),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1038),
.B(n_1045),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_803),
.B(n_1029),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_803),
.B(n_1029),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_842),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_819),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_803),
.B(n_1029),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_803),
.B(n_1029),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1024),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1059),
.B(n_1099),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_803),
.B(n_1029),
.Y(n_1827)
);

NAND2xp33_ASAP7_75t_L g1828 ( 
.A(n_880),
.B(n_818),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_805),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1044),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_803),
.B(n_1029),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_842),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_803),
.B(n_1029),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_805),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_803),
.A2(n_1049),
.B1(n_1072),
.B2(n_1029),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_805),
.Y(n_1836)
);

NAND2xp33_ASAP7_75t_SL g1837 ( 
.A(n_991),
.B(n_707),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_859),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_803),
.B(n_1029),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_803),
.B(n_1029),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_L g1841 ( 
.A(n_837),
.B(n_371),
.C(n_362),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_803),
.B(n_1029),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_803),
.B(n_1029),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1044),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_803),
.B(n_1029),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_842),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_805),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_842),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_842),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1851)
);

INVx4_ASAP7_75t_L g1852 ( 
.A(n_1059),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_803),
.B(n_1029),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_805),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_805),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_842),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_805),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_805),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_842),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1038),
.B(n_1045),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_859),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1059),
.B(n_1099),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_803),
.B(n_1029),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_842),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1024),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_803),
.B(n_1029),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_807),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_842),
.Y(n_1873)
);

NOR2xp67_ASAP7_75t_L g1874 ( 
.A(n_1059),
.B(n_1099),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_803),
.A2(n_793),
.B1(n_1049),
.B2(n_1029),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_SL g1876 ( 
.A(n_990),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_803),
.B(n_1029),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1044),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_803),
.B(n_1029),
.Y(n_1879)
);

BUFx8_ASAP7_75t_L g1880 ( 
.A(n_1023),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_805),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_842),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_803),
.B(n_1029),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_803),
.B(n_1029),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_803),
.B(n_1029),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_803),
.B(n_1029),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_803),
.B(n_1029),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_803),
.B(n_1029),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_803),
.B(n_1029),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_803),
.B(n_1029),
.Y(n_1892)
);

NOR2xp67_ASAP7_75t_SL g1893 ( 
.A(n_1059),
.B(n_1099),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_803),
.B(n_1029),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_803),
.B(n_1029),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_803),
.A2(n_793),
.B1(n_1049),
.B2(n_1029),
.Y(n_1898)
);

OAI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_803),
.A2(n_1049),
.B1(n_1072),
.B2(n_1029),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_859),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_803),
.B(n_1029),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_805),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1024),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1116),
.B(n_1233),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_803),
.B(n_1029),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_859),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_803),
.B(n_1029),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1268),
.Y(n_1908)
);

NAND2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1336),
.B(n_1392),
.Y(n_1909)
);

AO22x2_ASAP7_75t_L g1910 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_1910)
);

AO22x2_ASAP7_75t_L g1911 ( 
.A1(n_1588),
.A2(n_1593),
.B1(n_1601),
.B2(n_1590),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1260),
.B(n_1381),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1246),
.B(n_1595),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1324),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1270),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1560),
.B(n_1565),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1287),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1712),
.A2(n_1687),
.B1(n_1685),
.B2(n_1576),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1289),
.Y(n_1919)
);

AO22x2_ASAP7_75t_L g1920 ( 
.A1(n_1608),
.A2(n_1617),
.B1(n_1633),
.B2(n_1612),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1291),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1300),
.Y(n_1922)
);

AND2x2_ASAP7_75t_SL g1923 ( 
.A(n_1255),
.B(n_1586),
.Y(n_1923)
);

NAND2x1p5_ASAP7_75t_L g1924 ( 
.A(n_1392),
.B(n_1350),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1300),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1611),
.B(n_1622),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1564),
.B(n_1578),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1257),
.B(n_1835),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1292),
.Y(n_1929)
);

AO22x2_ASAP7_75t_L g1930 ( 
.A1(n_1635),
.A2(n_1646),
.B1(n_1666),
.B2(n_1663),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1296),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1650),
.A2(n_1898),
.B1(n_1875),
.B2(n_1677),
.C(n_1640),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1300),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1304),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1355),
.Y(n_1935)
);

AO22x2_ASAP7_75t_L g1936 ( 
.A1(n_1679),
.A2(n_1701),
.B1(n_1719),
.B2(n_1707),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1300),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1615),
.B(n_1731),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1313),
.Y(n_1939)
);

NOR2xp67_ASAP7_75t_L g1940 ( 
.A(n_1580),
.B(n_1596),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1374),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1322),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1323),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1300),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1625),
.A2(n_1637),
.B1(n_1644),
.B2(n_1626),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1899),
.B(n_1265),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1348),
.Y(n_1947)
);

OR2x6_ASAP7_75t_L g1948 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1301),
.Y(n_1949)
);

OAI221xp5_ASAP7_75t_L g1950 ( 
.A1(n_1765),
.A2(n_1841),
.B1(n_1716),
.B2(n_1602),
.C(n_1589),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1672),
.B(n_1674),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1332),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1683),
.B(n_1686),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1263),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1693),
.B(n_1761),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1737),
.B(n_1753),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1780),
.A2(n_1806),
.B1(n_1807),
.B2(n_1801),
.C(n_1795),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1267),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1886),
.B(n_1888),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1575),
.Y(n_1960)
);

AO22x2_ASAP7_75t_L g1961 ( 
.A1(n_1720),
.A2(n_1788),
.B1(n_1789),
.B2(n_1758),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1754),
.B(n_1774),
.Y(n_1962)
);

OAI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1890),
.A2(n_1905),
.B1(n_1562),
.B2(n_1727),
.C(n_1567),
.Y(n_1963)
);

OR2x6_ASAP7_75t_SL g1964 ( 
.A(n_1310),
.B(n_1664),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1577),
.Y(n_1965)
);

BUFx8_ASAP7_75t_L g1966 ( 
.A(n_1515),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_SL g1967 ( 
.A(n_1779),
.Y(n_1967)
);

AO22x2_ASAP7_75t_L g1968 ( 
.A1(n_1802),
.A2(n_1810),
.B1(n_1812),
.B2(n_1803),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1585),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1273),
.B(n_1269),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1605),
.Y(n_1971)
);

AO22x2_ASAP7_75t_L g1972 ( 
.A1(n_1818),
.A2(n_1851),
.B1(n_1853),
.B2(n_1826),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1604),
.Y(n_1973)
);

AO22x2_ASAP7_75t_L g1974 ( 
.A1(n_1856),
.A2(n_1858),
.B1(n_1864),
.B2(n_1857),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1616),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1620),
.Y(n_1976)
);

AO22x2_ASAP7_75t_L g1977 ( 
.A1(n_1887),
.A2(n_1897),
.B1(n_1894),
.B2(n_1314),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1624),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1629),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1359),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1632),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1638),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1563),
.A2(n_1566),
.B1(n_1581),
.B2(n_1570),
.C(n_1568),
.Y(n_1983)
);

CKINVDCx16_ASAP7_75t_R g1984 ( 
.A(n_1730),
.Y(n_1984)
);

NAND2x1p5_ASAP7_75t_L g1985 ( 
.A(n_1893),
.B(n_1275),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1654),
.Y(n_1986)
);

OR2x6_ASAP7_75t_L g1987 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1987)
);

OAI21xp33_ASAP7_75t_L g1988 ( 
.A1(n_1582),
.A2(n_1587),
.B(n_1583),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1618),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1657),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1827),
.B(n_1833),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1667),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1675),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1253),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1692),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1503),
.Y(n_1996)
);

AO22x2_ASAP7_75t_L g1997 ( 
.A1(n_1847),
.A2(n_1885),
.B1(n_1259),
.B2(n_1256),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1383),
.Y(n_1998)
);

BUFx8_ASAP7_75t_L g1999 ( 
.A(n_1515),
.Y(n_1999)
);

BUFx8_ASAP7_75t_L g2000 ( 
.A(n_1518),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1698),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1700),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1845),
.B(n_1258),
.Y(n_2004)
);

AO22x2_ASAP7_75t_L g2005 ( 
.A1(n_1254),
.A2(n_1599),
.B1(n_1600),
.B2(n_1594),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1710),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1603),
.B(n_1609),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1721),
.Y(n_2008)
);

CKINVDCx20_ASAP7_75t_R g2009 ( 
.A(n_1880),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1315),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1396),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1733),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1740),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1779),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1741),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1610),
.B(n_1613),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1746),
.Y(n_2017)
);

AO22x2_ASAP7_75t_L g2018 ( 
.A1(n_1623),
.A2(n_1636),
.B1(n_1641),
.B2(n_1631),
.Y(n_2018)
);

OAI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_1642),
.A2(n_1647),
.B1(n_1648),
.B2(n_1645),
.C(n_1643),
.Y(n_2019)
);

OAI221xp5_ASAP7_75t_L g2020 ( 
.A1(n_1649),
.A2(n_1659),
.B1(n_1661),
.B2(n_1653),
.C(n_1652),
.Y(n_2020)
);

OA22x2_ASAP7_75t_L g2021 ( 
.A1(n_1662),
.A2(n_1673),
.B1(n_1684),
.B2(n_1665),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1759),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1278),
.A2(n_1346),
.B1(n_1378),
.B2(n_1345),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1266),
.Y(n_2024)
);

AO22x2_ASAP7_75t_L g2025 ( 
.A1(n_1690),
.A2(n_1694),
.B1(n_1696),
.B2(n_1691),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_SL g2026 ( 
.A1(n_1247),
.A2(n_1250),
.B1(n_1702),
.B2(n_1699),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1573),
.A2(n_1711),
.B1(n_1699),
.B2(n_1702),
.C(n_1247),
.Y(n_2027)
);

INVxp67_ASAP7_75t_L g2028 ( 
.A(n_1747),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1347),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1777),
.Y(n_2030)
);

AND2x6_ASAP7_75t_L g2031 ( 
.A(n_1326),
.B(n_1327),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1264),
.B(n_1250),
.Y(n_2032)
);

AO22x2_ASAP7_75t_L g2033 ( 
.A1(n_1704),
.A2(n_1708),
.B1(n_1715),
.B2(n_1713),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1704),
.B(n_1708),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1786),
.Y(n_2035)
);

OAI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1713),
.A2(n_1715),
.B1(n_1732),
.B2(n_1722),
.C(n_1717),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1678),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1717),
.A2(n_1722),
.B1(n_1742),
.B2(n_1736),
.C(n_1732),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_1275),
.Y(n_2039)
);

AO22x2_ASAP7_75t_L g2040 ( 
.A1(n_1736),
.A2(n_1742),
.B1(n_1745),
.B2(n_1743),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1391),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1743),
.A2(n_1752),
.B1(n_1755),
.B2(n_1745),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1271),
.B(n_1272),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1799),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1811),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1820),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1302),
.B(n_1303),
.Y(n_2047)
);

NOR2x1p5_ASAP7_75t_L g2048 ( 
.A(n_1492),
.B(n_1748),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1271),
.B(n_1272),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1382),
.B(n_1406),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1832),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1253),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1846),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_1880),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1849),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1850),
.Y(n_2056)
);

AO22x2_ASAP7_75t_L g2057 ( 
.A1(n_1752),
.A2(n_1756),
.B1(n_1760),
.B2(n_1755),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1860),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1275),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1863),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1869),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_1796),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1274),
.B(n_1281),
.Y(n_2063)
);

AO22x2_ASAP7_75t_L g2064 ( 
.A1(n_1756),
.A2(n_1767),
.B1(n_1768),
.B2(n_1760),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1873),
.Y(n_2065)
);

AO22x2_ASAP7_75t_L g2066 ( 
.A1(n_1767),
.A2(n_1772),
.B1(n_1773),
.B2(n_1768),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1772),
.B(n_1773),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1882),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_1872),
.Y(n_2069)
);

OAI21xp33_ASAP7_75t_L g2070 ( 
.A1(n_1775),
.A2(n_1778),
.B(n_1776),
.Y(n_2070)
);

AO22x2_ASAP7_75t_L g2071 ( 
.A1(n_1775),
.A2(n_1778),
.B1(n_1781),
.B2(n_1776),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1423),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1365),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1779),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_SL g2075 ( 
.A(n_1556),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1366),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1369),
.Y(n_2077)
);

AO22x2_ASAP7_75t_L g2078 ( 
.A1(n_1781),
.A2(n_1794),
.B1(n_1800),
.B2(n_1793),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1793),
.B(n_1794),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1371),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1274),
.B(n_1281),
.Y(n_2081)
);

BUFx8_ASAP7_75t_L g2082 ( 
.A(n_1518),
.Y(n_2082)
);

AO22x2_ASAP7_75t_L g2083 ( 
.A1(n_1907),
.A2(n_1800),
.B1(n_1815),
.B2(n_1814),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1372),
.Y(n_2084)
);

AO22x2_ASAP7_75t_L g2085 ( 
.A1(n_1907),
.A2(n_1814),
.B1(n_1817),
.B2(n_1815),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1817),
.B(n_1819),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1373),
.Y(n_2087)
);

OAI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_1819),
.A2(n_1831),
.B1(n_1839),
.B2(n_1823),
.C(n_1822),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1678),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1379),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1245),
.Y(n_2091)
);

AO22x2_ASAP7_75t_L g2092 ( 
.A1(n_1822),
.A2(n_1823),
.B1(n_1839),
.B2(n_1831),
.Y(n_2092)
);

AO22x2_ASAP7_75t_L g2093 ( 
.A1(n_1840),
.A2(n_1842),
.B1(n_1854),
.B2(n_1843),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1382),
.B(n_1406),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1678),
.Y(n_2095)
);

BUFx8_ASAP7_75t_L g2096 ( 
.A(n_1556),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1384),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1840),
.B(n_1842),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1678),
.Y(n_2099)
);

AO22x2_ASAP7_75t_L g2100 ( 
.A1(n_1843),
.A2(n_1854),
.B1(n_1871),
.B2(n_1868),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1388),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1393),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1397),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1572),
.B(n_1530),
.Y(n_2104)
);

AO22x2_ASAP7_75t_L g2105 ( 
.A1(n_1868),
.A2(n_1871),
.B1(n_1879),
.B2(n_1877),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1402),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1286),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1877),
.B(n_1879),
.Y(n_2108)
);

BUFx8_ASAP7_75t_L g2109 ( 
.A(n_1556),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1298),
.B(n_1337),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1411),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_1398),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1413),
.Y(n_2113)
);

OAI22xp33_ASAP7_75t_SL g2114 ( 
.A1(n_1883),
.A2(n_1884),
.B1(n_1891),
.B2(n_1889),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1757),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1282),
.B(n_1592),
.Y(n_2116)
);

AO22x2_ASAP7_75t_L g2117 ( 
.A1(n_1883),
.A2(n_1884),
.B1(n_1891),
.B2(n_1889),
.Y(n_2117)
);

AO22x2_ASAP7_75t_L g2118 ( 
.A1(n_1892),
.A2(n_1895),
.B1(n_1901),
.B2(n_1896),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1419),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1356),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1892),
.B(n_1895),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1364),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1370),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_1446),
.Y(n_2124)
);

BUFx8_ASAP7_75t_L g2125 ( 
.A(n_1630),
.Y(n_2125)
);

OAI21xp33_ASAP7_75t_L g2126 ( 
.A1(n_1896),
.A2(n_1901),
.B(n_1282),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_1572),
.B(n_1533),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1386),
.Y(n_2128)
);

NAND2x1p5_ASAP7_75t_L g2129 ( 
.A(n_1325),
.B(n_1844),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1400),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1655),
.B(n_1734),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_1401),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1404),
.Y(n_2133)
);

OAI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_1307),
.A2(n_1362),
.B1(n_1865),
.B2(n_1816),
.C(n_1689),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1534),
.B(n_1536),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1283),
.B(n_1293),
.Y(n_2136)
);

INVxp67_ASAP7_75t_L g2137 ( 
.A(n_1368),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1408),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1445),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1253),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1458),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1305),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1757),
.Y(n_2143)
);

AO22x2_ASAP7_75t_L g2144 ( 
.A1(n_1771),
.A2(n_1279),
.B1(n_1444),
.B2(n_1394),
.Y(n_2144)
);

AO22x2_ASAP7_75t_L g2145 ( 
.A1(n_1437),
.A2(n_1298),
.B1(n_1327),
.B2(n_1326),
.Y(n_2145)
);

INVxp67_ASAP7_75t_L g2146 ( 
.A(n_1537),
.Y(n_2146)
);

OAI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_1376),
.A2(n_1493),
.B1(n_1528),
.B2(n_1377),
.C(n_1299),
.Y(n_2147)
);

AO22x1_ASAP7_75t_L g2148 ( 
.A1(n_1809),
.A2(n_1407),
.B1(n_1417),
.B2(n_1316),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1458),
.Y(n_2149)
);

NAND2x1p5_ASAP7_75t_L g2150 ( 
.A(n_1325),
.B(n_1844),
.Y(n_2150)
);

NAND2x1p5_ASAP7_75t_L g2151 ( 
.A(n_1325),
.B(n_1844),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_1509),
.Y(n_2152)
);

AO22x2_ASAP7_75t_L g2153 ( 
.A1(n_1437),
.A2(n_1335),
.B1(n_1431),
.B2(n_1328),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1294),
.B(n_1309),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_1276),
.Y(n_2155)
);

OAI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_1277),
.A2(n_1306),
.B1(n_1303),
.B2(n_1302),
.C(n_1339),
.Y(n_2156)
);

AO22x2_ASAP7_75t_L g2157 ( 
.A1(n_1328),
.A2(n_1335),
.B1(n_1434),
.B2(n_1431),
.Y(n_2157)
);

OAI221xp5_ASAP7_75t_L g2158 ( 
.A1(n_1306),
.A2(n_1542),
.B1(n_1309),
.B2(n_1331),
.C(n_1341),
.Y(n_2158)
);

INVxp67_ASAP7_75t_L g2159 ( 
.A(n_1509),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1424),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1450),
.B(n_1334),
.Y(n_2161)
);

AO22x2_ASAP7_75t_L g2162 ( 
.A1(n_1434),
.A2(n_1435),
.B1(n_1321),
.B2(n_1478),
.Y(n_2162)
);

AO22x2_ASAP7_75t_L g2163 ( 
.A1(n_1435),
.A2(n_1478),
.B1(n_1442),
.B2(n_1439),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1472),
.B(n_1464),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_1462),
.B(n_1527),
.Y(n_2165)
);

OAI221xp5_ASAP7_75t_L g2166 ( 
.A1(n_1344),
.A2(n_1311),
.B1(n_1680),
.B2(n_1681),
.C(n_1607),
.Y(n_2166)
);

AO22x2_ASAP7_75t_L g2167 ( 
.A1(n_1439),
.A2(n_1442),
.B1(n_1320),
.B2(n_1329),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1449),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1453),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1757),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1757),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1527),
.B(n_1526),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1353),
.B(n_1479),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_1399),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1469),
.B(n_1474),
.Y(n_2175)
);

CKINVDCx16_ASAP7_75t_R g2176 ( 
.A(n_1427),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1249),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1797),
.Y(n_2178)
);

NAND2x1p5_ASAP7_75t_L g2179 ( 
.A(n_1878),
.B(n_1544),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1251),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1695),
.B(n_1706),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1261),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1454),
.B(n_1457),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1280),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_L g2185 ( 
.A(n_1545),
.B(n_1906),
.C(n_1791),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1284),
.Y(n_2186)
);

AOI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_1380),
.A2(n_1735),
.B1(n_1866),
.B2(n_1838),
.Y(n_2187)
);

AO22x2_ASAP7_75t_L g2188 ( 
.A1(n_1351),
.A2(n_1443),
.B1(n_1475),
.B2(n_1900),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1288),
.Y(n_2189)
);

BUFx8_ASAP7_75t_L g2190 ( 
.A(n_1630),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1330),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_1540),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1509),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1757),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1295),
.Y(n_2195)
);

AO22x2_ASAP7_75t_L g2196 ( 
.A1(n_1443),
.A2(n_1454),
.B1(n_1457),
.B2(n_1363),
.Y(n_2196)
);

CKINVDCx20_ASAP7_75t_R g2197 ( 
.A(n_1571),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1358),
.B(n_1432),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1333),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1757),
.Y(n_2200)
);

AOI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1502),
.A2(n_1308),
.B1(n_1426),
.B2(n_1440),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_1516),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1412),
.B(n_1465),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1340),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1441),
.B(n_1555),
.Y(n_2205)
);

CKINVDCx20_ASAP7_75t_R g2206 ( 
.A(n_1728),
.Y(n_2206)
);

OAI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_1422),
.A2(n_1338),
.B1(n_1455),
.B2(n_1447),
.C(n_1367),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1342),
.Y(n_2208)
);

AO22x2_ASAP7_75t_L g2209 ( 
.A1(n_1552),
.A2(n_1460),
.B1(n_1554),
.B2(n_1482),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1471),
.A2(n_1361),
.B1(n_1460),
.B2(n_1354),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1357),
.Y(n_2211)
);

AO22x2_ASAP7_75t_L g2212 ( 
.A1(n_1471),
.A2(n_1375),
.B1(n_1390),
.B2(n_1387),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_1276),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1395),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1403),
.Y(n_2215)
);

AO22x2_ASAP7_75t_L g2216 ( 
.A1(n_1405),
.A2(n_1703),
.B1(n_1705),
.B2(n_1902),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1448),
.B(n_1459),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1555),
.B(n_1414),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1420),
.Y(n_2219)
);

AND2x2_ASAP7_75t_SL g2220 ( 
.A(n_1544),
.B(n_1312),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_1276),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1428),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1429),
.Y(n_2223)
);

NAND2x1p5_ASAP7_75t_L g2224 ( 
.A(n_1878),
.B(n_1262),
.Y(n_2224)
);

INVx4_ASAP7_75t_L g2225 ( 
.A(n_1878),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1430),
.Y(n_2226)
);

BUFx8_ASAP7_75t_L g2227 ( 
.A(n_1784),
.Y(n_2227)
);

AO22x2_ASAP7_75t_L g2228 ( 
.A1(n_1433),
.A2(n_1792),
.B1(n_1658),
.B2(n_1628),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_1385),
.A2(n_1409),
.B1(n_1421),
.B2(n_1763),
.C(n_1621),
.Y(n_2229)
);

BUFx2_ASAP7_75t_L g2230 ( 
.A(n_1540),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1526),
.B(n_1549),
.Y(n_2231)
);

BUFx8_ASAP7_75t_L g2232 ( 
.A(n_1784),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1438),
.Y(n_2233)
);

CKINVDCx20_ASAP7_75t_R g2234 ( 
.A(n_1821),
.Y(n_2234)
);

AO22x2_ASAP7_75t_L g2235 ( 
.A1(n_1559),
.A2(n_1639),
.B1(n_1627),
.B2(n_1606),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1569),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1813),
.Y(n_2237)
);

AO22x2_ASAP7_75t_L g2238 ( 
.A1(n_1584),
.A2(n_1798),
.B1(n_1671),
.B2(n_1597),
.Y(n_2238)
);

CKINVDCx16_ASAP7_75t_R g2239 ( 
.A(n_1813),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1555),
.B(n_1591),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1676),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1682),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1688),
.B(n_1709),
.Y(n_2243)
);

OAI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_1837),
.A2(n_1548),
.B1(n_1551),
.B2(n_1550),
.C(n_1352),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1714),
.B(n_1718),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1725),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1729),
.B(n_1751),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1555),
.B(n_1762),
.Y(n_2248)
);

BUFx8_ASAP7_75t_L g2249 ( 
.A(n_1876),
.Y(n_2249)
);

AOI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_1876),
.A2(n_1416),
.B1(n_1468),
.B2(n_1496),
.Y(n_2250)
);

NAND2x1p5_ASAP7_75t_L g2251 ( 
.A(n_1262),
.B(n_1290),
.Y(n_2251)
);

BUFx8_ASAP7_75t_L g2252 ( 
.A(n_1516),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1770),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1782),
.B(n_1785),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1549),
.B(n_1790),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1804),
.Y(n_2256)
);

NAND2x1p5_ASAP7_75t_L g2257 ( 
.A(n_1290),
.B(n_1418),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1805),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1829),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1834),
.B(n_1836),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1555),
.B(n_1848),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1855),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_1540),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1859),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1861),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1862),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1466),
.B(n_1467),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_1555),
.B(n_1881),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1473),
.B(n_1488),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1538),
.B(n_1531),
.Y(n_2270)
);

NAND2x1p5_ASAP7_75t_L g2271 ( 
.A(n_1418),
.B(n_1723),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_1516),
.Y(n_2272)
);

INVxp67_ASAP7_75t_SL g2273 ( 
.A(n_1480),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1476),
.Y(n_2274)
);

AO22x2_ASAP7_75t_L g2275 ( 
.A1(n_1535),
.A2(n_1456),
.B1(n_1461),
.B2(n_1521),
.Y(n_2275)
);

AO22x2_ASAP7_75t_L g2276 ( 
.A1(n_1349),
.A2(n_1498),
.B1(n_1481),
.B2(n_1491),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_1410),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_1561),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1504),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1497),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1499),
.Y(n_2281)
);

OAI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_1553),
.A2(n_1343),
.B1(n_1451),
.B2(n_1524),
.C(n_1539),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1519),
.Y(n_2283)
);

OAI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_1525),
.A2(n_1529),
.B1(n_1543),
.B2(n_1470),
.C(n_1463),
.Y(n_2284)
);

AO22x2_ASAP7_75t_L g2285 ( 
.A1(n_1508),
.A2(n_1513),
.B1(n_1514),
.B2(n_1512),
.Y(n_2285)
);

INVxp67_ASAP7_75t_L g2286 ( 
.A(n_1511),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_1252),
.A2(n_1769),
.B1(n_1614),
.B2(n_1744),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1360),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1506),
.B(n_1452),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_1561),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1520),
.Y(n_2291)
);

OAI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_1574),
.A2(n_1828),
.B1(n_1724),
.B2(n_1750),
.C(n_1505),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1285),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_1532),
.B(n_1285),
.Y(n_2294)
);

INVxp67_ASAP7_75t_L g2295 ( 
.A(n_1547),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_1723),
.B(n_1764),
.Y(n_2296)
);

NAND2x1p5_ASAP7_75t_L g2297 ( 
.A(n_1764),
.B(n_1852),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_1808),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_1317),
.B(n_1830),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1317),
.Y(n_2300)
);

NAND3xp33_ASAP7_75t_SL g2301 ( 
.A(n_1546),
.B(n_1541),
.C(n_1483),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1500),
.B(n_1830),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1619),
.Y(n_2303)
);

OA22x2_ASAP7_75t_L g2304 ( 
.A1(n_1485),
.A2(n_1495),
.B1(n_1490),
.B2(n_1486),
.Y(n_2304)
);

CKINVDCx11_ASAP7_75t_R g2305 ( 
.A(n_1519),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1619),
.B(n_1726),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_SL g2307 ( 
.A1(n_1557),
.A2(n_1852),
.B1(n_1523),
.B2(n_1507),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1519),
.Y(n_2308)
);

NOR2xp67_ASAP7_75t_L g2309 ( 
.A(n_1651),
.B(n_1874),
.Y(n_2309)
);

AO22x2_ASAP7_75t_L g2310 ( 
.A1(n_1660),
.A2(n_1726),
.B1(n_1410),
.B2(n_1522),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1480),
.B(n_1484),
.Y(n_2311)
);

AO22x2_ASAP7_75t_L g2312 ( 
.A1(n_1660),
.A2(n_1410),
.B1(n_1523),
.B2(n_1489),
.Y(n_2312)
);

NAND2x1p5_ASAP7_75t_L g2313 ( 
.A(n_1825),
.B(n_1867),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1410),
.Y(n_2314)
);

OAI221xp5_ASAP7_75t_L g2315 ( 
.A1(n_1510),
.A2(n_1487),
.B1(n_1477),
.B2(n_1870),
.C(n_1415),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1484),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1489),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1494),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1494),
.Y(n_2319)
);

CKINVDCx14_ASAP7_75t_R g2320 ( 
.A(n_1561),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1501),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1501),
.Y(n_2322)
);

HB1xp67_ASAP7_75t_L g2323 ( 
.A(n_1668),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_1598),
.B(n_1787),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1410),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1507),
.B(n_1766),
.Y(n_2326)
);

AND2x4_ASAP7_75t_L g2327 ( 
.A(n_1389),
.B(n_1670),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1668),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_1668),
.B(n_1766),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1297),
.B(n_1783),
.Y(n_2330)
);

NAND2x1p5_ASAP7_75t_L g2331 ( 
.A(n_1425),
.B(n_1436),
.Y(n_2331)
);

AO22x2_ASAP7_75t_L g2332 ( 
.A1(n_1634),
.A2(n_1739),
.B1(n_1656),
.B2(n_1669),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1766),
.Y(n_2333)
);

OAI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_1697),
.A2(n_1738),
.B1(n_1749),
.B2(n_1824),
.C(n_1903),
.Y(n_2334)
);

AO22x2_ASAP7_75t_L g2335 ( 
.A1(n_1517),
.A2(n_1687),
.B1(n_1685),
.B2(n_1558),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1517),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_1517),
.B(n_1260),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_1355),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_L g2340 ( 
.A(n_1562),
.B(n_1567),
.Y(n_2340)
);

AO22x2_ASAP7_75t_L g2341 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1268),
.Y(n_2342)
);

AO22x2_ASAP7_75t_L g2343 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2344)
);

OAI221xp5_ASAP7_75t_L g2345 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2345)
);

AO22x2_ASAP7_75t_L g2346 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1268),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2348)
);

OAI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2349)
);

AO22x2_ASAP7_75t_L g2350 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1560),
.B(n_803),
.Y(n_2351)
);

OR2x6_ASAP7_75t_L g2352 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1560),
.B(n_803),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1268),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1268),
.Y(n_2355)
);

AO22x2_ASAP7_75t_L g2356 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_1359),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1560),
.B(n_803),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1268),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1560),
.B(n_803),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1268),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1560),
.B(n_803),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1560),
.B(n_803),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1560),
.B(n_803),
.Y(n_2365)
);

AO22x2_ASAP7_75t_L g2366 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1268),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1300),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1268),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1300),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1300),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_1336),
.Y(n_2372)
);

AO22x2_ASAP7_75t_L g2373 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1268),
.Y(n_2374)
);

AND2x6_ASAP7_75t_L g2375 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1268),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_1374),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1268),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1268),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1300),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_SL g2382 ( 
.A(n_1779),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2383)
);

NAND2x1p5_ASAP7_75t_L g2384 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1300),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1268),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_1374),
.Y(n_2387)
);

AO22x2_ASAP7_75t_L g2388 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1268),
.Y(n_2389)
);

AO22x2_ASAP7_75t_L g2390 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2390)
);

AO22x2_ASAP7_75t_L g2391 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1300),
.Y(n_2392)
);

AO22x2_ASAP7_75t_L g2393 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1560),
.B(n_803),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1268),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1268),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_1355),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1268),
.Y(n_2398)
);

AO22x2_ASAP7_75t_L g2399 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1560),
.B(n_803),
.Y(n_2400)
);

BUFx8_ASAP7_75t_L g2401 ( 
.A(n_1515),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1268),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_1273),
.B(n_1269),
.Y(n_2404)
);

NAND2x1p5_ASAP7_75t_L g2405 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_1391),
.Y(n_2406)
);

OAI221xp5_ASAP7_75t_L g2407 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1268),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_1779),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1268),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1268),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1268),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1268),
.Y(n_2415)
);

AO22x2_ASAP7_75t_L g2416 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1268),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1560),
.B(n_803),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1268),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2421)
);

INVxp67_ASAP7_75t_SL g2422 ( 
.A(n_1347),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1268),
.Y(n_2423)
);

AND2x6_ASAP7_75t_L g2424 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2424)
);

NOR2xp67_ASAP7_75t_L g2425 ( 
.A(n_1564),
.B(n_941),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1268),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2427)
);

NAND2x1p5_ASAP7_75t_L g2428 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1268),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1268),
.Y(n_2430)
);

OAI221xp5_ASAP7_75t_L g2431 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_1300),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_1300),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1268),
.Y(n_2434)
);

NAND2x1p5_ASAP7_75t_L g2435 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1268),
.Y(n_2436)
);

INVxp67_ASAP7_75t_SL g2437 ( 
.A(n_1347),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1268),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_1324),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1268),
.Y(n_2440)
);

INVxp67_ASAP7_75t_L g2441 ( 
.A(n_1355),
.Y(n_2441)
);

INVx2_ASAP7_75t_SL g2442 ( 
.A(n_1374),
.Y(n_2442)
);

AO22x2_ASAP7_75t_L g2443 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2443)
);

OAI221xp5_ASAP7_75t_L g2444 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2444)
);

AOI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_1336),
.Y(n_2446)
);

NAND2x1p5_ASAP7_75t_L g2447 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1268),
.Y(n_2448)
);

INVxp67_ASAP7_75t_L g2449 ( 
.A(n_1355),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1268),
.Y(n_2450)
);

OAI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_1391),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_1560),
.B(n_803),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1268),
.Y(n_2455)
);

OAI221xp5_ASAP7_75t_L g2456 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2456)
);

NOR2xp67_ASAP7_75t_L g2457 ( 
.A(n_1564),
.B(n_941),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2458)
);

NAND2x1p5_ASAP7_75t_L g2459 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1560),
.B(n_803),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1268),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1268),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_1268),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1268),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1268),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1560),
.B(n_803),
.Y(n_2468)
);

NAND2x1p5_ASAP7_75t_L g2469 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_1300),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_1268),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_1560),
.B(n_803),
.Y(n_2472)
);

AND2x2_ASAP7_75t_SL g2473 ( 
.A(n_1255),
.B(n_803),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_1268),
.Y(n_2474)
);

AO22x2_ASAP7_75t_L g2475 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2475)
);

OAI221xp5_ASAP7_75t_L g2476 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1560),
.B(n_803),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_1355),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_1268),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_1268),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2481)
);

OAI22xp33_ASAP7_75t_SL g2482 ( 
.A1(n_1712),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2482)
);

INVxp67_ASAP7_75t_L g2483 ( 
.A(n_1355),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_1355),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_1300),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1268),
.Y(n_2487)
);

AO22x2_ASAP7_75t_L g2488 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2488)
);

NOR2xp67_ASAP7_75t_L g2489 ( 
.A(n_1564),
.B(n_941),
.Y(n_2489)
);

NAND2xp33_ASAP7_75t_L g2490 ( 
.A(n_1562),
.B(n_1567),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_1268),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1268),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_1273),
.B(n_1269),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_1268),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_1300),
.Y(n_2496)
);

NAND2x1p5_ASAP7_75t_L g2497 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2497)
);

NAND2x1p5_ASAP7_75t_L g2498 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1268),
.Y(n_2500)
);

NAND2x1p5_ASAP7_75t_L g2501 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2501)
);

AO22x2_ASAP7_75t_L g2502 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_SL g2503 ( 
.A(n_1779),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1268),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_1268),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1268),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1560),
.B(n_803),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1560),
.B(n_803),
.Y(n_2508)
);

CKINVDCx11_ASAP7_75t_R g2509 ( 
.A(n_1503),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_1268),
.Y(n_2510)
);

OAI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_1650),
.A2(n_803),
.B1(n_1049),
.B2(n_1029),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1268),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1268),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1268),
.Y(n_2515)
);

OAI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_1268),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_1560),
.B(n_803),
.Y(n_2518)
);

OAI221xp5_ASAP7_75t_L g2519 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1268),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_1268),
.Y(n_2522)
);

NAND2x1p5_ASAP7_75t_L g2523 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2523)
);

AO22x2_ASAP7_75t_L g2524 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2524)
);

INVxp67_ASAP7_75t_L g2525 ( 
.A(n_1355),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1300),
.Y(n_2526)
);

AO22x2_ASAP7_75t_L g2527 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_1560),
.B(n_803),
.Y(n_2529)
);

INVxp33_ASAP7_75t_L g2530 ( 
.A(n_1355),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_1300),
.Y(n_2531)
);

INVx1_ASAP7_75t_SL g2532 ( 
.A(n_1324),
.Y(n_2532)
);

NAND2x1p5_ASAP7_75t_L g2533 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2533)
);

AO22x2_ASAP7_75t_L g2534 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1268),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_1336),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_1268),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_1268),
.Y(n_2538)
);

AO22x2_ASAP7_75t_L g2539 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1268),
.Y(n_2540)
);

INVx3_ASAP7_75t_L g2541 ( 
.A(n_1336),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_1268),
.Y(n_2542)
);

AO22x2_ASAP7_75t_L g2543 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_1300),
.Y(n_2544)
);

NAND2x1p5_ASAP7_75t_L g2545 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2545)
);

AO22x2_ASAP7_75t_L g2546 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_1268),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_1300),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2549)
);

AO22x2_ASAP7_75t_L g2550 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_1268),
.Y(n_2551)
);

AO22x2_ASAP7_75t_L g2552 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_1359),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_1300),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1391),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1268),
.Y(n_2556)
);

XNOR2x2_ASAP7_75t_SL g2557 ( 
.A(n_1310),
.B(n_1589),
.Y(n_2557)
);

AO22x2_ASAP7_75t_L g2558 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_1300),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_1268),
.Y(n_2560)
);

CKINVDCx20_ASAP7_75t_R g2561 ( 
.A(n_1503),
.Y(n_2561)
);

AO22x2_ASAP7_75t_L g2562 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_1324),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1300),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_1268),
.Y(n_2565)
);

AOI22xp33_ASAP7_75t_L g2566 ( 
.A1(n_1712),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_1268),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_1779),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_1268),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1268),
.Y(n_2571)
);

INVxp67_ASAP7_75t_L g2572 ( 
.A(n_1355),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_1300),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_1268),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_1391),
.Y(n_2575)
);

NOR2x1p5_ASAP7_75t_L g2576 ( 
.A(n_1492),
.B(n_451),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_1268),
.Y(n_2577)
);

NAND2x1p5_ASAP7_75t_L g2578 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2578)
);

NAND2x1p5_ASAP7_75t_L g2579 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_1268),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1268),
.Y(n_2581)
);

AO22x2_ASAP7_75t_L g2582 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1268),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1268),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_1268),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_1268),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_1268),
.Y(n_2589)
);

INVxp67_ASAP7_75t_L g2590 ( 
.A(n_1355),
.Y(n_2590)
);

AO22x2_ASAP7_75t_L g2591 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_1268),
.Y(n_2592)
);

BUFx8_ASAP7_75t_L g2593 ( 
.A(n_1515),
.Y(n_2593)
);

AO22x2_ASAP7_75t_L g2594 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_1268),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_1300),
.Y(n_2596)
);

OAI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_1589),
.A2(n_1716),
.B1(n_1602),
.B2(n_1029),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_1268),
.Y(n_2598)
);

OR2x6_ASAP7_75t_L g2599 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_1268),
.Y(n_2600)
);

AO22x2_ASAP7_75t_L g2601 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2601)
);

AO22x2_ASAP7_75t_L g2602 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2602)
);

AO22x2_ASAP7_75t_L g2603 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2603)
);

BUFx2_ASAP7_75t_L g2604 ( 
.A(n_1359),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_1560),
.B(n_803),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_1268),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_1560),
.B(n_803),
.Y(n_2607)
);

AO22x2_ASAP7_75t_L g2608 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_1560),
.B(n_803),
.Y(n_2609)
);

AOI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1268),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1268),
.Y(n_2612)
);

NAND2x1p5_ASAP7_75t_L g2613 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_1560),
.B(n_803),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_1268),
.Y(n_2615)
);

NOR2xp67_ASAP7_75t_L g2616 ( 
.A(n_1564),
.B(n_941),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_1300),
.Y(n_2617)
);

AO22x2_ASAP7_75t_L g2618 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2618)
);

OAI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_1300),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1268),
.Y(n_2621)
);

INVxp67_ASAP7_75t_L g2622 ( 
.A(n_1355),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_1300),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_1300),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1268),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_1300),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_1268),
.Y(n_2627)
);

CKINVDCx20_ASAP7_75t_R g2628 ( 
.A(n_1503),
.Y(n_2628)
);

BUFx8_ASAP7_75t_L g2629 ( 
.A(n_1515),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_1560),
.B(n_803),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1560),
.B(n_803),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_1300),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_1268),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_1268),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_1779),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_1268),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_1268),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_1268),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_1268),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_SL g2644 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_1268),
.Y(n_2645)
);

NAND2x1p5_ASAP7_75t_L g2646 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2646)
);

AO22x2_ASAP7_75t_L g2647 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_1268),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_1268),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2650)
);

INVx2_ASAP7_75t_SL g2651 ( 
.A(n_1374),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_1560),
.B(n_803),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_1268),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_1268),
.Y(n_2656)
);

OAI221xp5_ASAP7_75t_L g2657 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_1268),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_1268),
.Y(n_2659)
);

OAI221xp5_ASAP7_75t_L g2660 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2660)
);

INVxp67_ASAP7_75t_L g2661 ( 
.A(n_1355),
.Y(n_2661)
);

AO22x2_ASAP7_75t_L g2662 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2662)
);

INVxp67_ASAP7_75t_L g2663 ( 
.A(n_1355),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_1560),
.B(n_803),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_1268),
.Y(n_2665)
);

OAI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_1650),
.A2(n_803),
.B1(n_1049),
.B2(n_1029),
.Y(n_2666)
);

AOI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_1268),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_R g2669 ( 
.A(n_1730),
.B(n_493),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_1560),
.B(n_803),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_1268),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_1336),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_1560),
.B(n_803),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_1391),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_1268),
.Y(n_2676)
);

CKINVDCx11_ASAP7_75t_R g2677 ( 
.A(n_1503),
.Y(n_2677)
);

AOI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_1268),
.Y(n_2679)
);

AO22x2_ASAP7_75t_L g2680 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_1300),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_1391),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_1560),
.B(n_803),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_1268),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_1268),
.Y(n_2685)
);

AO22x2_ASAP7_75t_L g2686 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1268),
.Y(n_2687)
);

AO22x2_ASAP7_75t_L g2688 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_1268),
.Y(n_2689)
);

AO22x2_ASAP7_75t_L g2690 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_1268),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_1268),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_1268),
.Y(n_2693)
);

AO22x2_ASAP7_75t_L g2694 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2694)
);

AO21x1_ASAP7_75t_L g2695 ( 
.A1(n_1248),
.A2(n_1579),
.B(n_1558),
.Y(n_2695)
);

AO22x2_ASAP7_75t_L g2696 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_1560),
.B(n_803),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_1268),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_1712),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2699)
);

HB1xp67_ASAP7_75t_L g2700 ( 
.A(n_1324),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_1300),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_1268),
.Y(n_2702)
);

NOR2xp67_ASAP7_75t_L g2703 ( 
.A(n_1564),
.B(n_941),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_1560),
.B(n_803),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_1268),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_1300),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_SL g2707 ( 
.A1(n_1560),
.A2(n_675),
.B1(n_837),
.B2(n_1565),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2708)
);

AOI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_1268),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_L g2711 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_1391),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_1560),
.B(n_803),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_1268),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_1268),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_1268),
.Y(n_2717)
);

AND2x4_ASAP7_75t_L g2718 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2719)
);

AO22x2_ASAP7_75t_L g2720 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1560),
.B(n_803),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_1560),
.B(n_803),
.Y(n_2723)
);

AO22x2_ASAP7_75t_L g2724 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2724)
);

AND2x6_ASAP7_75t_SL g2725 ( 
.A(n_1557),
.B(n_967),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_1560),
.B(n_803),
.Y(n_2726)
);

AO22x2_ASAP7_75t_L g2727 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2727)
);

OAI221xp5_ASAP7_75t_L g2728 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2728)
);

OR2x6_ASAP7_75t_L g2729 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2729)
);

AO22x2_ASAP7_75t_L g2730 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_1391),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_1268),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_1268),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_1779),
.Y(n_2734)
);

AO22x2_ASAP7_75t_L g2735 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_1268),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_1355),
.Y(n_2737)
);

BUFx8_ASAP7_75t_L g2738 ( 
.A(n_1515),
.Y(n_2738)
);

INVx4_ASAP7_75t_L g2739 ( 
.A(n_1275),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2740)
);

INVxp67_ASAP7_75t_SL g2741 ( 
.A(n_1347),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_1355),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_1391),
.Y(n_2743)
);

AO22x2_ASAP7_75t_L g2744 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_1268),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_1324),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2747)
);

AO22x2_ASAP7_75t_L g2748 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2748)
);

INVx3_ASAP7_75t_L g2749 ( 
.A(n_1336),
.Y(n_2749)
);

AOI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2750)
);

AND2x4_ASAP7_75t_L g2751 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_1560),
.B(n_803),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_1268),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_1300),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_1268),
.Y(n_2755)
);

AO22x2_ASAP7_75t_L g2756 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2756)
);

NAND2x1p5_ASAP7_75t_L g2757 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_1268),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_1268),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_1560),
.B(n_803),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_1268),
.Y(n_2762)
);

AO22x2_ASAP7_75t_L g2763 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2763)
);

NAND2x1p5_ASAP7_75t_L g2764 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2764)
);

INVxp67_ASAP7_75t_L g2765 ( 
.A(n_1355),
.Y(n_2765)
);

NAND2x1p5_ASAP7_75t_L g2766 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2767)
);

AO22x2_ASAP7_75t_L g2768 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_1268),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_1300),
.Y(n_2770)
);

NAND2x1p5_ASAP7_75t_L g2771 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_1268),
.Y(n_2772)
);

BUFx8_ASAP7_75t_L g2773 ( 
.A(n_1515),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_1268),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_1268),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_1268),
.Y(n_2776)
);

OAI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_1300),
.Y(n_2778)
);

INVxp67_ASAP7_75t_L g2779 ( 
.A(n_1355),
.Y(n_2779)
);

BUFx8_ASAP7_75t_L g2780 ( 
.A(n_1515),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_1268),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_1268),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_1268),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_1268),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_1324),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_1324),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_1268),
.Y(n_2788)
);

AO22x2_ASAP7_75t_L g2789 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_1268),
.Y(n_2791)
);

BUFx8_ASAP7_75t_L g2792 ( 
.A(n_1515),
.Y(n_2792)
);

OAI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_1300),
.Y(n_2794)
);

AO22x2_ASAP7_75t_L g2795 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_1268),
.Y(n_2796)
);

AO22x2_ASAP7_75t_L g2797 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2797)
);

AO22x2_ASAP7_75t_L g2798 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2798)
);

AO22x2_ASAP7_75t_L g2799 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2799)
);

AO22x2_ASAP7_75t_L g2800 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_1268),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_1560),
.B(n_803),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_1300),
.Y(n_2803)
);

NAND2x1p5_ASAP7_75t_L g2804 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_1300),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_1560),
.B(n_803),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_1560),
.B(n_803),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_1560),
.B(n_803),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_1268),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_1560),
.B(n_803),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2811)
);

AOI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_1268),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_1300),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_1268),
.Y(n_2815)
);

CKINVDCx20_ASAP7_75t_R g2816 ( 
.A(n_1503),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_1560),
.B(n_803),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_1560),
.B(n_803),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_SL g2819 ( 
.A(n_1650),
.B(n_1875),
.C(n_1677),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_1560),
.B(n_803),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_1268),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_1268),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_1560),
.B(n_803),
.Y(n_2823)
);

NAND2x1p5_ASAP7_75t_L g2824 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2824)
);

AO22x2_ASAP7_75t_L g2825 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1268),
.Y(n_2826)
);

NAND2x1_ASAP7_75t_L g2827 ( 
.A(n_1392),
.B(n_871),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2828)
);

AO22x2_ASAP7_75t_L g2829 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_1268),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_1268),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_1779),
.Y(n_2833)
);

AO22x2_ASAP7_75t_L g2834 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_1560),
.B(n_803),
.Y(n_2835)
);

INVxp67_ASAP7_75t_L g2836 ( 
.A(n_1355),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_1268),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_1268),
.Y(n_2838)
);

AO22x2_ASAP7_75t_L g2839 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_1560),
.B(n_803),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1268),
.Y(n_2841)
);

AND2x4_ASAP7_75t_L g2842 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_1268),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_1268),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2846)
);

AO22x2_ASAP7_75t_L g2847 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_1300),
.Y(n_2848)
);

AND2x6_ASAP7_75t_L g2849 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2849)
);

OR2x6_ASAP7_75t_L g2850 ( 
.A(n_1318),
.B(n_1319),
.Y(n_2850)
);

AOI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_1560),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2851)
);

NAND2x1p5_ASAP7_75t_L g2852 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_1300),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_1560),
.B(n_803),
.Y(n_2854)
);

OAI221xp5_ASAP7_75t_L g2855 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2855)
);

AO22x2_ASAP7_75t_L g2856 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2856)
);

OAI221xp5_ASAP7_75t_L g2857 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2857)
);

INVx2_ASAP7_75t_SL g2858 ( 
.A(n_1374),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_1268),
.Y(n_2859)
);

AO22x2_ASAP7_75t_L g2860 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2860)
);

AO22x2_ASAP7_75t_L g2861 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2861)
);

AO22x2_ASAP7_75t_L g2862 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2862)
);

OAI221xp5_ASAP7_75t_L g2863 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2864)
);

AND2x4_ASAP7_75t_L g2865 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2865)
);

BUFx8_ASAP7_75t_L g2866 ( 
.A(n_1515),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_1257),
.B(n_1116),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_1268),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_1324),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_1300),
.Y(n_2871)
);

AO22x2_ASAP7_75t_L g2872 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1558),
.B2(n_1579),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_R g2873 ( 
.A(n_1730),
.B(n_493),
.Y(n_2873)
);

OAI221xp5_ASAP7_75t_L g2874 ( 
.A1(n_1650),
.A2(n_1677),
.B1(n_1898),
.B2(n_1875),
.C(n_1255),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_1779),
.Y(n_2875)
);

AO22x2_ASAP7_75t_L g2876 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_1268),
.Y(n_2877)
);

NAND2x1p5_ASAP7_75t_L g2878 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_1905),
.B(n_1560),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_1300),
.Y(n_2880)
);

INVxp67_ASAP7_75t_L g2881 ( 
.A(n_1355),
.Y(n_2881)
);

INVxp67_ASAP7_75t_L g2882 ( 
.A(n_1355),
.Y(n_2882)
);

INVxp67_ASAP7_75t_L g2883 ( 
.A(n_1355),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_1268),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_1268),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_1560),
.B(n_803),
.Y(n_2886)
);

AO22x2_ASAP7_75t_L g2887 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_1268),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_1246),
.B(n_1595),
.Y(n_2889)
);

OAI22xp33_ASAP7_75t_SL g2890 ( 
.A1(n_1712),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_2890)
);

AO22x2_ASAP7_75t_L g2891 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_1268),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_1268),
.Y(n_2894)
);

INVxp67_ASAP7_75t_L g2895 ( 
.A(n_1355),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_1268),
.Y(n_2896)
);

AO22x2_ASAP7_75t_L g2897 ( 
.A1(n_1904),
.A2(n_1558),
.B1(n_1579),
.B2(n_1248),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_1268),
.Y(n_2898)
);

HB1xp67_ASAP7_75t_L g2899 ( 
.A(n_1324),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_1260),
.B(n_1381),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_1268),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_1355),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_1300),
.Y(n_2903)
);

NAND2x1p5_ASAP7_75t_L g2904 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2904)
);

INVxp67_ASAP7_75t_L g2905 ( 
.A(n_1355),
.Y(n_2905)
);

NAND2x1p5_ASAP7_75t_L g2906 ( 
.A(n_1336),
.B(n_1392),
.Y(n_2906)
);

NOR2xp67_ASAP7_75t_L g2907 ( 
.A(n_1564),
.B(n_941),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_1273),
.B(n_1269),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_1268),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_SL g2910 ( 
.A(n_1984),
.B(n_2511),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2043),
.B(n_2049),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2388),
.B(n_2390),
.Y(n_2912)
);

AND2x2_ASAP7_75t_SL g2913 ( 
.A(n_2340),
.B(n_2490),
.Y(n_2913)
);

NOR3xp33_ASAP7_75t_L g2914 ( 
.A(n_1950),
.B(n_2666),
.C(n_1957),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2043),
.B(n_2049),
.Y(n_2915)
);

BUFx12f_ASAP7_75t_L g2916 ( 
.A(n_2305),
.Y(n_2916)
);

AOI21xp33_ASAP7_75t_L g2917 ( 
.A1(n_1928),
.A2(n_1963),
.B(n_2482),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2023),
.B(n_2597),
.Y(n_2918)
);

INVxp67_ASAP7_75t_L g2919 ( 
.A(n_1914),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_2920)
);

AND2x4_ASAP7_75t_L g2921 ( 
.A(n_1948),
.B(n_1987),
.Y(n_2921)
);

AND2x2_ASAP7_75t_SL g2922 ( 
.A(n_2340),
.B(n_2490),
.Y(n_2922)
);

OAI21x1_ASAP7_75t_L g2923 ( 
.A1(n_2277),
.A2(n_2325),
.B(n_2314),
.Y(n_2923)
);

AOI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2212),
.Y(n_2925)
);

OAI22x1_ASAP7_75t_L g2926 ( 
.A1(n_2344),
.A2(n_2348),
.B1(n_2445),
.B2(n_2383),
.Y(n_2926)
);

OAI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2463),
.A2(n_2570),
.B1(n_2610),
.B2(n_2512),
.Y(n_2927)
);

NOR2xp67_ASAP7_75t_L g2928 ( 
.A(n_2156),
.B(n_2229),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_1945),
.B(n_2410),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2063),
.B(n_2081),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2063),
.B(n_2081),
.Y(n_2931)
);

O2A1O1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2890),
.A2(n_1928),
.B(n_2481),
.C(n_2419),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2014),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2212),
.Y(n_2934)
);

O2A1O1Ixp5_ASAP7_75t_L g2935 ( 
.A1(n_2419),
.A2(n_2481),
.B(n_2644),
.C(n_2485),
.Y(n_2935)
);

OAI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2650),
.A2(n_2653),
.B1(n_2678),
.B2(n_2667),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2410),
.A2(n_2634),
.B1(n_2654),
.B2(n_2467),
.Y(n_2937)
);

HB1xp67_ASAP7_75t_L g2938 ( 
.A(n_2212),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2485),
.A2(n_2719),
.B(n_2644),
.Y(n_2939)
);

INVx4_ASAP7_75t_L g2940 ( 
.A(n_1948),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2212),
.Y(n_2941)
);

AOI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2719),
.A2(n_2867),
.B(n_2785),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2014),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_1918),
.B(n_2116),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2467),
.B(n_2634),
.Y(n_2945)
);

AOI21xp33_ASAP7_75t_L g2946 ( 
.A1(n_2785),
.A2(n_2867),
.B(n_1946),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2277),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2110),
.A2(n_1911),
.B(n_1910),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2110),
.A2(n_1911),
.B(n_1910),
.Y(n_2949)
);

INVxp67_ASAP7_75t_SL g2950 ( 
.A(n_2695),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2216),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_1946),
.A2(n_2345),
.B(n_2407),
.C(n_2349),
.Y(n_2952)
);

OAI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_1918),
.A2(n_2699),
.B(n_2566),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2388),
.B(n_2390),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_L g2955 ( 
.A(n_2654),
.B(n_2711),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_1910),
.A2(n_1920),
.B(n_1911),
.Y(n_2956)
);

BUFx4f_ASAP7_75t_L g2957 ( 
.A(n_2031),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_1910),
.A2(n_1920),
.B(n_1911),
.Y(n_2958)
);

BUFx4f_ASAP7_75t_L g2959 ( 
.A(n_2031),
.Y(n_2959)
);

OAI21xp33_ASAP7_75t_L g2960 ( 
.A1(n_2708),
.A2(n_2747),
.B(n_2709),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2116),
.B(n_2121),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2711),
.B(n_2879),
.Y(n_2962)
);

AOI22xp5_ASAP7_75t_L g2963 ( 
.A1(n_2879),
.A2(n_2819),
.B1(n_2812),
.B2(n_2750),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_SL g2964 ( 
.A(n_2201),
.B(n_1923),
.Y(n_2964)
);

AOI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_1920),
.A2(n_1936),
.B(n_1930),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2121),
.B(n_2042),
.Y(n_2966)
);

OAI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2566),
.A2(n_2699),
.B(n_2027),
.Y(n_2967)
);

AOI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_1920),
.A2(n_1936),
.B(n_1930),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2388),
.B(n_2390),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2126),
.B(n_2070),
.Y(n_2970)
);

INVxp67_ASAP7_75t_L g2971 ( 
.A(n_2439),
.Y(n_2971)
);

O2A1O1Ixp33_ASAP7_75t_L g2972 ( 
.A1(n_2431),
.A2(n_2444),
.B(n_2456),
.C(n_2451),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_1916),
.B(n_1926),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2228),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2228),
.Y(n_2975)
);

AOI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2828),
.A2(n_2851),
.B1(n_2846),
.B2(n_2476),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_1930),
.A2(n_2341),
.B(n_1936),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_1951),
.B(n_1953),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_1932),
.A2(n_2516),
.B(n_2619),
.C(n_2519),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2032),
.B(n_2047),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_1955),
.B(n_1959),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_1930),
.A2(n_2341),
.B(n_1936),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2341),
.A2(n_2346),
.B(n_2343),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_1923),
.B(n_2187),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2047),
.B(n_2391),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2391),
.B(n_2393),
.Y(n_2986)
);

BUFx4f_ASAP7_75t_L g2987 ( 
.A(n_2031),
.Y(n_2987)
);

AOI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2341),
.A2(n_2346),
.B(n_2343),
.Y(n_2988)
);

AOI21xp33_ASAP7_75t_L g2989 ( 
.A1(n_2391),
.A2(n_2399),
.B(n_2393),
.Y(n_2989)
);

BUFx4f_ASAP7_75t_L g2990 ( 
.A(n_2031),
.Y(n_2990)
);

OAI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_1970),
.A2(n_2493),
.B(n_2404),
.Y(n_2991)
);

BUFx4f_ASAP7_75t_L g2992 ( 
.A(n_2031),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2351),
.A2(n_2359),
.B1(n_2361),
.B2(n_2353),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_2669),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2363),
.A2(n_2365),
.B1(n_2394),
.B2(n_2364),
.Y(n_2995)
);

AOI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2343),
.A2(n_2350),
.B(n_2346),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2393),
.B(n_2399),
.Y(n_2997)
);

INVx3_ASAP7_75t_L g2998 ( 
.A(n_2277),
.Y(n_2998)
);

AOI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2343),
.A2(n_2350),
.B(n_2346),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2350),
.A2(n_2366),
.B(n_2356),
.Y(n_3000)
);

AO21x2_ASAP7_75t_L g3001 ( 
.A1(n_2173),
.A2(n_2695),
.B(n_2325),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2399),
.B(n_2416),
.Y(n_3002)
);

OAI21xp5_ASAP7_75t_L g3003 ( 
.A1(n_1970),
.A2(n_2493),
.B(n_2404),
.Y(n_3003)
);

INVx2_ASAP7_75t_SL g3004 ( 
.A(n_2314),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2228),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_1922),
.Y(n_3006)
);

CKINVDCx16_ASAP7_75t_R g3007 ( 
.A(n_2669),
.Y(n_3007)
);

INVx11_ASAP7_75t_L g3008 ( 
.A(n_2252),
.Y(n_3008)
);

AOI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2657),
.A2(n_2660),
.B1(n_2777),
.B2(n_2728),
.Y(n_3009)
);

BUFx3_ASAP7_75t_L g3010 ( 
.A(n_2074),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2908),
.A2(n_2173),
.B(n_2114),
.Y(n_3011)
);

O2A1O1Ixp33_ASAP7_75t_SL g3012 ( 
.A1(n_2034),
.A2(n_2079),
.B(n_2086),
.C(n_2067),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2235),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2400),
.B(n_2418),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2416),
.B(n_2443),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2416),
.B(n_2443),
.Y(n_3016)
);

OAI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2908),
.A2(n_2855),
.B(n_2793),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2443),
.B(n_2475),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2475),
.B(n_2488),
.Y(n_3019)
);

INVxp67_ASAP7_75t_L g3020 ( 
.A(n_2563),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2350),
.A2(n_2366),
.B(n_2356),
.Y(n_3021)
);

AOI22x1_ASAP7_75t_L g3022 ( 
.A1(n_2475),
.A2(n_2686),
.B1(n_2688),
.B2(n_2488),
.Y(n_3022)
);

INVx4_ASAP7_75t_L g3023 ( 
.A(n_1948),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2488),
.B(n_2686),
.Y(n_3024)
);

NAND2x1p5_ASAP7_75t_L g3025 ( 
.A(n_2220),
.B(n_2287),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2356),
.A2(n_2373),
.B(n_2366),
.Y(n_3026)
);

BUFx6f_ASAP7_75t_L g3027 ( 
.A(n_1948),
.Y(n_3027)
);

OR2x6_ASAP7_75t_L g3028 ( 
.A(n_2310),
.B(n_2312),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2686),
.B(n_2688),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2356),
.A2(n_2373),
.B(n_2366),
.Y(n_3030)
);

OAI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2857),
.A2(n_2874),
.B(n_2863),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2688),
.B(n_2690),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2373),
.A2(n_2524),
.B(n_2502),
.Y(n_3033)
);

AOI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2473),
.A2(n_2454),
.B1(n_2468),
.B2(n_2460),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2690),
.B(n_2694),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2373),
.A2(n_2524),
.B(n_2502),
.Y(n_3036)
);

OAI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_2472),
.A2(n_2507),
.B1(n_2508),
.B2(n_2477),
.Y(n_3037)
);

OAI321xp33_ASAP7_75t_L g3038 ( 
.A1(n_2019),
.A2(n_2020),
.A3(n_1983),
.B1(n_2036),
.B2(n_2088),
.C(n_2038),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_1987),
.B(n_2352),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_L g3040 ( 
.A(n_2518),
.B(n_2529),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2235),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_1988),
.A2(n_2707),
.B(n_2026),
.C(n_2147),
.Y(n_3042)
);

CKINVDCx10_ASAP7_75t_R g3043 ( 
.A(n_2075),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2690),
.B(n_2694),
.Y(n_3044)
);

A2O1A1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_2473),
.A2(n_2607),
.B(n_2609),
.C(n_2605),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2502),
.A2(n_2527),
.B(n_2524),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2694),
.B(n_2696),
.Y(n_3047)
);

OAI22xp5_ASAP7_75t_L g3048 ( 
.A1(n_2614),
.A2(n_2633),
.B1(n_2652),
.B2(n_2631),
.Y(n_3048)
);

BUFx8_ASAP7_75t_L g3049 ( 
.A(n_2075),
.Y(n_3049)
);

NAND3xp33_ASAP7_75t_SL g3050 ( 
.A(n_2664),
.B(n_2673),
.C(n_2670),
.Y(n_3050)
);

A2O1A1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_2683),
.A2(n_2704),
.B(n_2714),
.C(n_2697),
.Y(n_3051)
);

AOI21x1_ASAP7_75t_L g3052 ( 
.A1(n_2005),
.A2(n_2524),
.B(n_2502),
.Y(n_3052)
);

O2A1O1Ixp33_ASAP7_75t_L g3053 ( 
.A1(n_2722),
.A2(n_2726),
.B(n_2752),
.C(n_2723),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2527),
.A2(n_2539),
.B(n_2534),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2696),
.B(n_2720),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2696),
.B(n_2720),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2873),
.B(n_2161),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2527),
.A2(n_2539),
.B(n_2534),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2873),
.B(n_2004),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2720),
.B(n_2724),
.Y(n_3060)
);

OAI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2021),
.A2(n_2136),
.B(n_2210),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2527),
.A2(n_2539),
.B(n_2534),
.Y(n_3062)
);

BUFx3_ASAP7_75t_L g3063 ( 
.A(n_2074),
.Y(n_3063)
);

NAND3xp33_ASAP7_75t_L g3064 ( 
.A(n_2761),
.B(n_2806),
.C(n_2802),
.Y(n_3064)
);

OAI321xp33_ASAP7_75t_L g3065 ( 
.A1(n_2807),
.A2(n_2808),
.A3(n_2810),
.B1(n_2820),
.B2(n_2818),
.C(n_2817),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_2004),
.B(n_1947),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_1922),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2238),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2534),
.A2(n_2543),
.B(n_2539),
.Y(n_3069)
);

OA21x2_ASAP7_75t_L g3070 ( 
.A1(n_2183),
.A2(n_2240),
.B(n_2218),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2543),
.A2(n_2550),
.B(n_2546),
.Y(n_3071)
);

HB1xp67_ASAP7_75t_L g3072 ( 
.A(n_2238),
.Y(n_3072)
);

OAI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2179),
.A2(n_2183),
.B(n_2021),
.Y(n_3073)
);

AOI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2543),
.A2(n_2550),
.B(n_2546),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2823),
.B(n_2835),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2724),
.B(n_2727),
.Y(n_3076)
);

O2A1O1Ixp33_ASAP7_75t_SL g3077 ( 
.A1(n_2098),
.A2(n_2108),
.B(n_2016),
.C(n_2007),
.Y(n_3077)
);

BUFx6f_ASAP7_75t_L g3078 ( 
.A(n_1987),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2840),
.A2(n_2854),
.B1(n_2886),
.B2(n_1977),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2543),
.A2(n_2550),
.B(n_2546),
.Y(n_3080)
);

OAI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2724),
.A2(n_2730),
.B1(n_2735),
.B2(n_2727),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_1964),
.B(n_2134),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_L g3083 ( 
.A1(n_1977),
.A2(n_2730),
.B1(n_2735),
.B2(n_2727),
.Y(n_3083)
);

AOI21x1_ASAP7_75t_L g3084 ( 
.A1(n_2005),
.A2(n_2550),
.B(n_2546),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2558),
.Y(n_3085)
);

OR2x6_ASAP7_75t_SL g3086 ( 
.A(n_2185),
.B(n_2557),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2558),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2530),
.B(n_2131),
.Y(n_3088)
);

AOI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2558),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2558),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2730),
.B(n_2735),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2582),
.A2(n_2594),
.B(n_2591),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2744),
.B(n_2748),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2163),
.Y(n_3094)
);

OR2x6_ASAP7_75t_L g3095 ( 
.A(n_2310),
.B(n_2312),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2530),
.B(n_2124),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2582),
.A2(n_2594),
.B(n_2591),
.Y(n_3097)
);

CKINVDCx5p33_ASAP7_75t_R g3098 ( 
.A(n_2509),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2146),
.B(n_2166),
.Y(n_3099)
);

BUFx4f_ASAP7_75t_L g3100 ( 
.A(n_2031),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2744),
.B(n_2748),
.Y(n_3101)
);

O2A1O1Ixp5_ASAP7_75t_L g3102 ( 
.A1(n_2205),
.A2(n_2311),
.B(n_2240),
.C(n_2248),
.Y(n_3102)
);

AOI22xp33_ASAP7_75t_SL g3103 ( 
.A1(n_1977),
.A2(n_2797),
.B1(n_2748),
.B2(n_2756),
.Y(n_3103)
);

OAI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2292),
.A2(n_2203),
.B(n_2154),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2744),
.A2(n_2763),
.B1(n_2768),
.B2(n_2756),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_L g3106 ( 
.A(n_1987),
.Y(n_3106)
);

AOI21x1_ASAP7_75t_L g3107 ( 
.A1(n_2005),
.A2(n_2594),
.B(n_2591),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2591),
.A2(n_2601),
.B(n_2594),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2158),
.A2(n_2198),
.B(n_2220),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2601),
.A2(n_2603),
.B(n_2602),
.Y(n_3110)
);

NAND2x1p5_ASAP7_75t_L g3111 ( 
.A(n_2205),
.B(n_2218),
.Y(n_3111)
);

O2A1O1Ixp33_ASAP7_75t_L g3112 ( 
.A1(n_2207),
.A2(n_2437),
.B(n_2741),
.C(n_2422),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2601),
.A2(n_2603),
.B(n_2602),
.Y(n_3113)
);

AOI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2601),
.A2(n_2603),
.B(n_2602),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2756),
.B(n_2763),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2163),
.Y(n_3116)
);

BUFx12f_ASAP7_75t_L g3117 ( 
.A(n_2305),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_L g3118 ( 
.A(n_1935),
.B(n_2339),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2602),
.A2(n_2608),
.B(n_2603),
.Y(n_3119)
);

O2A1O1Ixp33_ASAP7_75t_L g3120 ( 
.A1(n_1998),
.A2(n_2029),
.B(n_2244),
.C(n_2330),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2763),
.B(n_2768),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2608),
.A2(n_2647),
.B(n_2618),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2608),
.A2(n_2647),
.B(n_2618),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2768),
.B(n_2789),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2608),
.A2(n_2647),
.B(n_2618),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2789),
.B(n_2795),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2618),
.A2(n_2662),
.B(n_2647),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2163),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2789),
.B(n_2795),
.Y(n_3129)
);

OR2x2_ASAP7_75t_L g3130 ( 
.A(n_2352),
.B(n_2599),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2795),
.B(n_2797),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2411),
.Y(n_3132)
);

CKINVDCx20_ASAP7_75t_R g3133 ( 
.A(n_2509),
.Y(n_3133)
);

AOI21x1_ASAP7_75t_L g3134 ( 
.A1(n_2662),
.A2(n_2876),
.B(n_2680),
.Y(n_3134)
);

INVx3_ASAP7_75t_L g3135 ( 
.A(n_1925),
.Y(n_3135)
);

INVx4_ASAP7_75t_L g3136 ( 
.A(n_2352),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2662),
.A2(n_2876),
.B(n_2680),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2662),
.A2(n_2876),
.B(n_2680),
.Y(n_3138)
);

AO22x1_ASAP7_75t_L g3139 ( 
.A1(n_2273),
.A2(n_2316),
.B1(n_2318),
.B2(n_2317),
.Y(n_3139)
);

AOI21x1_ASAP7_75t_L g3140 ( 
.A1(n_2876),
.A2(n_2891),
.B(n_2887),
.Y(n_3140)
);

INVxp67_ASAP7_75t_L g3141 ( 
.A(n_2700),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_2887),
.A2(n_2897),
.B(n_2891),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2887),
.A2(n_2897),
.B(n_2891),
.Y(n_3143)
);

AOI21x1_ASAP7_75t_L g3144 ( 
.A1(n_2887),
.A2(n_2897),
.B(n_2891),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2897),
.A2(n_1968),
.B(n_1961),
.Y(n_3145)
);

A2O1A1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_2072),
.A2(n_2076),
.B(n_2077),
.C(n_2073),
.Y(n_3146)
);

AOI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_1961),
.A2(n_1972),
.B(n_1968),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2797),
.B(n_2798),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2798),
.B(n_2799),
.Y(n_3149)
);

AOI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2798),
.A2(n_2800),
.B1(n_2825),
.B2(n_2799),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2799),
.B(n_2800),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2800),
.B(n_2825),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_1961),
.A2(n_1972),
.B(n_1968),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_1964),
.B(n_1913),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2825),
.B(n_2829),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_1972),
.A2(n_1974),
.B(n_2829),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_2301),
.B(n_2248),
.Y(n_3157)
);

OAI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_2829),
.A2(n_2839),
.B1(n_2847),
.B2(n_2834),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_L g3159 ( 
.A(n_1913),
.B(n_1938),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2834),
.B(n_2839),
.Y(n_3160)
);

AOI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_2834),
.A2(n_2839),
.B1(n_2856),
.B2(n_2847),
.Y(n_3161)
);

NOR2xp33_ASAP7_75t_L g3162 ( 
.A(n_1938),
.B(n_1956),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_2352),
.B(n_2599),
.Y(n_3163)
);

AOI22xp5_ASAP7_75t_L g3164 ( 
.A1(n_2847),
.A2(n_2856),
.B1(n_2861),
.B2(n_2860),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_2599),
.B(n_2729),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_1974),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_2179),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_1974),
.A2(n_2860),
.B(n_2856),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2599),
.Y(n_3169)
);

OAI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2175),
.A2(n_2311),
.B(n_2268),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2860),
.B(n_2861),
.Y(n_3171)
);

O2A1O1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_2010),
.A2(n_1980),
.B(n_2441),
.C(n_2397),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_1956),
.B(n_1962),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2861),
.A2(n_2872),
.B(n_2862),
.Y(n_3174)
);

OAI21x1_ASAP7_75t_L g3175 ( 
.A1(n_2261),
.A2(n_2268),
.B(n_1933),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2163),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2862),
.A2(n_2872),
.B(n_2261),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2862),
.A2(n_2872),
.B(n_2335),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_1997),
.B(n_2131),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2141),
.A2(n_2149),
.B(n_2304),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2145),
.Y(n_3181)
);

BUFx6f_ASAP7_75t_L g3182 ( 
.A(n_2729),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2335),
.A2(n_1997),
.B(n_2312),
.Y(n_3183)
);

NAND2x1p5_ASAP7_75t_L g3184 ( 
.A(n_1925),
.B(n_1933),
.Y(n_3184)
);

BUFx6f_ASAP7_75t_L g3185 ( 
.A(n_2729),
.Y(n_3185)
);

OR2x6_ASAP7_75t_L g3186 ( 
.A(n_2310),
.B(n_2162),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_1937),
.Y(n_3187)
);

A2O1A1Ixp33_ASAP7_75t_L g3188 ( 
.A1(n_2080),
.A2(n_2087),
.B(n_2090),
.C(n_2084),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_1997),
.B(n_2335),
.Y(n_3189)
);

INVx2_ASAP7_75t_SL g3190 ( 
.A(n_2729),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2145),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_1937),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_1944),
.Y(n_3193)
);

OAI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2097),
.A2(n_2102),
.B1(n_2103),
.B2(n_2101),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2018),
.A2(n_2025),
.B(n_2083),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2018),
.A2(n_2025),
.B(n_2083),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2162),
.B(n_2083),
.Y(n_3197)
);

OAI321xp33_ASAP7_75t_L g3198 ( 
.A1(n_2091),
.A2(n_2421),
.A3(n_1991),
.B1(n_2427),
.B2(n_2338),
.C(n_1962),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2145),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2106),
.B(n_2111),
.Y(n_3200)
);

NAND3xp33_ASAP7_75t_L g3201 ( 
.A(n_2148),
.B(n_2478),
.C(n_2449),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2037),
.Y(n_3202)
);

OAI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2304),
.A2(n_2321),
.B(n_2319),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2113),
.B(n_2119),
.Y(n_3204)
);

OAI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2322),
.A2(n_2424),
.B(n_2375),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_2018),
.A2(n_2025),
.B(n_2083),
.Y(n_3206)
);

OR2x2_ASAP7_75t_L g3207 ( 
.A(n_2850),
.B(n_2358),
.Y(n_3207)
);

A2O1A1Ixp33_ASAP7_75t_L g3208 ( 
.A1(n_2160),
.A2(n_2425),
.B(n_2489),
.C(n_2457),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2037),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2085),
.A2(n_2093),
.B(n_2092),
.Y(n_3210)
);

OAI22xp5_ASAP7_75t_L g3211 ( 
.A1(n_1991),
.A2(n_2421),
.B1(n_2427),
.B2(n_2338),
.Y(n_3211)
);

CKINVDCx8_ASAP7_75t_R g3212 ( 
.A(n_2725),
.Y(n_3212)
);

AND2x4_ASAP7_75t_L g3213 ( 
.A(n_2850),
.B(n_2375),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2850),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2085),
.A2(n_2093),
.B(n_2092),
.Y(n_3215)
);

INVx6_ASAP7_75t_L g3216 ( 
.A(n_2252),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2033),
.B(n_2040),
.Y(n_3217)
);

CKINVDCx8_ASAP7_75t_R g3218 ( 
.A(n_2192),
.Y(n_3218)
);

NOR2x1p5_ASAP7_75t_SL g3219 ( 
.A(n_2089),
.B(n_2095),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2085),
.A2(n_2093),
.B(n_2092),
.Y(n_3220)
);

NAND3xp33_ASAP7_75t_SL g3221 ( 
.A(n_2112),
.B(n_2289),
.C(n_1941),
.Y(n_3221)
);

OR2x6_ASAP7_75t_L g3222 ( 
.A(n_2162),
.B(n_2850),
.Y(n_3222)
);

AOI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_2085),
.A2(n_2093),
.B(n_2092),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2033),
.B(n_2040),
.Y(n_3224)
);

A2O1A1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_2616),
.A2(n_2703),
.B(n_2907),
.C(n_2288),
.Y(n_3225)
);

OAI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2375),
.A2(n_2849),
.B(n_2424),
.Y(n_3226)
);

O2A1O1Ixp5_ASAP7_75t_L g3227 ( 
.A1(n_2269),
.A2(n_2326),
.B(n_2095),
.C(n_2099),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2145),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2153),
.Y(n_3229)
);

A2O1A1Ixp33_ASAP7_75t_L g3230 ( 
.A1(n_2164),
.A2(n_2307),
.B(n_2267),
.C(n_2181),
.Y(n_3230)
);

AO22x1_ASAP7_75t_L g3231 ( 
.A1(n_2164),
.A2(n_2109),
.B1(n_2096),
.B2(n_2125),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2411),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2033),
.B(n_2040),
.Y(n_3233)
);

OAI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2375),
.A2(n_2849),
.B(n_2424),
.Y(n_3234)
);

AOI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2452),
.A2(n_2494),
.B1(n_2499),
.B2(n_2458),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_2162),
.B(n_2100),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_2100),
.A2(n_2117),
.B(n_2105),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_2375),
.B(n_2424),
.Y(n_3238)
);

INVx1_ASAP7_75t_SL g3239 ( 
.A(n_2358),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2089),
.Y(n_3240)
);

O2A1O1Ixp33_ASAP7_75t_L g3241 ( 
.A1(n_2483),
.A2(n_2525),
.B(n_2572),
.C(n_2484),
.Y(n_3241)
);

AND3x2_ASAP7_75t_L g3242 ( 
.A(n_2192),
.B(n_2263),
.C(n_2230),
.Y(n_3242)
);

INVx11_ASAP7_75t_L g3243 ( 
.A(n_2252),
.Y(n_3243)
);

CKINVDCx5p33_ASAP7_75t_R g3244 ( 
.A(n_2677),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2452),
.A2(n_2494),
.B1(n_2499),
.B2(n_2458),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_1927),
.B(n_1940),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_2375),
.B(n_2424),
.Y(n_3247)
);

AOI22x1_ASAP7_75t_L g3248 ( 
.A1(n_2144),
.A2(n_2064),
.B1(n_2066),
.B2(n_2057),
.Y(n_3248)
);

A2O1A1Ixp33_ASAP7_75t_L g3249 ( 
.A1(n_2164),
.A2(n_2267),
.B(n_2181),
.C(n_2528),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2057),
.B(n_2064),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_2100),
.A2(n_2117),
.B(n_2105),
.Y(n_3251)
);

AND2x2_ASAP7_75t_SL g3252 ( 
.A(n_2100),
.B(n_2105),
.Y(n_3252)
);

OR2x2_ASAP7_75t_L g3253 ( 
.A(n_2553),
.B(n_2604),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2057),
.B(n_2064),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2105),
.B(n_2117),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_2553),
.Y(n_3256)
);

O2A1O1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_2590),
.A2(n_2661),
.B(n_2663),
.C(n_2622),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2737),
.B(n_2742),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2099),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_2424),
.Y(n_3260)
);

NAND3xp33_ASAP7_75t_L g3261 ( 
.A(n_2765),
.B(n_2836),
.C(n_2779),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_2117),
.A2(n_2118),
.B(n_2269),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2066),
.B(n_2071),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_2118),
.B(n_2066),
.Y(n_3264)
);

A2O1A1Ixp33_ASAP7_75t_L g3265 ( 
.A1(n_2528),
.A2(n_2588),
.B(n_2630),
.C(n_2549),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_2118),
.B(n_2071),
.Y(n_3266)
);

AND2x4_ASAP7_75t_L g3267 ( 
.A(n_2849),
.B(n_2143),
.Y(n_3267)
);

A2O1A1Ixp33_ASAP7_75t_L g3268 ( 
.A1(n_2549),
.A2(n_2630),
.B(n_2632),
.C(n_2588),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2118),
.A2(n_2903),
.B(n_2143),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2903),
.A2(n_2170),
.B(n_2115),
.Y(n_3270)
);

INVxp33_ASAP7_75t_SL g3271 ( 
.A(n_2142),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2153),
.Y(n_3272)
);

AOI21x1_ASAP7_75t_L g3273 ( 
.A1(n_2071),
.A2(n_2078),
.B(n_2157),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_2115),
.A2(n_2171),
.B(n_2170),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_2881),
.B(n_2882),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2171),
.A2(n_2200),
.B(n_2194),
.Y(n_3276)
);

INVx2_ASAP7_75t_SL g3277 ( 
.A(n_2194),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_2078),
.B(n_2153),
.Y(n_3278)
);

OAI21xp33_ASAP7_75t_L g3279 ( 
.A1(n_2632),
.A2(n_2721),
.B(n_2638),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2078),
.B(n_2638),
.Y(n_3280)
);

OAI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_2849),
.A2(n_2256),
.B(n_2246),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2200),
.A2(n_2370),
.B(n_2368),
.Y(n_3282)
);

AOI21xp33_ASAP7_75t_L g3283 ( 
.A1(n_2144),
.A2(n_2188),
.B(n_2167),
.Y(n_3283)
);

INVx3_ASAP7_75t_L g3284 ( 
.A(n_2368),
.Y(n_3284)
);

O2A1O1Ixp33_ASAP7_75t_L g3285 ( 
.A1(n_2883),
.A2(n_2902),
.B(n_2905),
.C(n_2895),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_2370),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2721),
.B(n_2740),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2371),
.A2(n_2385),
.B(n_2381),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2740),
.A2(n_2790),
.B1(n_2843),
.B2(n_2811),
.Y(n_3289)
);

BUFx2_ASAP7_75t_L g3290 ( 
.A(n_2285),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_2371),
.A2(n_2385),
.B(n_2381),
.Y(n_3291)
);

OAI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2849),
.A2(n_2256),
.B(n_2246),
.Y(n_3292)
);

NAND2xp33_ASAP7_75t_L g3293 ( 
.A(n_2107),
.B(n_2142),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2790),
.B(n_2811),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2843),
.B(n_2889),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2889),
.B(n_2144),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_2604),
.B(n_2378),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2157),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_2392),
.A2(n_2433),
.B(n_2432),
.Y(n_3299)
);

BUFx4f_ASAP7_75t_L g3300 ( 
.A(n_2849),
.Y(n_3300)
);

OAI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_2262),
.A2(n_2432),
.B(n_2392),
.Y(n_3301)
);

OAI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2262),
.A2(n_2470),
.B(n_2433),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2144),
.B(n_2196),
.Y(n_3303)
);

NOR2xp33_ASAP7_75t_L g3304 ( 
.A(n_2532),
.B(n_1949),
.Y(n_3304)
);

BUFx2_ASAP7_75t_L g3305 ( 
.A(n_2285),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_SL g3306 ( 
.A(n_2378),
.B(n_2387),
.Y(n_3306)
);

AOI21x1_ASAP7_75t_L g3307 ( 
.A1(n_2157),
.A2(n_2188),
.B(n_2167),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2470),
.Y(n_3308)
);

OAI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_2486),
.A2(n_2526),
.B(n_2496),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_SL g3310 ( 
.A(n_2387),
.B(n_2442),
.Y(n_3310)
);

BUFx6f_ASAP7_75t_L g3311 ( 
.A(n_2486),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2496),
.A2(n_2531),
.B(n_2526),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2174),
.B(n_2028),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2531),
.A2(n_2548),
.B(n_2544),
.Y(n_3314)
);

NAND2x1p5_ASAP7_75t_L g3315 ( 
.A(n_2544),
.B(n_2548),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_2554),
.A2(n_2564),
.B(n_2559),
.Y(n_3316)
);

NAND2xp33_ASAP7_75t_L g3317 ( 
.A(n_2107),
.B(n_2191),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2196),
.B(n_2167),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2554),
.A2(n_2564),
.B(n_2559),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2157),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2196),
.B(n_2167),
.Y(n_3321)
);

A2O1A1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_2286),
.A2(n_2270),
.B(n_2282),
.C(n_2326),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2573),
.A2(n_2617),
.B(n_2596),
.Y(n_3323)
);

A2O1A1Ixp33_ASAP7_75t_L g3324 ( 
.A1(n_2270),
.A2(n_2137),
.B(n_2231),
.C(n_2024),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2442),
.B(n_2651),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2196),
.B(n_1908),
.Y(n_3326)
);

CKINVDCx10_ASAP7_75t_R g3327 ( 
.A(n_2075),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_1915),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2573),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2011),
.A2(n_2858),
.B1(n_2651),
.B2(n_2069),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_1917),
.B(n_1919),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_2858),
.A2(n_2188),
.B1(n_2209),
.B2(n_2169),
.Y(n_3332)
);

AOI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_2596),
.A2(n_2620),
.B(n_2617),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_1921),
.B(n_1929),
.Y(n_3334)
);

AOI22xp5_ASAP7_75t_L g3335 ( 
.A1(n_2062),
.A2(n_2250),
.B1(n_2270),
.B2(n_1967),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_1931),
.B(n_1934),
.Y(n_3336)
);

OAI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_1939),
.A2(n_1943),
.B1(n_1952),
.B2(n_1942),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_1954),
.B(n_1958),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_1960),
.B(n_1965),
.Y(n_3339)
);

BUFx8_ASAP7_75t_SL g3340 ( 
.A(n_1996),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2620),
.Y(n_3341)
);

INVx11_ASAP7_75t_L g3342 ( 
.A(n_2096),
.Y(n_3342)
);

NAND3xp33_ASAP7_75t_L g3343 ( 
.A(n_2746),
.B(n_2787),
.C(n_2786),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2870),
.B(n_2899),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_2623),
.A2(n_2626),
.B(n_2624),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_1969),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_1973),
.B(n_1975),
.Y(n_3347)
);

BUFx6f_ASAP7_75t_L g3348 ( 
.A(n_2623),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_1967),
.A2(n_2382),
.B1(n_2503),
.B2(n_2165),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_2295),
.B(n_2176),
.Y(n_3350)
);

OAI22xp5_ASAP7_75t_L g3351 ( 
.A1(n_1976),
.A2(n_1978),
.B1(n_1981),
.B2(n_1979),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2624),
.A2(n_2635),
.B(n_2626),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_2635),
.A2(n_2701),
.B(n_2681),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_2681),
.A2(n_2706),
.B(n_2701),
.Y(n_3354)
);

NOR2xp67_ASAP7_75t_L g3355 ( 
.A(n_2372),
.B(n_2446),
.Y(n_3355)
);

O2A1O1Ixp33_ASAP7_75t_L g3356 ( 
.A1(n_1971),
.A2(n_2132),
.B(n_1989),
.C(n_2315),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_2706),
.A2(n_2770),
.B(n_2754),
.Y(n_3357)
);

AOI21x1_ASAP7_75t_L g3358 ( 
.A1(n_2188),
.A2(n_2276),
.B(n_2275),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2754),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_2778),
.A2(n_2803),
.B(n_2794),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_2803),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_1989),
.B(n_2255),
.Y(n_3362)
);

NOR2x1_ASAP7_75t_L g3363 ( 
.A(n_2805),
.B(n_2814),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_1982),
.B(n_1986),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_2805),
.A2(n_2848),
.B(n_2814),
.Y(n_3365)
);

BUFx2_ASAP7_75t_L g3366 ( 
.A(n_2276),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_2848),
.A2(n_2871),
.B(n_2853),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_1990),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_1992),
.B(n_1993),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_1995),
.Y(n_3370)
);

O2A1O1Ixp33_ASAP7_75t_L g3371 ( 
.A1(n_2120),
.A2(n_2123),
.B(n_2128),
.C(n_2122),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2853),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_2001),
.B(n_2002),
.Y(n_3373)
);

NAND3xp33_ASAP7_75t_L g3374 ( 
.A(n_2177),
.B(n_2182),
.C(n_2180),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_2677),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2006),
.B(n_2008),
.Y(n_3376)
);

BUFx6f_ASAP7_75t_L g3377 ( 
.A(n_2871),
.Y(n_3377)
);

AOI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_2880),
.A2(n_2275),
.B(n_2302),
.Y(n_3378)
);

BUFx6f_ASAP7_75t_L g3379 ( 
.A(n_2880),
.Y(n_3379)
);

OAI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_2012),
.A2(n_2015),
.B1(n_2017),
.B2(n_2013),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_L g3381 ( 
.A(n_2165),
.B(n_2191),
.Y(n_3381)
);

AOI222xp33_ASAP7_75t_L g3382 ( 
.A1(n_2022),
.A2(n_2030),
.B1(n_2044),
.B2(n_2046),
.C1(n_2045),
.C2(n_2035),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_2165),
.B(n_2298),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2051),
.Y(n_3384)
);

NOR3xp33_ASAP7_75t_L g3385 ( 
.A(n_2284),
.B(n_2334),
.C(n_2239),
.Y(n_3385)
);

INVx4_ASAP7_75t_L g3386 ( 
.A(n_2372),
.Y(n_3386)
);

AOI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_1967),
.A2(n_2382),
.B1(n_2503),
.B2(n_2209),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_2255),
.B(n_2294),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_2276),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2275),
.A2(n_2209),
.B(n_2827),
.Y(n_3390)
);

CKINVDCx14_ASAP7_75t_R g3391 ( 
.A(n_2009),
.Y(n_3391)
);

INVx3_ASAP7_75t_L g3392 ( 
.A(n_2372),
.Y(n_3392)
);

NOR3xp33_ASAP7_75t_L g3393 ( 
.A(n_2329),
.B(n_2263),
.C(n_2230),
.Y(n_3393)
);

OR2x2_ASAP7_75t_L g3394 ( 
.A(n_2130),
.B(n_2133),
.Y(n_3394)
);

OAI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_2172),
.A2(n_2186),
.B(n_2184),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2197),
.B(n_2206),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_2197),
.B(n_2206),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_2209),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2053),
.B(n_2055),
.Y(n_3399)
);

OAI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_2172),
.A2(n_2195),
.B(n_2189),
.Y(n_3400)
);

OAI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_2172),
.A2(n_2204),
.B(n_2199),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2056),
.B(n_2058),
.Y(n_3402)
);

A2O1A1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_2231),
.A2(n_2061),
.B(n_2065),
.C(n_2060),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_2068),
.B(n_2342),
.Y(n_3404)
);

O2A1O1Ixp5_ASAP7_75t_L g3405 ( 
.A1(n_2138),
.A2(n_2139),
.B(n_2536),
.C(n_2446),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2347),
.B(n_2354),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2355),
.Y(n_3407)
);

BUFx6f_ASAP7_75t_L g3408 ( 
.A(n_2446),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2360),
.B(n_2362),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2367),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_2369),
.B(n_2374),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2376),
.B(n_2379),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2380),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_1924),
.A2(n_2389),
.B(n_2386),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2395),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_2382),
.A2(n_2503),
.B1(n_2003),
.B2(n_2050),
.Y(n_3416)
);

BUFx6f_ASAP7_75t_L g3417 ( 
.A(n_2536),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2396),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2398),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_1924),
.A2(n_2909),
.B(n_2408),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_2231),
.B(n_1912),
.Y(n_3421)
);

NOR2xp33_ASAP7_75t_L g3422 ( 
.A(n_1912),
.B(n_2003),
.Y(n_3422)
);

NOR2xp33_ASAP7_75t_L g3423 ( 
.A(n_1912),
.B(n_2003),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2403),
.B(n_2412),
.Y(n_3424)
);

AND2x6_ASAP7_75t_L g3425 ( 
.A(n_2536),
.B(n_2541),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2413),
.B(n_2414),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_2415),
.B(n_2417),
.Y(n_3427)
);

OAI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_2420),
.A2(n_2423),
.B1(n_2429),
.B2(n_2426),
.Y(n_3428)
);

AO32x2_ASAP7_75t_L g3429 ( 
.A1(n_2039),
.A2(n_2739),
.A3(n_2225),
.B1(n_2052),
.B2(n_2155),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_2430),
.A2(n_2436),
.B(n_2434),
.Y(n_3430)
);

A2O1A1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_2438),
.A2(n_2440),
.B(n_2450),
.C(n_2448),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_2455),
.A2(n_2462),
.B(n_2461),
.Y(n_3432)
);

BUFx3_ASAP7_75t_L g3433 ( 
.A(n_2568),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_2464),
.A2(n_2466),
.B(n_2465),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_L g3435 ( 
.A(n_2050),
.B(n_2094),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_SL g3436 ( 
.A(n_2255),
.B(n_2294),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_2471),
.Y(n_3437)
);

NOR3xp33_ASAP7_75t_L g3438 ( 
.A(n_2329),
.B(n_2245),
.C(n_2217),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_2474),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_2479),
.A2(n_2487),
.B(n_2480),
.Y(n_3440)
);

AOI21x1_ASAP7_75t_L g3441 ( 
.A1(n_2168),
.A2(n_2294),
.B(n_2491),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_2492),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_2495),
.A2(n_2504),
.B(n_2500),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2505),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_2309),
.B(n_2050),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_SL g3446 ( 
.A(n_2096),
.B(n_2109),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_2094),
.B(n_2377),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2506),
.A2(n_2513),
.B(n_2510),
.Y(n_3448)
);

A2O1A1Ixp33_ASAP7_75t_L g3449 ( 
.A1(n_2514),
.A2(n_2517),
.B(n_2521),
.C(n_2515),
.Y(n_3449)
);

BUFx6f_ASAP7_75t_L g3450 ( 
.A(n_2541),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_2522),
.A2(n_2537),
.B(n_2535),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_2538),
.B(n_2540),
.Y(n_3452)
);

INVx4_ASAP7_75t_L g3453 ( 
.A(n_2541),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_2094),
.B(n_2377),
.Y(n_3454)
);

AND2x6_ASAP7_75t_SL g3455 ( 
.A(n_2324),
.B(n_2327),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_2234),
.B(n_2377),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2542),
.B(n_2547),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_2551),
.Y(n_3458)
);

OAI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_2208),
.A2(n_2214),
.B(n_2211),
.Y(n_3459)
);

AND2x4_ASAP7_75t_L g3460 ( 
.A(n_2520),
.B(n_2584),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_2556),
.B(n_2560),
.Y(n_3461)
);

BUFx6f_ASAP7_75t_L g3462 ( 
.A(n_2672),
.Y(n_3462)
);

NOR2x1p5_ASAP7_75t_SL g3463 ( 
.A(n_2215),
.B(n_2219),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2565),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_2567),
.B(n_2569),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2571),
.A2(n_2577),
.B(n_2574),
.Y(n_3466)
);

AOI22x1_ASAP7_75t_L g3467 ( 
.A1(n_2672),
.A2(n_2749),
.B1(n_2384),
.B2(n_2405),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_2580),
.A2(n_2583),
.B(n_2581),
.Y(n_3468)
);

O2A1O1Ixp5_ASAP7_75t_L g3469 ( 
.A1(n_2672),
.A2(n_2749),
.B(n_2586),
.C(n_2587),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_2234),
.B(n_2520),
.Y(n_3470)
);

NAND2xp33_ASAP7_75t_L g3471 ( 
.A(n_2333),
.B(n_2251),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_2585),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_2520),
.B(n_2584),
.Y(n_3473)
);

O2A1O1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_2589),
.A2(n_2595),
.B(n_2598),
.C(n_2592),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_2600),
.A2(n_2611),
.B(n_2606),
.Y(n_3475)
);

BUFx6f_ASAP7_75t_L g3476 ( 
.A(n_2749),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_2584),
.B(n_2675),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2612),
.B(n_2615),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_2621),
.A2(n_2627),
.B(n_2625),
.Y(n_3479)
);

O2A1O1Ixp33_ASAP7_75t_L g3480 ( 
.A1(n_2636),
.A2(n_2640),
.B(n_2641),
.C(n_2637),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_2642),
.B(n_2643),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2645),
.B(n_2648),
.Y(n_3482)
);

O2A1O1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_2649),
.A2(n_2656),
.B(n_2658),
.C(n_2655),
.Y(n_3483)
);

AO21x1_ASAP7_75t_L g3484 ( 
.A1(n_2659),
.A2(n_2668),
.B(n_2665),
.Y(n_3484)
);

INVx1_ASAP7_75t_SL g3485 ( 
.A(n_2243),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_2671),
.B(n_2676),
.Y(n_3486)
);

BUFx12f_ASAP7_75t_L g3487 ( 
.A(n_2109),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_2679),
.B(n_2684),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_2675),
.B(n_2712),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2685),
.A2(n_2689),
.B(n_2687),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_2691),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_2675),
.B(n_2712),
.Y(n_3492)
);

OR2x6_ASAP7_75t_L g3493 ( 
.A(n_1909),
.B(n_2384),
.Y(n_3493)
);

INVx3_ASAP7_75t_L g3494 ( 
.A(n_1909),
.Y(n_3494)
);

AOI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_2692),
.A2(n_2698),
.B(n_2693),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_2712),
.B(n_2718),
.Y(n_3496)
);

INVx3_ASAP7_75t_L g3497 ( 
.A(n_2405),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_2702),
.A2(n_2710),
.B(n_2705),
.Y(n_3498)
);

BUFx2_ASAP7_75t_SL g3499 ( 
.A(n_2039),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2715),
.B(n_2716),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_2717),
.A2(n_2733),
.B(n_2732),
.Y(n_3501)
);

NOR3xp33_ASAP7_75t_L g3502 ( 
.A(n_2247),
.B(n_2333),
.C(n_2328),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_2736),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_2718),
.B(n_2751),
.Y(n_3504)
);

OAI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_2745),
.A2(n_2901),
.B1(n_2837),
.B2(n_2832),
.Y(n_3505)
);

OR2x6_ASAP7_75t_L g3506 ( 
.A(n_2428),
.B(n_2435),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_2753),
.B(n_2755),
.Y(n_3507)
);

NOR2xp33_ASAP7_75t_L g3508 ( 
.A(n_2718),
.B(n_2751),
.Y(n_3508)
);

CKINVDCx8_ASAP7_75t_R g3509 ( 
.A(n_2278),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_2759),
.Y(n_3510)
);

AO21x1_ASAP7_75t_L g3511 ( 
.A1(n_2760),
.A2(n_2769),
.B(n_2762),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2772),
.B(n_2774),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_2775),
.A2(n_2781),
.B(n_2776),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_2782),
.B(n_2783),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2784),
.B(n_2788),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2791),
.B(n_2796),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_2801),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2809),
.B(n_2813),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_2751),
.B(n_2758),
.Y(n_3519)
);

NOR2xp67_ASAP7_75t_L g3520 ( 
.A(n_2222),
.B(n_2223),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_2758),
.B(n_2767),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2815),
.B(n_2821),
.Y(n_3522)
);

NAND3xp33_ASAP7_75t_L g3523 ( 
.A(n_2226),
.B(n_2236),
.C(n_2233),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_2822),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2826),
.B(n_2830),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_2838),
.A2(n_2844),
.B(n_2841),
.Y(n_3526)
);

AND2x2_ASAP7_75t_SL g3527 ( 
.A(n_2324),
.B(n_2758),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_SL g3528 ( 
.A(n_2767),
.B(n_2842),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_SL g3529 ( 
.A(n_2767),
.B(n_2842),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2845),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2859),
.A2(n_2877),
.B(n_2868),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_2884),
.A2(n_2888),
.B(n_2885),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_2892),
.A2(n_2896),
.B(n_2894),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_2898),
.B(n_2243),
.Y(n_3534)
);

A2O1A1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_2241),
.A2(n_2242),
.B(n_2253),
.C(n_2266),
.Y(n_3535)
);

BUFx4f_ASAP7_75t_L g3536 ( 
.A(n_2428),
.Y(n_3536)
);

AND2x4_ASAP7_75t_L g3537 ( 
.A(n_2842),
.B(n_2864),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_2435),
.A2(n_2459),
.B(n_2447),
.Y(n_3538)
);

AND2x6_ASAP7_75t_SL g3539 ( 
.A(n_2324),
.B(n_2327),
.Y(n_3539)
);

OAI21xp33_ASAP7_75t_L g3540 ( 
.A1(n_2254),
.A2(n_2260),
.B(n_2258),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_2259),
.Y(n_3541)
);

OAI21x1_ASAP7_75t_L g3542 ( 
.A1(n_2447),
.A2(n_2906),
.B(n_2469),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_SL g3543 ( 
.A(n_2125),
.B(n_2190),
.Y(n_3543)
);

AOI21x1_ASAP7_75t_L g3544 ( 
.A1(n_2293),
.A2(n_2300),
.B(n_2303),
.Y(n_3544)
);

AOI22x1_ASAP7_75t_L g3545 ( 
.A1(n_2906),
.A2(n_2904),
.B1(n_2459),
.B2(n_2469),
.Y(n_3545)
);

NOR2xp33_ASAP7_75t_L g3546 ( 
.A(n_2864),
.B(n_2865),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_2264),
.B(n_2265),
.Y(n_3547)
);

AOI21x1_ASAP7_75t_L g3548 ( 
.A1(n_2291),
.A2(n_2299),
.B(n_2306),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2497),
.A2(n_2904),
.B(n_2501),
.Y(n_3549)
);

OR2x6_ASAP7_75t_L g3550 ( 
.A(n_2497),
.B(n_2498),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_2254),
.B(n_2260),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_2299),
.B(n_2306),
.Y(n_3552)
);

NOR2x1_ASAP7_75t_L g3553 ( 
.A(n_2568),
.B(n_2639),
.Y(n_3553)
);

OAI321xp33_ASAP7_75t_L g3554 ( 
.A1(n_2280),
.A2(n_2281),
.A3(n_2313),
.B1(n_1985),
.B2(n_2274),
.C(n_2279),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_2864),
.B(n_2865),
.Y(n_3555)
);

A2O1A1Ixp33_ASAP7_75t_L g3556 ( 
.A1(n_2104),
.A2(n_2127),
.B(n_2135),
.C(n_2900),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_2865),
.B(n_2869),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_2104),
.B(n_2127),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_2498),
.A2(n_2501),
.B(n_2771),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_2523),
.Y(n_3560)
);

NOR2xp67_ASAP7_75t_L g3561 ( 
.A(n_1994),
.B(n_2052),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2523),
.A2(n_2824),
.B(n_2766),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_2869),
.B(n_2893),
.Y(n_3563)
);

INVx4_ASAP7_75t_L g3564 ( 
.A(n_2533),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2533),
.A2(n_2764),
.B(n_2804),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_2104),
.B(n_2127),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_2545),
.Y(n_3567)
);

OAI321xp33_ASAP7_75t_L g3568 ( 
.A1(n_2313),
.A2(n_1985),
.A3(n_2297),
.B1(n_2296),
.B2(n_2257),
.C(n_2271),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_2869),
.B(n_2893),
.Y(n_3569)
);

NAND3xp33_ASAP7_75t_SL g3570 ( 
.A(n_2237),
.B(n_2308),
.C(n_2283),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_2545),
.A2(n_2824),
.B(n_2578),
.Y(n_3571)
);

BUFx6f_ASAP7_75t_L g3572 ( 
.A(n_2578),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_2893),
.B(n_2900),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_2579),
.Y(n_3574)
);

OAI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_2332),
.A2(n_2639),
.B1(n_2734),
.B2(n_2875),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_2579),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2900),
.B(n_2613),
.Y(n_3577)
);

O2A1O1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_2193),
.A2(n_2272),
.B(n_2159),
.C(n_2202),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2613),
.A2(n_2878),
.B(n_2646),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_2646),
.B(n_2757),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2757),
.Y(n_3581)
);

BUFx6f_ASAP7_75t_L g3582 ( 
.A(n_2764),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_2766),
.B(n_2771),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_2178),
.B(n_2041),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_2804),
.B(n_2831),
.Y(n_3585)
);

OAI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_2831),
.A2(n_2878),
.B(n_2852),
.Y(n_3586)
);

OAI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_2852),
.A2(n_2135),
.B(n_2251),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_2332),
.Y(n_3588)
);

BUFx2_ASAP7_75t_L g3589 ( 
.A(n_2875),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_2059),
.Y(n_3590)
);

BUFx2_ASAP7_75t_L g3591 ( 
.A(n_2734),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_2178),
.B(n_2041),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_2129),
.A2(n_2150),
.B(n_2151),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_2237),
.A2(n_2337),
.B1(n_2320),
.B2(n_1996),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_2135),
.Y(n_3595)
);

A2O1A1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_1994),
.A2(n_2213),
.B(n_2221),
.C(n_2140),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_2129),
.A2(n_2151),
.B(n_2150),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_2039),
.A2(n_2225),
.B(n_2739),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_2833),
.B(n_2249),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_2833),
.A2(n_2278),
.B1(n_2290),
.B2(n_2221),
.Y(n_3600)
);

NAND2x1p5_ASAP7_75t_L g3601 ( 
.A(n_2225),
.B(n_2739),
.Y(n_3601)
);

NOR2x1_ASAP7_75t_L g3602 ( 
.A(n_2290),
.B(n_2576),
.Y(n_3602)
);

OAI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2257),
.A2(n_2271),
.B(n_2296),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_2059),
.B(n_2224),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_SL g3605 ( 
.A(n_2125),
.B(n_2190),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_2224),
.A2(n_2059),
.B(n_2213),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2059),
.A2(n_2155),
.B(n_2140),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_2152),
.B(n_2337),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_2190),
.B(n_2249),
.Y(n_3609)
);

AOI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_2337),
.A2(n_2320),
.B1(n_2628),
.B2(n_2561),
.Y(n_3610)
);

A2O1A1Ixp33_ASAP7_75t_L g3611 ( 
.A1(n_2336),
.A2(n_2323),
.B(n_2327),
.C(n_2048),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_2297),
.A2(n_2331),
.B(n_2308),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_2283),
.A2(n_2331),
.B1(n_2575),
.B2(n_2743),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_2227),
.B(n_2249),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_2406),
.A2(n_2674),
.B(n_2743),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_2406),
.B(n_2555),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_2453),
.B(n_2575),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2453),
.A2(n_2674),
.B(n_2555),
.Y(n_3618)
);

OAI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_2682),
.A2(n_2713),
.B1(n_2731),
.B2(n_2816),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_2227),
.B(n_2232),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_2561),
.A2(n_2628),
.B1(n_2816),
.B2(n_2232),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2682),
.A2(n_2731),
.B(n_2713),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2227),
.A2(n_2232),
.B(n_2054),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_2009),
.A2(n_2054),
.B(n_1999),
.Y(n_3624)
);

O2A1O1Ixp5_ASAP7_75t_L g3625 ( 
.A1(n_1966),
.A2(n_1999),
.B(n_2000),
.C(n_2082),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_1966),
.A2(n_1999),
.B(n_2000),
.Y(n_3626)
);

INVx2_ASAP7_75t_SL g3627 ( 
.A(n_1966),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_2000),
.Y(n_3628)
);

BUFx8_ASAP7_75t_L g3629 ( 
.A(n_2082),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_2082),
.A2(n_2401),
.B(n_2593),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_SL g3631 ( 
.A(n_2401),
.B(n_2593),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_2401),
.A2(n_2593),
.B(n_2629),
.Y(n_3632)
);

INVx3_ASAP7_75t_L g3633 ( 
.A(n_2629),
.Y(n_3633)
);

AOI22xp5_ASAP7_75t_L g3634 ( 
.A1(n_2629),
.A2(n_2738),
.B1(n_2773),
.B2(n_2780),
.Y(n_3634)
);

OAI21x1_ASAP7_75t_L g3635 ( 
.A1(n_2738),
.A2(n_2773),
.B(n_2780),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_2738),
.A2(n_2773),
.B(n_2780),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_2792),
.A2(n_818),
.B(n_793),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_2792),
.B(n_2866),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_2792),
.Y(n_3639)
);

AOI21x1_ASAP7_75t_L g3640 ( 
.A1(n_2866),
.A2(n_2110),
.B(n_1558),
.Y(n_3640)
);

OAI22xp5_ASAP7_75t_L g3641 ( 
.A1(n_2866),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3641)
);

INVx3_ASAP7_75t_L g3642 ( 
.A(n_2277),
.Y(n_3642)
);

AOI22x1_ASAP7_75t_L g3643 ( 
.A1(n_2388),
.A2(n_2391),
.B1(n_2393),
.B2(n_2390),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3646)
);

AOI21xp5_ASAP7_75t_L g3647 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3647)
);

BUFx2_ASAP7_75t_L g3648 ( 
.A(n_2216),
.Y(n_3648)
);

OAI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3649)
);

AOI22x1_ASAP7_75t_L g3650 ( 
.A1(n_2388),
.A2(n_2391),
.B1(n_2393),
.B2(n_2390),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3651)
);

NAND3xp33_ASAP7_75t_L g3652 ( 
.A(n_2344),
.B(n_793),
.C(n_803),
.Y(n_3652)
);

A2O1A1Ixp33_ASAP7_75t_L g3653 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3653)
);

AOI33xp33_ASAP7_75t_L g3654 ( 
.A1(n_2566),
.A2(n_1677),
.A3(n_1875),
.B1(n_1898),
.B2(n_1650),
.B3(n_2699),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_1957),
.B(n_837),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3656)
);

BUFx3_ASAP7_75t_L g3657 ( 
.A(n_2014),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2212),
.Y(n_3659)
);

NAND2x1_ASAP7_75t_L g3660 ( 
.A(n_2277),
.B(n_1961),
.Y(n_3660)
);

AO21x1_ASAP7_75t_L g3661 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_2212),
.Y(n_3662)
);

BUFx2_ASAP7_75t_L g3663 ( 
.A(n_2216),
.Y(n_3663)
);

AOI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3665)
);

AOI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_2212),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_2014),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_2216),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_2212),
.Y(n_3673)
);

OAI22xp5_ASAP7_75t_L g3674 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3674)
);

INVx2_ASAP7_75t_SL g3675 ( 
.A(n_2277),
.Y(n_3675)
);

A2O1A1Ixp33_ASAP7_75t_L g3676 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3677)
);

OR2x2_ASAP7_75t_L g3678 ( 
.A(n_2908),
.B(n_1970),
.Y(n_3678)
);

OAI22xp5_ASAP7_75t_L g3679 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3679)
);

BUFx2_ASAP7_75t_SL g3680 ( 
.A(n_1967),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3681)
);

CKINVDCx10_ASAP7_75t_R g3682 ( 
.A(n_2075),
.Y(n_3682)
);

INVx3_ASAP7_75t_L g3683 ( 
.A(n_2277),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3685)
);

A2O1A1Ixp33_ASAP7_75t_L g3686 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3686)
);

OAI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3688)
);

AND2x6_ASAP7_75t_SL g3689 ( 
.A(n_2330),
.B(n_837),
.Y(n_3689)
);

O2A1O1Ixp33_ASAP7_75t_SL g3690 ( 
.A1(n_1928),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3690)
);

INVxp67_ASAP7_75t_L g3691 ( 
.A(n_1914),
.Y(n_3691)
);

OAI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_1957),
.B(n_837),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3696)
);

OAI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3697)
);

INVx1_ASAP7_75t_SL g3698 ( 
.A(n_1941),
.Y(n_3698)
);

NOR2x1_ASAP7_75t_L g3699 ( 
.A(n_2185),
.B(n_2301),
.Y(n_3699)
);

INVx2_ASAP7_75t_SL g3700 ( 
.A(n_2277),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_2212),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3702)
);

OR2x6_ASAP7_75t_L g3703 ( 
.A(n_2314),
.B(n_2325),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3704)
);

AOI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3705)
);

A2O1A1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3707)
);

AO22x1_ASAP7_75t_L g3708 ( 
.A1(n_2511),
.A2(n_803),
.B1(n_1049),
.B2(n_1029),
.Y(n_3708)
);

AOI21xp5_ASAP7_75t_L g3709 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3709)
);

AOI221x1_ASAP7_75t_L g3710 ( 
.A1(n_2018),
.A2(n_2025),
.B1(n_1977),
.B2(n_1911),
.C(n_1930),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_R g3711 ( 
.A(n_2197),
.B(n_493),
.Y(n_3711)
);

AND2x4_ASAP7_75t_L g3712 ( 
.A(n_1948),
.B(n_1987),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_2212),
.Y(n_3714)
);

NAND3xp33_ASAP7_75t_SL g3715 ( 
.A(n_2344),
.B(n_793),
.C(n_1255),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_2216),
.Y(n_3716)
);

INVx3_ASAP7_75t_L g3717 ( 
.A(n_2277),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3718)
);

OR2x2_ASAP7_75t_SL g3719 ( 
.A(n_2819),
.B(n_1984),
.Y(n_3719)
);

A2O1A1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3723)
);

OAI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3724)
);

NAND3xp33_ASAP7_75t_L g3725 ( 
.A(n_2344),
.B(n_793),
.C(n_803),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3728)
);

INVxp67_ASAP7_75t_L g3729 ( 
.A(n_1914),
.Y(n_3729)
);

O2A1O1Ixp33_ASAP7_75t_L g3730 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3730)
);

BUFx4f_ASAP7_75t_L g3731 ( 
.A(n_2031),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_2212),
.Y(n_3733)
);

AOI21xp5_ASAP7_75t_L g3734 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_2212),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_L g3736 ( 
.A(n_1957),
.B(n_837),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3737)
);

OAI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3738)
);

OAI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3740)
);

CKINVDCx16_ASAP7_75t_R g3741 ( 
.A(n_2669),
.Y(n_3741)
);

NOR3xp33_ASAP7_75t_L g3742 ( 
.A(n_1950),
.B(n_793),
.C(n_721),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3743)
);

AO21x1_ASAP7_75t_L g3744 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3745)
);

NAND2xp33_ASAP7_75t_L g3746 ( 
.A(n_2669),
.B(n_993),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_SL g3749 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3749)
);

AOI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3752)
);

A2O1A1Ixp33_ASAP7_75t_L g3753 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3755)
);

BUFx12f_ASAP7_75t_L g3756 ( 
.A(n_2305),
.Y(n_3756)
);

HB1xp67_ASAP7_75t_L g3757 ( 
.A(n_2212),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3759)
);

AOI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3760)
);

NOR3xp33_ASAP7_75t_L g3761 ( 
.A(n_1950),
.B(n_793),
.C(n_721),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3764)
);

NOR3xp33_ASAP7_75t_L g3765 ( 
.A(n_1950),
.B(n_793),
.C(n_721),
.Y(n_3765)
);

BUFx8_ASAP7_75t_L g3766 ( 
.A(n_2075),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_2216),
.Y(n_3768)
);

AOI21x1_ASAP7_75t_L g3769 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_SL g3771 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3772)
);

A2O1A1Ixp33_ASAP7_75t_L g3773 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_2212),
.Y(n_3774)
);

O2A1O1Ixp33_ASAP7_75t_L g3775 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3775)
);

NAND3xp33_ASAP7_75t_SL g3776 ( 
.A(n_2344),
.B(n_793),
.C(n_1255),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3777)
);

OAI21xp33_ASAP7_75t_L g3778 ( 
.A1(n_2344),
.A2(n_1029),
.B(n_803),
.Y(n_3778)
);

INVxp67_ASAP7_75t_L g3779 ( 
.A(n_1914),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3780)
);

NAND2x1p5_ASAP7_75t_L g3781 ( 
.A(n_2277),
.B(n_2314),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3782)
);

HB1xp67_ASAP7_75t_L g3783 ( 
.A(n_2212),
.Y(n_3783)
);

BUFx12f_ASAP7_75t_L g3784 ( 
.A(n_2305),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_2216),
.Y(n_3785)
);

AOI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_1957),
.B(n_837),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_1957),
.B(n_837),
.Y(n_3790)
);

AOI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3792)
);

NOR2x1p5_ASAP7_75t_SL g3793 ( 
.A(n_2314),
.B(n_1300),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_2212),
.Y(n_3795)
);

BUFx6f_ASAP7_75t_L g3796 ( 
.A(n_2277),
.Y(n_3796)
);

OAI22xp5_ASAP7_75t_L g3797 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3798)
);

AOI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3801)
);

AOI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3805)
);

AOI21xp33_ASAP7_75t_L g3806 ( 
.A1(n_1928),
.A2(n_793),
.B(n_803),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_2212),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3808)
);

A2O1A1Ixp33_ASAP7_75t_L g3809 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3809)
);

AOI22xp5_ASAP7_75t_L g3810 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3812)
);

CKINVDCx11_ASAP7_75t_R g3813 ( 
.A(n_2009),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_2212),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_2216),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3816)
);

O2A1O1Ixp33_ASAP7_75t_L g3817 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_2212),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3820)
);

OAI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3822)
);

BUFx6f_ASAP7_75t_L g3823 ( 
.A(n_2277),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3824)
);

O2A1O1Ixp33_ASAP7_75t_L g3825 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3825)
);

INVx2_ASAP7_75t_SL g3826 ( 
.A(n_2277),
.Y(n_3826)
);

A2O1A1Ixp33_ASAP7_75t_L g3827 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3829)
);

AO21x2_ASAP7_75t_L g3830 ( 
.A1(n_2409),
.A2(n_2402),
.B(n_2357),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3831)
);

NOR2xp67_ASAP7_75t_SL g3832 ( 
.A(n_1963),
.B(n_2357),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3838)
);

AOI21xp5_ASAP7_75t_L g3839 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3839)
);

OAI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3840)
);

OAI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3843)
);

BUFx6f_ASAP7_75t_L g3844 ( 
.A(n_2277),
.Y(n_3844)
);

OAI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3845)
);

NOR2xp33_ASAP7_75t_L g3846 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3848)
);

AO22x1_ASAP7_75t_L g3849 ( 
.A1(n_2511),
.A2(n_803),
.B1(n_1049),
.B2(n_1029),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_2277),
.Y(n_3851)
);

NOR2xp33_ASAP7_75t_L g3852 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3853)
);

NOR2xp33_ASAP7_75t_L g3854 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3856)
);

A2O1A1Ixp33_ASAP7_75t_L g3857 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3859)
);

BUFx6f_ASAP7_75t_L g3860 ( 
.A(n_2277),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_2216),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3862)
);

AOI22xp5_ASAP7_75t_L g3863 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_SL g3864 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3864)
);

INVx3_ASAP7_75t_L g3865 ( 
.A(n_2277),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3866)
);

NOR2x1_ASAP7_75t_R g3867 ( 
.A(n_2305),
.B(n_493),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_2212),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3871)
);

BUFx6f_ASAP7_75t_L g3872 ( 
.A(n_2277),
.Y(n_3872)
);

CKINVDCx10_ASAP7_75t_R g3873 ( 
.A(n_2075),
.Y(n_3873)
);

A2O1A1Ixp33_ASAP7_75t_L g3874 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_1948),
.B(n_1987),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3877)
);

AOI21x1_ASAP7_75t_L g3878 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3881)
);

O2A1O1Ixp33_ASAP7_75t_L g3882 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3883)
);

INVx1_ASAP7_75t_SL g3884 ( 
.A(n_1941),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_2212),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3887)
);

NAND3xp33_ASAP7_75t_L g3888 ( 
.A(n_2344),
.B(n_793),
.C(n_803),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3890)
);

O2A1O1Ixp33_ASAP7_75t_L g3891 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3892)
);

BUFx6f_ASAP7_75t_L g3893 ( 
.A(n_2277),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3894)
);

INVx2_ASAP7_75t_SL g3895 ( 
.A(n_2277),
.Y(n_3895)
);

A2O1A1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_2216),
.Y(n_3898)
);

INVx11_ASAP7_75t_L g3899 ( 
.A(n_2252),
.Y(n_3899)
);

CKINVDCx16_ASAP7_75t_R g3900 ( 
.A(n_2669),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_2216),
.Y(n_3903)
);

NOR2xp33_ASAP7_75t_L g3904 ( 
.A(n_1957),
.B(n_1945),
.Y(n_3904)
);

NOR2xp67_ASAP7_75t_SL g3905 ( 
.A(n_1963),
.B(n_2357),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3906)
);

AOI21x1_ASAP7_75t_L g3907 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3910)
);

A2O1A1Ixp33_ASAP7_75t_L g3911 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3911)
);

AOI21xp5_ASAP7_75t_L g3912 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3912)
);

A2O1A1Ixp33_ASAP7_75t_L g3913 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3913)
);

BUFx2_ASAP7_75t_L g3914 ( 
.A(n_2216),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_2212),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_1957),
.B(n_837),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_2212),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_2212),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_2212),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_1957),
.B(n_837),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_2212),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_1957),
.B(n_837),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_2216),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_1957),
.B(n_837),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_2819),
.A2(n_2511),
.B1(n_2666),
.B2(n_1932),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_2216),
.Y(n_3939)
);

AND2x4_ASAP7_75t_L g3940 ( 
.A(n_1948),
.B(n_1987),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_2216),
.Y(n_3942)
);

AOI21x1_ASAP7_75t_L g3943 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_SL g3944 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3944)
);

A2O1A1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3946)
);

AOI21x1_ASAP7_75t_L g3947 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3947)
);

AND2x2_ASAP7_75t_L g3948 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3948)
);

OAI21xp33_ASAP7_75t_L g3949 ( 
.A1(n_2344),
.A2(n_1029),
.B(n_803),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_2277),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_2277),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3955)
);

BUFx6f_ASAP7_75t_L g3956 ( 
.A(n_2277),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_2908),
.B(n_1970),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_2216),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_2216),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3962)
);

CKINVDCx10_ASAP7_75t_R g3963 ( 
.A(n_2075),
.Y(n_3963)
);

AOI21x1_ASAP7_75t_L g3964 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3966)
);

AOI21xp5_ASAP7_75t_L g3967 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3967)
);

INVx11_ASAP7_75t_L g3968 ( 
.A(n_2252),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3969)
);

OAI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_3970)
);

AOI22xp33_ASAP7_75t_L g3971 ( 
.A1(n_2819),
.A2(n_2511),
.B1(n_2666),
.B2(n_1932),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3972)
);

O2A1O1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3975)
);

BUFx3_ASAP7_75t_L g3976 ( 
.A(n_2014),
.Y(n_3976)
);

O2A1O1Ixp33_ASAP7_75t_SL g3977 ( 
.A1(n_1928),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3979)
);

AOI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_2388),
.B(n_2390),
.Y(n_3981)
);

BUFx6f_ASAP7_75t_L g3982 ( 
.A(n_2277),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3983)
);

OAI321xp33_ASAP7_75t_L g3984 ( 
.A1(n_2511),
.A2(n_1899),
.A3(n_1835),
.B1(n_1712),
.B2(n_1687),
.C(n_1685),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_SL g3988 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_L g3989 ( 
.A(n_1957),
.B(n_837),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_2277),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_1957),
.B(n_837),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_3993)
);

OAI22xp5_ASAP7_75t_L g3994 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_2023),
.B(n_1278),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_2043),
.B(n_2049),
.Y(n_3996)
);

INVx4_ASAP7_75t_L g3997 ( 
.A(n_1948),
.Y(n_3997)
);

AOI21x1_ASAP7_75t_L g3998 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_3998)
);

NOR3xp33_ASAP7_75t_L g3999 ( 
.A(n_1950),
.B(n_793),
.C(n_721),
.Y(n_3999)
);

O2A1O1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_4000)
);

AOI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4001)
);

OA22x2_ASAP7_75t_L g4002 ( 
.A1(n_2344),
.A2(n_2383),
.B1(n_2445),
.B2(n_2348),
.Y(n_4002)
);

INVxp67_ASAP7_75t_L g4003 ( 
.A(n_1914),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4006)
);

AOI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_1945),
.A2(n_1029),
.B1(n_1049),
.B2(n_803),
.Y(n_4007)
);

NAND3xp33_ASAP7_75t_SL g4008 ( 
.A(n_2344),
.B(n_793),
.C(n_1255),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_2388),
.B(n_2390),
.Y(n_4012)
);

AO21x1_ASAP7_75t_L g4013 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_4013)
);

AOI21x1_ASAP7_75t_L g4014 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_4014)
);

OAI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_4015)
);

OAI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4017)
);

AOI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_2819),
.A2(n_2511),
.B1(n_2666),
.B2(n_1932),
.Y(n_4019)
);

HB1xp67_ASAP7_75t_L g4020 ( 
.A(n_2212),
.Y(n_4020)
);

OAI22x1_ASAP7_75t_L g4021 ( 
.A1(n_2344),
.A2(n_2348),
.B1(n_2445),
.B2(n_2383),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4022)
);

OAI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_2344),
.A2(n_1602),
.B1(n_1716),
.B2(n_1589),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4024)
);

AOI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_SL g4026 ( 
.A1(n_1928),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_2216),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4028)
);

AOI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_1957),
.B(n_837),
.Y(n_4030)
);

AOI21x1_ASAP7_75t_L g4031 ( 
.A1(n_2110),
.A2(n_1558),
.B(n_1248),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_2212),
.Y(n_4033)
);

NAND3xp33_ASAP7_75t_L g4034 ( 
.A(n_2344),
.B(n_793),
.C(n_803),
.Y(n_4034)
);

NOR2xp33_ASAP7_75t_L g4035 ( 
.A(n_1957),
.B(n_837),
.Y(n_4035)
);

OAI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_2023),
.B(n_1278),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4038)
);

A2O1A1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_1957),
.B(n_837),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_2023),
.B(n_1278),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_2212),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4045)
);

A2O1A1Ixp33_ASAP7_75t_L g4046 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_4046)
);

BUFx3_ASAP7_75t_L g4047 ( 
.A(n_2014),
.Y(n_4047)
);

BUFx4f_ASAP7_75t_L g4048 ( 
.A(n_2031),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_1948),
.B(n_1987),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4050)
);

NOR2xp67_ASAP7_75t_L g4051 ( 
.A(n_2156),
.B(n_2229),
.Y(n_4051)
);

A2O1A1Ixp33_ASAP7_75t_L g4052 ( 
.A1(n_2344),
.A2(n_803),
.B(n_1049),
.C(n_1029),
.Y(n_4052)
);

OAI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_2357),
.A2(n_2409),
.B(n_2402),
.Y(n_4053)
);

O2A1O1Ixp33_ASAP7_75t_L g4054 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_4054)
);

O2A1O1Ixp33_ASAP7_75t_L g4055 ( 
.A1(n_2482),
.A2(n_1567),
.B(n_1727),
.C(n_1562),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_2388),
.B(n_2390),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_1957),
.B(n_1945),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4059)
);

INVx3_ASAP7_75t_L g4060 ( 
.A(n_2277),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_2043),
.B(n_2049),
.Y(n_4061)
);

AND2x6_ASAP7_75t_L g4062 ( 
.A(n_2277),
.B(n_1922),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_SL g4063 ( 
.A(n_2023),
.B(n_1278),
.Y(n_4063)
);

AOI21xp5_ASAP7_75t_L g4064 ( 
.A1(n_2357),
.A2(n_818),
.B(n_793),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_2212),
.Y(n_4065)
);

NOR3xp33_ASAP7_75t_SL g4066 ( 
.A(n_3715),
.B(n_4008),
.C(n_3776),
.Y(n_4066)
);

NOR2x1_ASAP7_75t_L g4067 ( 
.A(n_3112),
.B(n_3699),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3742),
.B(n_3761),
.Y(n_4068)
);

OAI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3810),
.A2(n_3705),
.B1(n_3732),
.B2(n_3666),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3197),
.B(n_3236),
.Y(n_4070)
);

AOI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3742),
.A2(n_3765),
.B1(n_3999),
.B2(n_3761),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3072),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_2951),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_2951),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3197),
.B(n_3236),
.Y(n_4075)
);

INVxp67_ASAP7_75t_L g4076 ( 
.A(n_3343),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3863),
.A2(n_3705),
.B1(n_3732),
.B2(n_3666),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3765),
.B(n_3999),
.Y(n_4078)
);

BUFx6f_ASAP7_75t_L g4079 ( 
.A(n_2957),
.Y(n_4079)
);

INVx4_ASAP7_75t_L g4080 ( 
.A(n_3425),
.Y(n_4080)
);

NOR2xp33_ASAP7_75t_L g4081 ( 
.A(n_3760),
.B(n_3810),
.Y(n_4081)
);

BUFx3_ASAP7_75t_L g4082 ( 
.A(n_3509),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_2974),
.Y(n_4083)
);

INVx2_ASAP7_75t_SL g4084 ( 
.A(n_3027),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_2974),
.Y(n_4085)
);

NOR3xp33_ASAP7_75t_SL g4086 ( 
.A(n_3715),
.B(n_4008),
.C(n_3776),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_3863),
.A2(n_3760),
.B1(n_4007),
.B2(n_3706),
.Y(n_4087)
);

AOI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_3646),
.A2(n_3664),
.B(n_3647),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_3094),
.B(n_3116),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_L g4090 ( 
.A1(n_3646),
.A2(n_3664),
.B(n_3647),
.Y(n_4090)
);

CKINVDCx20_ASAP7_75t_R g4091 ( 
.A(n_3340),
.Y(n_4091)
);

BUFx3_ASAP7_75t_L g4092 ( 
.A(n_3509),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_2975),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_2966),
.B(n_2980),
.Y(n_4094)
);

A2O1A1Ixp33_ASAP7_75t_L g4095 ( 
.A1(n_3655),
.A2(n_3736),
.B(n_3788),
.C(n_3694),
.Y(n_4095)
);

BUFx6f_ASAP7_75t_L g4096 ( 
.A(n_2957),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_3425),
.Y(n_4097)
);

AOI21xp5_ASAP7_75t_L g4098 ( 
.A1(n_3667),
.A2(n_3670),
.B(n_3668),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_2975),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_4007),
.B(n_2918),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_SL g4101 ( 
.A(n_2937),
.B(n_3790),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_3667),
.A2(n_3670),
.B(n_3668),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_3677),
.A2(n_3684),
.B(n_3681),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_2966),
.B(n_2980),
.Y(n_4104)
);

HB1xp67_ASAP7_75t_L g4105 ( 
.A(n_3072),
.Y(n_4105)
);

NOR3xp33_ASAP7_75t_SL g4106 ( 
.A(n_3652),
.B(n_3888),
.C(n_3725),
.Y(n_4106)
);

INVx1_ASAP7_75t_SL g4107 ( 
.A(n_3239),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3677),
.A2(n_3684),
.B(n_3681),
.Y(n_4108)
);

NOR3xp33_ASAP7_75t_L g4109 ( 
.A(n_4063),
.B(n_3759),
.C(n_3749),
.Y(n_4109)
);

NOR3xp33_ASAP7_75t_L g4110 ( 
.A(n_3767),
.B(n_3853),
.C(n_3771),
.Y(n_4110)
);

AOI21x1_ASAP7_75t_L g4111 ( 
.A1(n_3832),
.A2(n_3905),
.B(n_3640),
.Y(n_4111)
);

INVx1_ASAP7_75t_SL g4112 ( 
.A(n_3239),
.Y(n_4112)
);

AOI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3693),
.A2(n_3709),
.B(n_3696),
.Y(n_4113)
);

NOR2xp67_ASAP7_75t_SL g4114 ( 
.A(n_3693),
.B(n_3696),
.Y(n_4114)
);

AOI22x1_ASAP7_75t_L g4115 ( 
.A1(n_3709),
.A2(n_3718),
.B1(n_3734),
.B2(n_3723),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_L g4116 ( 
.A1(n_3718),
.A2(n_3734),
.B(n_3723),
.Y(n_4116)
);

OAI21xp33_ASAP7_75t_L g4117 ( 
.A1(n_3653),
.A2(n_3686),
.B(n_3676),
.Y(n_4117)
);

AND2x6_ASAP7_75t_SL g4118 ( 
.A(n_3638),
.B(n_3919),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_R g4119 ( 
.A(n_3007),
.B(n_3741),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_2957),
.Y(n_4120)
);

XNOR2xp5_ASAP7_75t_L g4121 ( 
.A(n_2937),
.B(n_3621),
.Y(n_4121)
);

INVx5_ASAP7_75t_L g4122 ( 
.A(n_3260),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3745),
.A2(n_3750),
.B(n_3748),
.Y(n_4123)
);

BUFx4f_ASAP7_75t_L g4124 ( 
.A(n_2913),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_3255),
.B(n_3278),
.Y(n_4125)
);

OAI22x1_ASAP7_75t_L g4126 ( 
.A1(n_3248),
.A2(n_3387),
.B1(n_3643),
.B2(n_3022),
.Y(n_4126)
);

CKINVDCx5p33_ASAP7_75t_R g4127 ( 
.A(n_3711),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3079),
.B(n_2961),
.Y(n_4128)
);

AOI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_3745),
.A2(n_3750),
.B(n_3748),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_3005),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3009),
.B(n_2911),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3009),
.B(n_2911),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_3924),
.B(n_3926),
.Y(n_4133)
);

NOR2xp33_ASAP7_75t_L g4134 ( 
.A(n_3933),
.B(n_3989),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_3013),
.Y(n_4135)
);

OR2x2_ASAP7_75t_L g4136 ( 
.A(n_3094),
.B(n_3116),
.Y(n_4136)
);

OAI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_3751),
.A2(n_3780),
.B(n_3772),
.Y(n_4137)
);

NOR2xp67_ASAP7_75t_SL g4138 ( 
.A(n_3751),
.B(n_3772),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_2915),
.B(n_2930),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3780),
.A2(n_3786),
.B(n_3782),
.Y(n_4140)
);

AOI22xp5_ASAP7_75t_L g4141 ( 
.A1(n_3992),
.A2(n_4035),
.B1(n_4040),
.B2(n_4030),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_2915),
.B(n_2930),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3013),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_L g4144 ( 
.A(n_2945),
.B(n_3057),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_3637),
.B(n_3038),
.Y(n_4145)
);

A2O1A1Ixp33_ASAP7_75t_L g4146 ( 
.A1(n_3728),
.A2(n_3846),
.B(n_3848),
.C(n_3843),
.Y(n_4146)
);

NOR2xp33_ASAP7_75t_L g4147 ( 
.A(n_3864),
.B(n_3886),
.Y(n_4147)
);

A2O1A1Ixp33_ASAP7_75t_SL g4148 ( 
.A1(n_3728),
.A2(n_3843),
.B(n_3848),
.C(n_3846),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_3637),
.B(n_3038),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_2957),
.Y(n_4150)
);

INVx5_ASAP7_75t_L g4151 ( 
.A(n_3260),
.Y(n_4151)
);

BUFx8_ASAP7_75t_L g4152 ( 
.A(n_2916),
.Y(n_4152)
);

BUFx3_ASAP7_75t_L g4153 ( 
.A(n_3509),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_2931),
.B(n_3644),
.Y(n_4154)
);

NAND2x1p5_ASAP7_75t_L g4155 ( 
.A(n_2959),
.B(n_2987),
.Y(n_4155)
);

O2A1O1Ixp33_ASAP7_75t_L g4156 ( 
.A1(n_3707),
.A2(n_3720),
.B(n_3773),
.C(n_3753),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_SL g4157 ( 
.A(n_3806),
.B(n_3778),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_3652),
.B(n_3725),
.Y(n_4158)
);

INVx3_ASAP7_75t_SL g4159 ( 
.A(n_2994),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_2931),
.B(n_3644),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3658),
.B(n_3665),
.Y(n_4161)
);

AOI22xp5_ASAP7_75t_L g4162 ( 
.A1(n_2914),
.A2(n_2960),
.B1(n_3854),
.B2(n_3852),
.Y(n_4162)
);

AOI21xp5_ASAP7_75t_L g4163 ( 
.A1(n_3782),
.A2(n_3787),
.B(n_3786),
.Y(n_4163)
);

BUFx6f_ASAP7_75t_L g4164 ( 
.A(n_2959),
.Y(n_4164)
);

O2A1O1Ixp33_ASAP7_75t_L g4165 ( 
.A1(n_3809),
.A2(n_3857),
.B(n_3874),
.C(n_3827),
.Y(n_4165)
);

AOI21xp5_ASAP7_75t_L g4166 ( 
.A1(n_3787),
.A2(n_3791),
.B(n_3789),
.Y(n_4166)
);

NOR2xp33_ASAP7_75t_L g4167 ( 
.A(n_3888),
.B(n_4034),
.Y(n_4167)
);

INVx6_ASAP7_75t_L g4168 ( 
.A(n_3049),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3658),
.B(n_3665),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3806),
.B(n_3778),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3685),
.B(n_3688),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_3789),
.A2(n_3794),
.B(n_3791),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3685),
.B(n_3688),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3695),
.B(n_3702),
.Y(n_4174)
);

OAI22xp5_ASAP7_75t_L g4175 ( 
.A1(n_4052),
.A2(n_3911),
.B1(n_3913),
.B2(n_3896),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_3255),
.B(n_3278),
.Y(n_4176)
);

AOI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_3794),
.A2(n_3799),
.B(n_3798),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_3798),
.A2(n_3800),
.B(n_3799),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3695),
.B(n_3702),
.Y(n_4179)
);

NAND2xp33_ASAP7_75t_R g4180 ( 
.A(n_3271),
.B(n_3098),
.Y(n_4180)
);

NOR2xp33_ASAP7_75t_R g4181 ( 
.A(n_3007),
.B(n_3741),
.Y(n_4181)
);

OR2x6_ASAP7_75t_SL g4182 ( 
.A(n_3081),
.B(n_3105),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4039),
.A2(n_3945),
.B1(n_4046),
.B2(n_4034),
.Y(n_4183)
);

O2A1O1Ixp33_ASAP7_75t_L g4184 ( 
.A1(n_3906),
.A2(n_3928),
.B(n_3979),
.C(n_3944),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3713),
.B(n_3721),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_SL g4186 ( 
.A(n_2929),
.B(n_3900),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_3713),
.B(n_3721),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_L g4188 ( 
.A(n_3949),
.B(n_2960),
.Y(n_4188)
);

O2A1O1Ixp5_ASAP7_75t_L g4189 ( 
.A1(n_3708),
.A2(n_3849),
.B(n_3802),
.C(n_3804),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_R g4190 ( 
.A(n_3900),
.B(n_3043),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3722),
.B(n_3737),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3722),
.B(n_3737),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_L g4193 ( 
.A1(n_2914),
.A2(n_4002),
.B1(n_2936),
.B2(n_2927),
.Y(n_4193)
);

NOR2xp67_ASAP7_75t_SL g4194 ( 
.A(n_3800),
.B(n_3802),
.Y(n_4194)
);

INVxp67_ASAP7_75t_L g4195 ( 
.A(n_3343),
.Y(n_4195)
);

O2A1O1Ixp5_ASAP7_75t_SL g4196 ( 
.A1(n_3283),
.A2(n_2917),
.B(n_3995),
.C(n_3988),
.Y(n_4196)
);

OAI22xp5_ASAP7_75t_L g4197 ( 
.A1(n_3935),
.A2(n_4019),
.B1(n_3971),
.B2(n_2962),
.Y(n_4197)
);

A2O1A1Ixp33_ASAP7_75t_L g4198 ( 
.A1(n_3852),
.A2(n_3866),
.B(n_3904),
.C(n_3854),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_3866),
.A2(n_4058),
.B1(n_3904),
.B2(n_2927),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3740),
.B(n_3743),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_SL g4201 ( 
.A(n_3949),
.B(n_2963),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3740),
.B(n_3743),
.Y(n_4202)
);

CKINVDCx5p33_ASAP7_75t_R g4203 ( 
.A(n_3813),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_3804),
.A2(n_3812),
.B(n_3805),
.Y(n_4204)
);

AOI21xp5_ASAP7_75t_L g4205 ( 
.A1(n_3805),
.A2(n_3822),
.B(n_3812),
.Y(n_4205)
);

INVx4_ASAP7_75t_L g4206 ( 
.A(n_3425),
.Y(n_4206)
);

AOI21xp33_ASAP7_75t_L g4207 ( 
.A1(n_2952),
.A2(n_3905),
.B(n_3832),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_SL g4208 ( 
.A(n_2929),
.B(n_3446),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_4058),
.B(n_4037),
.Y(n_4209)
);

O2A1O1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_4042),
.A2(n_2979),
.B(n_3042),
.C(n_2936),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3255),
.B(n_3278),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3747),
.B(n_3752),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3747),
.B(n_3752),
.Y(n_4213)
);

BUFx2_ASAP7_75t_L g4214 ( 
.A(n_3588),
.Y(n_4214)
);

OR2x6_ASAP7_75t_L g4215 ( 
.A(n_3226),
.B(n_3234),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_3822),
.A2(n_3828),
.B(n_3824),
.Y(n_4216)
);

O2A1O1Ixp33_ASAP7_75t_L g4217 ( 
.A1(n_3649),
.A2(n_3674),
.B(n_3692),
.C(n_3679),
.Y(n_4217)
);

BUFx4f_ASAP7_75t_L g4218 ( 
.A(n_2913),
.Y(n_4218)
);

OAI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_2976),
.A2(n_4002),
.B1(n_2910),
.B2(n_2963),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3034),
.B(n_2976),
.Y(n_4220)
);

AOI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_3824),
.A2(n_3831),
.B(n_3828),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3754),
.B(n_3755),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_3831),
.A2(n_3835),
.B(n_3834),
.Y(n_4223)
);

BUFx2_ASAP7_75t_L g4224 ( 
.A(n_3588),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_3754),
.B(n_3755),
.Y(n_4225)
);

BUFx3_ASAP7_75t_L g4226 ( 
.A(n_3049),
.Y(n_4226)
);

OAI22xp5_ASAP7_75t_L g4227 ( 
.A1(n_3935),
.A2(n_4019),
.B1(n_3971),
.B2(n_2955),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3758),
.B(n_3762),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3758),
.B(n_3762),
.Y(n_4229)
);

O2A1O1Ixp33_ASAP7_75t_L g4230 ( 
.A1(n_3649),
.A2(n_3674),
.B(n_3692),
.C(n_3679),
.Y(n_4230)
);

AOI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_3834),
.A2(n_3838),
.B(n_3835),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3034),
.B(n_3120),
.Y(n_4232)
);

BUFx6f_ASAP7_75t_L g4233 ( 
.A(n_2959),
.Y(n_4233)
);

INVx3_ASAP7_75t_L g4234 ( 
.A(n_3238),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_2955),
.A2(n_2962),
.B1(n_3064),
.B2(n_3103),
.Y(n_4235)
);

A2O1A1Ixp33_ASAP7_75t_SL g4236 ( 
.A1(n_3082),
.A2(n_3065),
.B(n_3984),
.C(n_3031),
.Y(n_4236)
);

AOI21xp5_ASAP7_75t_L g4237 ( 
.A1(n_3838),
.A2(n_3850),
.B(n_3839),
.Y(n_4237)
);

AOI21x1_ASAP7_75t_L g4238 ( 
.A1(n_3640),
.A2(n_3878),
.B(n_3769),
.Y(n_4238)
);

BUFx2_ASAP7_75t_L g4239 ( 
.A(n_3588),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_3238),
.Y(n_4240)
);

AOI21xp33_ASAP7_75t_L g4241 ( 
.A1(n_2952),
.A2(n_2972),
.B(n_2932),
.Y(n_4241)
);

O2A1O1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_3697),
.A2(n_3797),
.B(n_3820),
.C(n_3739),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_SL g4243 ( 
.A(n_3120),
.B(n_3208),
.Y(n_4243)
);

OAI21xp5_ASAP7_75t_L g4244 ( 
.A1(n_3839),
.A2(n_3858),
.B(n_3850),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_SL g4245 ( 
.A(n_2910),
.B(n_3053),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_3238),
.B(n_3247),
.Y(n_4246)
);

NOR2xp33_ASAP7_75t_L g4247 ( 
.A(n_3984),
.B(n_3708),
.Y(n_4247)
);

CKINVDCx8_ASAP7_75t_R g4248 ( 
.A(n_3455),
.Y(n_4248)
);

AOI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_3858),
.A2(n_3868),
.B(n_3859),
.Y(n_4249)
);

NAND2x1p5_ASAP7_75t_L g4250 ( 
.A(n_2959),
.B(n_2987),
.Y(n_4250)
);

NOR2xp67_ASAP7_75t_SL g4251 ( 
.A(n_3859),
.B(n_3868),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_R g4252 ( 
.A(n_3043),
.B(n_3327),
.Y(n_4252)
);

O2A1O1Ixp33_ASAP7_75t_L g4253 ( 
.A1(n_3697),
.A2(n_3797),
.B(n_3820),
.C(n_3739),
.Y(n_4253)
);

AOI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_3870),
.A2(n_3875),
.B(n_3871),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_3870),
.A2(n_3875),
.B(n_3871),
.Y(n_4255)
);

OAI22xp5_ASAP7_75t_L g4256 ( 
.A1(n_3064),
.A2(n_3103),
.B1(n_3031),
.B2(n_3821),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_3763),
.B(n_3764),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_SL g4258 ( 
.A(n_3053),
.B(n_3225),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_3877),
.A2(n_3881),
.B(n_3879),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_3821),
.A2(n_3994),
.B1(n_4023),
.B2(n_4010),
.Y(n_4260)
);

O2A1O1Ixp33_ASAP7_75t_L g4261 ( 
.A1(n_3994),
.A2(n_4023),
.B(n_4010),
.C(n_3690),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_3877),
.A2(n_3881),
.B(n_3879),
.Y(n_4262)
);

BUFx6f_ASAP7_75t_L g4263 ( 
.A(n_2987),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3763),
.B(n_3764),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_3264),
.B(n_3266),
.Y(n_4265)
);

O2A1O1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_3977),
.A2(n_4026),
.B(n_2917),
.C(n_2972),
.Y(n_4266)
);

AND2x4_ASAP7_75t_L g4267 ( 
.A(n_3238),
.B(n_3247),
.Y(n_4267)
);

OA22x2_ASAP7_75t_L g4268 ( 
.A1(n_3387),
.A2(n_3335),
.B1(n_4021),
.B2(n_2926),
.Y(n_4268)
);

NOR2xp33_ASAP7_75t_L g4269 ( 
.A(n_3849),
.B(n_4002),
.Y(n_4269)
);

INVx4_ASAP7_75t_L g4270 ( 
.A(n_3425),
.Y(n_4270)
);

OAI21x1_ASAP7_75t_SL g4271 ( 
.A1(n_3180),
.A2(n_3203),
.B(n_3661),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3770),
.B(n_3777),
.Y(n_4272)
);

A2O1A1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4064),
.A2(n_3887),
.B(n_3897),
.C(n_3883),
.Y(n_4273)
);

OAI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_3086),
.A2(n_3083),
.B1(n_4002),
.B2(n_3075),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3770),
.B(n_3777),
.Y(n_4275)
);

INVx5_ASAP7_75t_L g4276 ( 
.A(n_3260),
.Y(n_4276)
);

AOI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_3883),
.A2(n_3897),
.B(n_3887),
.Y(n_4277)
);

INVx3_ASAP7_75t_L g4278 ( 
.A(n_3247),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3801),
.B(n_3803),
.Y(n_4279)
);

AOI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_3901),
.A2(n_3910),
.B(n_3908),
.Y(n_4280)
);

O2A1O1Ixp33_ASAP7_75t_L g4281 ( 
.A1(n_2967),
.A2(n_2953),
.B(n_2932),
.C(n_3901),
.Y(n_4281)
);

NAND3xp33_ASAP7_75t_SL g4282 ( 
.A(n_3910),
.B(n_3916),
.C(n_3912),
.Y(n_4282)
);

O2A1O1Ixp33_ASAP7_75t_L g4283 ( 
.A1(n_2967),
.A2(n_2953),
.B(n_3912),
.C(n_3908),
.Y(n_4283)
);

NOR3xp33_ASAP7_75t_L g4284 ( 
.A(n_3916),
.B(n_3929),
.C(n_3918),
.Y(n_4284)
);

NOR3xp33_ASAP7_75t_SL g4285 ( 
.A(n_3050),
.B(n_3641),
.C(n_3570),
.Y(n_4285)
);

BUFx12f_ASAP7_75t_L g4286 ( 
.A(n_3629),
.Y(n_4286)
);

O2A1O1Ixp33_ASAP7_75t_L g4287 ( 
.A1(n_3918),
.A2(n_3930),
.B(n_3938),
.C(n_3934),
.Y(n_4287)
);

BUFx8_ASAP7_75t_L g4288 ( 
.A(n_2916),
.Y(n_4288)
);

OAI22xp5_ASAP7_75t_L g4289 ( 
.A1(n_3086),
.A2(n_3083),
.B1(n_3075),
.B2(n_2978),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_3801),
.B(n_3803),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_3929),
.A2(n_3934),
.B(n_3930),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3808),
.B(n_3811),
.Y(n_4292)
);

BUFx6f_ASAP7_75t_L g4293 ( 
.A(n_2987),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_3808),
.B(n_3811),
.Y(n_4294)
);

AOI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_3938),
.A2(n_3951),
.B(n_3946),
.Y(n_4295)
);

INVxp67_ASAP7_75t_L g4296 ( 
.A(n_3253),
.Y(n_4296)
);

AOI22xp33_ASAP7_75t_L g4297 ( 
.A1(n_2926),
.A2(n_4021),
.B1(n_3017),
.B2(n_2964),
.Y(n_4297)
);

XNOR2xp5_ASAP7_75t_L g4298 ( 
.A(n_3621),
.B(n_3610),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_SL g4299 ( 
.A(n_3446),
.B(n_3867),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3068),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_L g4301 ( 
.A(n_2973),
.B(n_2981),
.Y(n_4301)
);

A2O1A1Ixp33_ASAP7_75t_L g4302 ( 
.A1(n_3946),
.A2(n_4064),
.B(n_4050),
.C(n_3959),
.Y(n_4302)
);

OAI22xp5_ASAP7_75t_L g4303 ( 
.A1(n_3086),
.A2(n_3051),
.B1(n_3040),
.B2(n_3014),
.Y(n_4303)
);

O2A1O1Ixp5_ASAP7_75t_L g4304 ( 
.A1(n_3951),
.A2(n_3960),
.B(n_3967),
.C(n_3959),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_3816),
.B(n_3819),
.Y(n_4305)
);

A2O1A1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_3960),
.A2(n_3974),
.B(n_3978),
.C(n_3967),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_3816),
.B(n_3819),
.Y(n_4307)
);

NOR2xp33_ASAP7_75t_SL g4308 ( 
.A(n_3867),
.B(n_3487),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_3264),
.B(n_3266),
.Y(n_4309)
);

BUFx2_ASAP7_75t_L g4310 ( 
.A(n_3207),
.Y(n_4310)
);

NOR3xp33_ASAP7_75t_SL g4311 ( 
.A(n_3050),
.B(n_3641),
.C(n_3570),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_L g4312 ( 
.A1(n_3974),
.A2(n_3980),
.B(n_3978),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_3264),
.B(n_3266),
.Y(n_4313)
);

CKINVDCx5p33_ASAP7_75t_R g4314 ( 
.A(n_3327),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_3829),
.B(n_3836),
.Y(n_4315)
);

AOI221xp5_ASAP7_75t_L g4316 ( 
.A1(n_2946),
.A2(n_3687),
.B1(n_3738),
.B2(n_3724),
.C(n_2920),
.Y(n_4316)
);

AOI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_3980),
.A2(n_3993),
.B(n_3983),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3829),
.B(n_3836),
.Y(n_4318)
);

BUFx6f_ASAP7_75t_L g4319 ( 
.A(n_2990),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3672),
.Y(n_4320)
);

AND2x4_ASAP7_75t_L g4321 ( 
.A(n_3247),
.B(n_3213),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_SL g4322 ( 
.A(n_3045),
.B(n_3112),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_SL g4323 ( 
.A(n_3201),
.B(n_2928),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_SL g4324 ( 
.A1(n_2913),
.A2(n_2922),
.B1(n_3643),
.B2(n_3022),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3837),
.B(n_3842),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_3837),
.B(n_3842),
.Y(n_4326)
);

OAI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_2922),
.A2(n_3188),
.B1(n_3146),
.B2(n_2995),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_SL g4328 ( 
.A(n_3201),
.B(n_2928),
.Y(n_4328)
);

NOR2xp33_ASAP7_75t_L g4329 ( 
.A(n_3082),
.B(n_2993),
.Y(n_4329)
);

INVx3_ASAP7_75t_SL g4330 ( 
.A(n_3216),
.Y(n_4330)
);

BUFx2_ASAP7_75t_L g4331 ( 
.A(n_3207),
.Y(n_4331)
);

CKINVDCx20_ASAP7_75t_R g4332 ( 
.A(n_3133),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_3682),
.Y(n_4333)
);

INVx3_ASAP7_75t_SL g4334 ( 
.A(n_3216),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_3983),
.A2(n_4001),
.B(n_3993),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_2993),
.B(n_2995),
.Y(n_4336)
);

NOR2xp33_ASAP7_75t_SL g4337 ( 
.A(n_3487),
.B(n_3049),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3716),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4001),
.A2(n_4006),
.B(n_4004),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3847),
.B(n_3855),
.Y(n_4340)
);

O2A1O1Ixp5_ASAP7_75t_L g4341 ( 
.A1(n_4004),
.A2(n_4009),
.B(n_4011),
.C(n_4006),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3847),
.B(n_3855),
.Y(n_4342)
);

A2O1A1Ixp33_ASAP7_75t_L g4343 ( 
.A1(n_4050),
.A2(n_4009),
.B(n_4017),
.C(n_4011),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_3247),
.B(n_3213),
.Y(n_4344)
);

A2O1A1Ixp33_ASAP7_75t_SL g4345 ( 
.A1(n_3065),
.A2(n_4018),
.B(n_4024),
.C(n_4017),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_3856),
.B(n_3862),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_3037),
.B(n_3048),
.Y(n_4347)
);

AOI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_4018),
.A2(n_4025),
.B(n_4024),
.Y(n_4348)
);

O2A1O1Ixp33_ASAP7_75t_L g4349 ( 
.A1(n_4025),
.A2(n_4029),
.B(n_4032),
.C(n_4028),
.Y(n_4349)
);

BUFx8_ASAP7_75t_L g4350 ( 
.A(n_2916),
.Y(n_4350)
);

NAND2x1p5_ASAP7_75t_L g4351 ( 
.A(n_2990),
.B(n_2992),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_SL g4352 ( 
.A(n_4051),
.B(n_3037),
.Y(n_4352)
);

AOI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_4028),
.A2(n_4032),
.B(n_4029),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_2922),
.A2(n_3048),
.B1(n_3164),
.B2(n_3150),
.Y(n_4354)
);

NAND3xp33_ASAP7_75t_L g4355 ( 
.A(n_4038),
.B(n_4045),
.C(n_4041),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_L g4356 ( 
.A(n_2984),
.B(n_3099),
.Y(n_4356)
);

AOI33xp33_ASAP7_75t_L g4357 ( 
.A1(n_3172),
.A2(n_3332),
.A3(n_3884),
.B1(n_3698),
.B2(n_3241),
.B3(n_3257),
.Y(n_4357)
);

INVxp67_ASAP7_75t_L g4358 ( 
.A(n_3253),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_3768),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_3856),
.B(n_3862),
.Y(n_4360)
);

BUFx3_ASAP7_75t_L g4361 ( 
.A(n_3049),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_3017),
.B(n_3249),
.Y(n_4362)
);

A2O1A1Ixp33_ASAP7_75t_L g4363 ( 
.A1(n_4038),
.A2(n_4041),
.B(n_4045),
.C(n_3654),
.Y(n_4363)
);

OAI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_2935),
.A2(n_2939),
.B(n_2924),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_3880),
.B(n_3889),
.Y(n_4365)
);

O2A1O1Ixp33_ASAP7_75t_L g4366 ( 
.A1(n_3730),
.A2(n_3817),
.B(n_3825),
.C(n_3775),
.Y(n_4366)
);

NOR2xp33_ASAP7_75t_L g4367 ( 
.A(n_3230),
.B(n_2944),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3768),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_3213),
.B(n_2921),
.Y(n_4369)
);

AOI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_2924),
.A2(n_2942),
.B(n_2939),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_SL g4371 ( 
.A(n_4051),
.B(n_3261),
.Y(n_4371)
);

OAI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_3150),
.A2(n_3164),
.B1(n_3161),
.B2(n_2958),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_2926),
.A2(n_4021),
.B1(n_2946),
.B2(n_3661),
.Y(n_4373)
);

HB1xp67_ASAP7_75t_L g4374 ( 
.A(n_3768),
.Y(n_4374)
);

AOI21xp5_ASAP7_75t_L g4375 ( 
.A1(n_2942),
.A2(n_2935),
.B(n_2920),
.Y(n_4375)
);

BUFx6f_ASAP7_75t_SL g4376 ( 
.A(n_3627),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_R g4377 ( 
.A(n_3682),
.B(n_3873),
.Y(n_4377)
);

O2A1O1Ixp33_ASAP7_75t_L g4378 ( 
.A1(n_3730),
.A2(n_3775),
.B(n_3825),
.C(n_3817),
.Y(n_4378)
);

AOI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_3154),
.A2(n_3744),
.B1(n_4013),
.B2(n_3661),
.Y(n_4379)
);

AOI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_3687),
.A2(n_3738),
.B(n_3724),
.Y(n_4380)
);

OR2x6_ASAP7_75t_SL g4381 ( 
.A(n_3081),
.B(n_3105),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_3880),
.B(n_3889),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_3792),
.A2(n_3841),
.B(n_3840),
.Y(n_4383)
);

AOI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_3154),
.A2(n_4013),
.B1(n_3744),
.B2(n_3840),
.Y(n_4384)
);

BUFx4f_ASAP7_75t_SL g4385 ( 
.A(n_3487),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_3892),
.B(n_3894),
.Y(n_4386)
);

AOI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_3792),
.A2(n_3845),
.B(n_3841),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_3892),
.B(n_3894),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_3815),
.Y(n_4389)
);

NOR2x1_ASAP7_75t_L g4390 ( 
.A(n_3699),
.B(n_3104),
.Y(n_4390)
);

AND2x4_ASAP7_75t_L g4391 ( 
.A(n_3213),
.B(n_2921),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_3161),
.A2(n_2958),
.B1(n_2965),
.B2(n_2956),
.Y(n_4392)
);

BUFx6f_ASAP7_75t_L g4393 ( 
.A(n_2990),
.Y(n_4393)
);

O2A1O1Ixp33_ASAP7_75t_L g4394 ( 
.A1(n_3882),
.A2(n_3891),
.B(n_4000),
.C(n_3973),
.Y(n_4394)
);

OAI22xp5_ASAP7_75t_L g4395 ( 
.A1(n_2956),
.A2(n_2968),
.B1(n_2977),
.B2(n_2965),
.Y(n_4395)
);

NOR2xp33_ASAP7_75t_L g4396 ( 
.A(n_2944),
.B(n_3279),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_3785),
.Y(n_4397)
);

BUFx3_ASAP7_75t_L g4398 ( 
.A(n_3049),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_3845),
.A2(n_3970),
.B(n_3955),
.Y(n_4399)
);

BUFx6f_ASAP7_75t_L g4400 ( 
.A(n_2990),
.Y(n_4400)
);

OR2x2_ASAP7_75t_L g4401 ( 
.A(n_3128),
.B(n_3176),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_3902),
.B(n_3909),
.Y(n_4402)
);

OAI22xp5_ASAP7_75t_L g4403 ( 
.A1(n_2968),
.A2(n_2982),
.B1(n_2983),
.B2(n_2977),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3815),
.Y(n_4404)
);

AO32x2_ASAP7_75t_L g4405 ( 
.A1(n_3158),
.A2(n_3575),
.A3(n_3190),
.B1(n_2940),
.B2(n_3169),
.Y(n_4405)
);

O2A1O1Ixp33_ASAP7_75t_L g4406 ( 
.A1(n_3882),
.A2(n_3891),
.B(n_4000),
.C(n_3973),
.Y(n_4406)
);

AOI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_3955),
.A2(n_4015),
.B(n_3970),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_SL g4408 ( 
.A(n_3766),
.B(n_3543),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_SL g4409 ( 
.A(n_3261),
.B(n_3385),
.Y(n_4409)
);

AOI21xp5_ASAP7_75t_L g4410 ( 
.A1(n_4015),
.A2(n_4036),
.B(n_4016),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_4016),
.A2(n_4053),
.B(n_4036),
.Y(n_4411)
);

AOI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4053),
.A2(n_3139),
.B(n_3744),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_3096),
.B(n_3059),
.Y(n_4413)
);

BUFx2_ASAP7_75t_L g4414 ( 
.A(n_3207),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_3139),
.A2(n_4013),
.B(n_2949),
.Y(n_4415)
);

A2O1A1Ixp33_ASAP7_75t_SL g4416 ( 
.A1(n_4054),
.A2(n_4055),
.B(n_3104),
.C(n_3061),
.Y(n_4416)
);

AND2x4_ASAP7_75t_L g4417 ( 
.A(n_3213),
.B(n_2921),
.Y(n_4417)
);

AOI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_2948),
.A2(n_2949),
.B(n_2950),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3861),
.Y(n_4419)
);

A2O1A1Ixp33_ASAP7_75t_SL g4420 ( 
.A1(n_4054),
.A2(n_4055),
.B(n_3061),
.C(n_3568),
.Y(n_4420)
);

O2A1O1Ixp33_ASAP7_75t_L g4421 ( 
.A1(n_3077),
.A2(n_3012),
.B(n_3322),
.C(n_3194),
.Y(n_4421)
);

AOI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_2948),
.A2(n_2950),
.B(n_3830),
.Y(n_4422)
);

BUFx6f_ASAP7_75t_L g4423 ( 
.A(n_2992),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_3830),
.A2(n_3469),
.B(n_3405),
.Y(n_4424)
);

O2A1O1Ixp33_ASAP7_75t_L g4425 ( 
.A1(n_3194),
.A2(n_2970),
.B(n_3356),
.C(n_3172),
.Y(n_4425)
);

INVx3_ASAP7_75t_L g4426 ( 
.A(n_3267),
.Y(n_4426)
);

AOI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_3221),
.A2(n_3279),
.B1(n_3066),
.B2(n_3385),
.Y(n_4427)
);

INVx4_ASAP7_75t_L g4428 ( 
.A(n_3425),
.Y(n_4428)
);

BUFx6f_ASAP7_75t_L g4429 ( 
.A(n_2992),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_3830),
.A2(n_3469),
.B(n_3405),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_3898),
.Y(n_4431)
);

AOI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_3830),
.A2(n_2996),
.B(n_2982),
.Y(n_4432)
);

NOR2xp33_ASAP7_75t_L g4433 ( 
.A(n_3902),
.B(n_3909),
.Y(n_4433)
);

AOI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_3221),
.A2(n_3088),
.B1(n_3335),
.B2(n_3211),
.Y(n_4434)
);

AOI21xp5_ASAP7_75t_L g4435 ( 
.A1(n_2983),
.A2(n_3030),
.B(n_3021),
.Y(n_4435)
);

AO22x1_ASAP7_75t_L g4436 ( 
.A1(n_3766),
.A2(n_3203),
.B1(n_3393),
.B2(n_3180),
.Y(n_4436)
);

INVx3_ASAP7_75t_SL g4437 ( 
.A(n_3216),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_3021),
.A2(n_3125),
.B(n_2996),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_3898),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_3917),
.B(n_3920),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_3917),
.B(n_3920),
.Y(n_4441)
);

AOI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_2999),
.A2(n_3054),
.B(n_3000),
.Y(n_4442)
);

OAI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_2988),
.A2(n_3000),
.B1(n_3026),
.B2(n_2999),
.Y(n_4443)
);

O2A1O1Ixp33_ASAP7_75t_L g4444 ( 
.A1(n_2970),
.A2(n_3356),
.B(n_3268),
.C(n_3265),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3898),
.Y(n_4445)
);

NOR3xp33_ASAP7_75t_SL g4446 ( 
.A(n_3244),
.B(n_3375),
.C(n_3605),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3903),
.Y(n_4447)
);

O2A1O1Ixp33_ASAP7_75t_L g4448 ( 
.A1(n_3158),
.A2(n_3611),
.B(n_2989),
.C(n_3011),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_3931),
.B(n_3936),
.Y(n_4449)
);

AOI22x1_ASAP7_75t_L g4450 ( 
.A1(n_3153),
.A2(n_3147),
.B1(n_3145),
.B2(n_3156),
.Y(n_4450)
);

NAND3xp33_ASAP7_75t_L g4451 ( 
.A(n_3011),
.B(n_3650),
.C(n_3109),
.Y(n_4451)
);

BUFx6f_ASAP7_75t_L g4452 ( 
.A(n_2992),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_3931),
.B(n_3936),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3937),
.B(n_3941),
.Y(n_4454)
);

INVx2_ASAP7_75t_SL g4455 ( 
.A(n_3027),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_3200),
.B(n_3204),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_3937),
.B(n_3941),
.Y(n_4457)
);

AOI21xp5_ASAP7_75t_L g4458 ( 
.A1(n_3089),
.A2(n_3114),
.B(n_3090),
.Y(n_4458)
);

HB1xp67_ASAP7_75t_L g4459 ( 
.A(n_3932),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_3089),
.A2(n_3114),
.B(n_3090),
.Y(n_4460)
);

BUFx3_ASAP7_75t_L g4461 ( 
.A(n_3766),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_3950),
.B(n_3952),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_3950),
.B(n_3952),
.Y(n_4463)
);

INVx1_ASAP7_75t_SL g4464 ( 
.A(n_3256),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_L g4465 ( 
.A1(n_2989),
.A2(n_3257),
.B(n_3285),
.C(n_3241),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_3962),
.B(n_3965),
.Y(n_4466)
);

BUFx6f_ASAP7_75t_L g4467 ( 
.A(n_3100),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_SL g4468 ( 
.A(n_3200),
.B(n_3204),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_SL g4469 ( 
.A(n_2991),
.B(n_3003),
.Y(n_4469)
);

OAI22xp5_ASAP7_75t_L g4470 ( 
.A1(n_2988),
.A2(n_3030),
.B1(n_3033),
.B2(n_3026),
.Y(n_4470)
);

OAI22x1_ASAP7_75t_L g4471 ( 
.A1(n_3248),
.A2(n_3650),
.B1(n_3140),
.B2(n_3142),
.Y(n_4471)
);

OAI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_3033),
.A2(n_3046),
.B1(n_3054),
.B2(n_3036),
.Y(n_4472)
);

O2A1O1Ixp33_ASAP7_75t_L g4473 ( 
.A1(n_3285),
.A2(n_3310),
.B(n_3325),
.C(n_3306),
.Y(n_4473)
);

NOR3xp33_ASAP7_75t_L g4474 ( 
.A(n_3246),
.B(n_3445),
.C(n_3769),
.Y(n_4474)
);

NOR2xp33_ASAP7_75t_L g4475 ( 
.A(n_3962),
.B(n_3965),
.Y(n_4475)
);

A2O1A1Ixp33_ASAP7_75t_SL g4476 ( 
.A1(n_3568),
.A2(n_3554),
.B(n_3109),
.C(n_3603),
.Y(n_4476)
);

O2A1O1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_3403),
.A2(n_3297),
.B(n_3324),
.C(n_3258),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_SL g4478 ( 
.A(n_2991),
.B(n_3003),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_SL g4479 ( 
.A(n_3349),
.B(n_3393),
.Y(n_4479)
);

O2A1O1Ixp33_ASAP7_75t_L g4480 ( 
.A1(n_3283),
.A2(n_3449),
.B(n_3431),
.C(n_3147),
.Y(n_4480)
);

NOR2xp33_ASAP7_75t_L g4481 ( 
.A(n_3966),
.B(n_3969),
.Y(n_4481)
);

OAI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_3036),
.A2(n_3058),
.B1(n_3062),
.B2(n_3046),
.Y(n_4482)
);

OAI22xp5_ASAP7_75t_L g4483 ( 
.A1(n_3058),
.A2(n_3069),
.B1(n_3071),
.B2(n_3062),
.Y(n_4483)
);

AND3x2_ASAP7_75t_L g4484 ( 
.A(n_3543),
.B(n_3638),
.C(n_3603),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_3287),
.B(n_3294),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_3966),
.B(n_3969),
.Y(n_4486)
);

AOI21xp5_ASAP7_75t_L g4487 ( 
.A1(n_3069),
.A2(n_3113),
.B(n_3074),
.Y(n_4487)
);

O2A1O1Ixp33_ASAP7_75t_L g4488 ( 
.A1(n_3153),
.A2(n_3296),
.B(n_3380),
.C(n_3156),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_3113),
.A2(n_3143),
.B(n_3125),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_3186),
.B(n_2912),
.Y(n_4490)
);

AOI22xp33_ASAP7_75t_L g4491 ( 
.A1(n_3159),
.A2(n_3173),
.B1(n_3162),
.B2(n_2912),
.Y(n_4491)
);

O2A1O1Ixp5_ASAP7_75t_SL g4492 ( 
.A1(n_2925),
.A2(n_2934),
.B(n_3659),
.C(n_2941),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_3287),
.B(n_3294),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_3071),
.A2(n_3127),
.B(n_3085),
.Y(n_4494)
);

OAI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_3074),
.A2(n_3085),
.B1(n_3087),
.B2(n_3080),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_3349),
.B(n_3527),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_3873),
.Y(n_4497)
);

AOI21xp5_ASAP7_75t_L g4498 ( 
.A1(n_3119),
.A2(n_3087),
.B(n_3080),
.Y(n_4498)
);

AOI21xp5_ASAP7_75t_L g4499 ( 
.A1(n_3108),
.A2(n_3123),
.B(n_3110),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_3092),
.A2(n_3108),
.B1(n_3110),
.B2(n_3097),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3296),
.A2(n_3380),
.B(n_3145),
.C(n_3179),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_3186),
.B(n_2912),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_3527),
.B(n_3416),
.Y(n_4503)
);

HB1xp67_ASAP7_75t_L g4504 ( 
.A(n_3939),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_SL g4505 ( 
.A(n_3527),
.B(n_3416),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_3972),
.B(n_3975),
.Y(n_4506)
);

NAND2x1_ASAP7_75t_L g4507 ( 
.A(n_3425),
.B(n_3493),
.Y(n_4507)
);

OAI22xp5_ASAP7_75t_L g4508 ( 
.A1(n_3092),
.A2(n_3119),
.B1(n_3122),
.B2(n_3097),
.Y(n_4508)
);

A2O1A1Ixp33_ASAP7_75t_L g4509 ( 
.A1(n_3122),
.A2(n_3127),
.B(n_3137),
.C(n_3123),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3939),
.Y(n_4510)
);

O2A1O1Ixp33_ASAP7_75t_L g4511 ( 
.A1(n_3179),
.A2(n_3168),
.B(n_2919),
.C(n_3020),
.Y(n_4511)
);

INVx3_ASAP7_75t_L g4512 ( 
.A(n_3267),
.Y(n_4512)
);

AOI22xp33_ASAP7_75t_SL g4513 ( 
.A1(n_2954),
.A2(n_2969),
.B1(n_3126),
.B2(n_3091),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_3235),
.B(n_3245),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_L g4515 ( 
.A(n_3972),
.B(n_3975),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_SL g4516 ( 
.A(n_3235),
.B(n_3245),
.Y(n_4516)
);

NOR2xp33_ASAP7_75t_SL g4517 ( 
.A(n_3766),
.B(n_3117),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_SL g4518 ( 
.A(n_3289),
.B(n_3381),
.Y(n_4518)
);

HB1xp67_ASAP7_75t_L g4519 ( 
.A(n_3942),
.Y(n_4519)
);

NAND2x1p5_ASAP7_75t_L g4520 ( 
.A(n_3100),
.B(n_3300),
.Y(n_4520)
);

NAND2xp33_ASAP7_75t_L g4521 ( 
.A(n_3602),
.B(n_3553),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_3958),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_3137),
.A2(n_3143),
.B(n_3138),
.Y(n_4523)
);

NOR2xp67_ASAP7_75t_SL g4524 ( 
.A(n_3212),
.B(n_3117),
.Y(n_4524)
);

NOR3xp33_ASAP7_75t_L g4525 ( 
.A(n_3878),
.B(n_3943),
.C(n_3907),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_SL g4526 ( 
.A(n_3289),
.B(n_3553),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_3138),
.A2(n_3549),
.B(n_3538),
.Y(n_4527)
);

O2A1O1Ixp33_ASAP7_75t_L g4528 ( 
.A1(n_3168),
.A2(n_2919),
.B(n_3020),
.C(n_2971),
.Y(n_4528)
);

AOI21xp5_ASAP7_75t_L g4529 ( 
.A1(n_3538),
.A2(n_3559),
.B(n_3549),
.Y(n_4529)
);

NOR2xp33_ASAP7_75t_R g4530 ( 
.A(n_3963),
.B(n_3746),
.Y(n_4530)
);

AOI22xp33_ASAP7_75t_L g4531 ( 
.A1(n_3159),
.A2(n_3173),
.B1(n_3162),
.B2(n_2969),
.Y(n_4531)
);

O2A1O1Ixp5_ASAP7_75t_L g4532 ( 
.A1(n_3195),
.A2(n_3196),
.B(n_3206),
.C(n_3174),
.Y(n_4532)
);

INVx3_ASAP7_75t_L g4533 ( 
.A(n_3267),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_3963),
.Y(n_4534)
);

A2O1A1Ixp33_ASAP7_75t_L g4535 ( 
.A1(n_3174),
.A2(n_3178),
.B(n_3177),
.C(n_3183),
.Y(n_4535)
);

CKINVDCx5p33_ASAP7_75t_R g4536 ( 
.A(n_3117),
.Y(n_4536)
);

AND3x1_ASAP7_75t_SL g4537 ( 
.A(n_3628),
.B(n_3639),
.C(n_3689),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_3559),
.A2(n_3565),
.B(n_3562),
.Y(n_4538)
);

AOI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_3562),
.A2(n_3571),
.B(n_3565),
.Y(n_4539)
);

AOI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_3211),
.A2(n_3330),
.B1(n_3118),
.B2(n_3275),
.Y(n_4540)
);

AOI22xp33_ASAP7_75t_L g4541 ( 
.A1(n_2954),
.A2(n_3091),
.B1(n_3126),
.B2(n_2969),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_3186),
.B(n_4056),
.Y(n_4542)
);

A2O1A1Ixp33_ASAP7_75t_L g4543 ( 
.A1(n_3178),
.A2(n_3177),
.B(n_3183),
.C(n_3414),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_3985),
.B(n_3986),
.Y(n_4544)
);

BUFx6f_ASAP7_75t_L g4545 ( 
.A(n_3100),
.Y(n_4545)
);

CKINVDCx16_ASAP7_75t_R g4546 ( 
.A(n_3756),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_3961),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3985),
.B(n_3986),
.Y(n_4548)
);

O2A1O1Ixp33_ASAP7_75t_L g4549 ( 
.A1(n_2971),
.A2(n_3691),
.B(n_3729),
.C(n_3141),
.Y(n_4549)
);

BUFx4f_ASAP7_75t_L g4550 ( 
.A(n_3425),
.Y(n_4550)
);

BUFx2_ASAP7_75t_L g4551 ( 
.A(n_3041),
.Y(n_4551)
);

AOI21xp5_ASAP7_75t_L g4552 ( 
.A1(n_3571),
.A2(n_3579),
.B(n_3420),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_3987),
.B(n_3990),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_3987),
.B(n_3990),
.Y(n_4554)
);

AOI22xp33_ASAP7_75t_L g4555 ( 
.A1(n_2954),
.A2(n_3126),
.B1(n_3131),
.B2(n_3091),
.Y(n_4555)
);

AND2x4_ASAP7_75t_L g4556 ( 
.A(n_2921),
.B(n_3039),
.Y(n_4556)
);

BUFx3_ASAP7_75t_L g4557 ( 
.A(n_3766),
.Y(n_4557)
);

INVx2_ASAP7_75t_SL g4558 ( 
.A(n_3027),
.Y(n_4558)
);

NOR3xp33_ASAP7_75t_SL g4559 ( 
.A(n_3609),
.B(n_3631),
.C(n_3613),
.Y(n_4559)
);

O2A1O1Ixp33_ASAP7_75t_L g4560 ( 
.A1(n_3141),
.A2(n_3691),
.B(n_3779),
.C(n_3729),
.Y(n_4560)
);

AOI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_3330),
.A2(n_3383),
.B1(n_3438),
.B2(n_3313),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3996),
.B(n_4005),
.Y(n_4562)
);

BUFx2_ASAP7_75t_L g4563 ( 
.A(n_3041),
.Y(n_4563)
);

O2A1O1Ixp33_ASAP7_75t_L g4564 ( 
.A1(n_3779),
.A2(n_4003),
.B(n_3189),
.C(n_3351),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4056),
.B(n_3131),
.Y(n_4565)
);

AOI22xp33_ASAP7_75t_L g4566 ( 
.A1(n_3131),
.A2(n_3645),
.B1(n_3656),
.B2(n_3651),
.Y(n_4566)
);

INVx5_ASAP7_75t_L g4567 ( 
.A(n_3260),
.Y(n_4567)
);

INVx6_ASAP7_75t_L g4568 ( 
.A(n_3455),
.Y(n_4568)
);

NAND2xp33_ASAP7_75t_L g4569 ( 
.A(n_3602),
.B(n_3438),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3996),
.B(n_4005),
.Y(n_4570)
);

OR2x6_ASAP7_75t_SL g4571 ( 
.A(n_3575),
.B(n_3303),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4022),
.B(n_4044),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_3579),
.A2(n_3420),
.B(n_3414),
.Y(n_4573)
);

A2O1A1Ixp33_ASAP7_75t_L g4574 ( 
.A1(n_3157),
.A2(n_3390),
.B(n_3612),
.C(n_3195),
.Y(n_4574)
);

AOI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_3100),
.A2(n_3731),
.B(n_3300),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_4022),
.B(n_4044),
.Y(n_4576)
);

NOR2xp33_ASAP7_75t_L g4577 ( 
.A(n_3295),
.B(n_3304),
.Y(n_4577)
);

A2O1A1Ixp33_ASAP7_75t_L g4578 ( 
.A1(n_3157),
.A2(n_3390),
.B(n_3612),
.C(n_3196),
.Y(n_4578)
);

AOI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_3678),
.A2(n_3957),
.B1(n_3698),
.B2(n_3884),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_3134),
.A2(n_3144),
.B1(n_3140),
.B2(n_3142),
.Y(n_4580)
);

NOR2xp67_ASAP7_75t_L g4581 ( 
.A(n_2940),
.B(n_3023),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_SL g4582 ( 
.A(n_3556),
.B(n_3212),
.Y(n_4582)
);

NOR2xp33_ASAP7_75t_L g4583 ( 
.A(n_3295),
.B(n_3350),
.Y(n_4583)
);

NOR2xp33_ASAP7_75t_L g4584 ( 
.A(n_3569),
.B(n_3344),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_SL g4585 ( 
.A(n_3212),
.B(n_3198),
.Y(n_4585)
);

OAI22xp5_ASAP7_75t_L g4586 ( 
.A1(n_3134),
.A2(n_3144),
.B1(n_4059),
.B2(n_4057),
.Y(n_4586)
);

AOI21xp5_ASAP7_75t_L g4587 ( 
.A1(n_3300),
.A2(n_4048),
.B(n_3731),
.Y(n_4587)
);

BUFx6f_ASAP7_75t_L g4588 ( 
.A(n_3300),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4027),
.Y(n_4589)
);

A2O1A1Ixp33_ASAP7_75t_SL g4590 ( 
.A1(n_3554),
.A2(n_3586),
.B(n_3205),
.C(n_3587),
.Y(n_4590)
);

AND2x4_ASAP7_75t_SL g4591 ( 
.A(n_3260),
.B(n_2940),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4057),
.B(n_4059),
.Y(n_4592)
);

OAI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_4061),
.A2(n_3256),
.B1(n_3253),
.B2(n_3719),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4061),
.B(n_3678),
.Y(n_4594)
);

AOI21xp5_ASAP7_75t_L g4595 ( 
.A1(n_3731),
.A2(n_4048),
.B(n_3471),
.Y(n_4595)
);

A2O1A1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_3206),
.A2(n_3189),
.B(n_3540),
.C(n_3463),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_2925),
.Y(n_4597)
);

NOR2xp33_ASAP7_75t_L g4598 ( 
.A(n_3198),
.B(n_3678),
.Y(n_4598)
);

BUFx2_ASAP7_75t_L g4599 ( 
.A(n_3648),
.Y(n_4599)
);

O2A1O1Ixp5_ASAP7_75t_SL g4600 ( 
.A1(n_2934),
.A2(n_3659),
.B(n_3662),
.C(n_2941),
.Y(n_4600)
);

AO21x1_ASAP7_75t_L g4601 ( 
.A1(n_3210),
.A2(n_3220),
.B(n_3215),
.Y(n_4601)
);

A2O1A1Ixp33_ASAP7_75t_L g4602 ( 
.A1(n_3540),
.A2(n_3463),
.B(n_3474),
.C(n_3371),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_3957),
.B(n_2985),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_3175),
.Y(n_4604)
);

AOI22xp5_ASAP7_75t_L g4605 ( 
.A1(n_3957),
.A2(n_3502),
.B1(n_3421),
.B2(n_3382),
.Y(n_4605)
);

O2A1O1Ixp33_ASAP7_75t_L g4606 ( 
.A1(n_4003),
.A2(n_3351),
.B(n_3428),
.C(n_3337),
.Y(n_4606)
);

AOI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_3731),
.A2(n_4048),
.B(n_3274),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_2985),
.B(n_3485),
.Y(n_4608)
);

BUFx2_ASAP7_75t_L g4609 ( 
.A(n_3648),
.Y(n_4609)
);

NAND2xp33_ASAP7_75t_SL g4610 ( 
.A(n_3614),
.B(n_3620),
.Y(n_4610)
);

OAI22xp5_ASAP7_75t_L g4611 ( 
.A1(n_3719),
.A2(n_3218),
.B1(n_3332),
.B2(n_3485),
.Y(n_4611)
);

BUFx6f_ASAP7_75t_L g4612 ( 
.A(n_4048),
.Y(n_4612)
);

BUFx2_ASAP7_75t_L g4613 ( 
.A(n_3663),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_L g4614 ( 
.A(n_3558),
.B(n_3566),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_3662),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_3645),
.B(n_3651),
.Y(n_4616)
);

AOI22xp33_ASAP7_75t_SL g4617 ( 
.A1(n_3645),
.A2(n_3656),
.B1(n_3704),
.B2(n_3651),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_3656),
.B(n_3704),
.Y(n_4618)
);

INVx1_ASAP7_75t_SL g4619 ( 
.A(n_3589),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_3669),
.Y(n_4620)
);

AOI22xp33_ASAP7_75t_L g4621 ( 
.A1(n_3704),
.A2(n_3727),
.B1(n_3833),
.B2(n_3726),
.Y(n_4621)
);

BUFx6f_ASAP7_75t_L g4622 ( 
.A(n_3027),
.Y(n_4622)
);

INVxp67_ASAP7_75t_SL g4623 ( 
.A(n_3484),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_3726),
.B(n_3727),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_SL g4625 ( 
.A(n_3382),
.B(n_3395),
.Y(n_4625)
);

O2A1O1Ixp33_ASAP7_75t_L g4626 ( 
.A1(n_3337),
.A2(n_3505),
.B(n_3428),
.C(n_2997),
.Y(n_4626)
);

AOI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_3502),
.A2(n_3421),
.B1(n_3566),
.B2(n_3558),
.Y(n_4627)
);

CKINVDCx20_ASAP7_75t_R g4628 ( 
.A(n_3391),
.Y(n_4628)
);

NAND3xp33_ASAP7_75t_SL g4629 ( 
.A(n_3578),
.B(n_3634),
.C(n_3625),
.Y(n_4629)
);

NOR3xp33_ASAP7_75t_SL g4630 ( 
.A(n_3613),
.B(n_3630),
.C(n_3626),
.Y(n_4630)
);

AOI21xp5_ASAP7_75t_L g4631 ( 
.A1(n_3270),
.A2(n_3276),
.B(n_3274),
.Y(n_4631)
);

OAI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_3218),
.A2(n_2997),
.B1(n_3002),
.B2(n_2986),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_3726),
.B(n_3727),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_L g4634 ( 
.A(n_3280),
.B(n_3551),
.Y(n_4634)
);

OAI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_3907),
.A2(n_3947),
.B(n_3943),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_3669),
.Y(n_4636)
);

O2A1O1Ixp5_ASAP7_75t_L g4637 ( 
.A1(n_3262),
.A2(n_3358),
.B(n_3084),
.C(n_3107),
.Y(n_4637)
);

AOI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_3270),
.A2(n_3282),
.B(n_3276),
.Y(n_4638)
);

A2O1A1Ixp33_ASAP7_75t_L g4639 ( 
.A1(n_3371),
.A2(n_3480),
.B(n_3483),
.C(n_3474),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_3833),
.B(n_3890),
.Y(n_4640)
);

AOI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_3447),
.A2(n_3489),
.B1(n_3496),
.B2(n_3454),
.Y(n_4641)
);

O2A1O1Ixp33_ASAP7_75t_L g4642 ( 
.A1(n_3505),
.A2(n_3002),
.B(n_3015),
.C(n_2986),
.Y(n_4642)
);

CKINVDCx5p33_ASAP7_75t_R g4643 ( 
.A(n_3756),
.Y(n_4643)
);

OAI22xp5_ASAP7_75t_L g4644 ( 
.A1(n_3218),
.A2(n_3015),
.B1(n_3018),
.B2(n_3016),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_2923),
.Y(n_4645)
);

INVx3_ASAP7_75t_L g4646 ( 
.A(n_3703),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_SL g4647 ( 
.A(n_3395),
.B(n_3400),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_3282),
.A2(n_3291),
.B(n_3288),
.Y(n_4648)
);

AOI22xp5_ASAP7_75t_L g4649 ( 
.A1(n_3528),
.A2(n_3557),
.B1(n_3529),
.B2(n_3600),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_3070),
.Y(n_4650)
);

OR2x6_ASAP7_75t_SL g4651 ( 
.A(n_3303),
.B(n_3280),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_L g4652 ( 
.A(n_3833),
.B(n_3890),
.Y(n_4652)
);

INVx4_ASAP7_75t_L g4653 ( 
.A(n_3425),
.Y(n_4653)
);

O2A1O1Ixp33_ASAP7_75t_L g4654 ( 
.A1(n_3016),
.A2(n_3018),
.B(n_3024),
.C(n_3019),
.Y(n_4654)
);

OA22x2_ASAP7_75t_L g4655 ( 
.A1(n_3710),
.A2(n_3242),
.B1(n_3095),
.B2(n_3028),
.Y(n_4655)
);

A2O1A1Ixp33_ASAP7_75t_SL g4656 ( 
.A1(n_3586),
.A2(n_3205),
.B(n_3587),
.C(n_3170),
.Y(n_4656)
);

AND2x6_ASAP7_75t_L g4657 ( 
.A(n_2947),
.B(n_3796),
.Y(n_4657)
);

AOI21xp5_ASAP7_75t_L g4658 ( 
.A1(n_3288),
.A2(n_3299),
.B(n_3291),
.Y(n_4658)
);

AOI22xp5_ASAP7_75t_L g4659 ( 
.A1(n_3600),
.A2(n_3890),
.B1(n_3948),
.B2(n_3927),
.Y(n_4659)
);

AOI21xp5_ASAP7_75t_L g4660 ( 
.A1(n_3299),
.A2(n_3314),
.B(n_3312),
.Y(n_4660)
);

O2A1O1Ixp33_ASAP7_75t_SL g4661 ( 
.A1(n_3596),
.A2(n_3614),
.B(n_3620),
.C(n_3599),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_3312),
.A2(n_3316),
.B(n_3314),
.Y(n_4662)
);

OAI22x1_ASAP7_75t_L g4663 ( 
.A1(n_3052),
.A2(n_3084),
.B1(n_3107),
.B2(n_3398),
.Y(n_4663)
);

NAND3xp33_ASAP7_75t_SL g4664 ( 
.A(n_3578),
.B(n_3634),
.C(n_3625),
.Y(n_4664)
);

BUFx8_ASAP7_75t_L g4665 ( 
.A(n_3756),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_SL g4666 ( 
.A(n_3400),
.B(n_3401),
.Y(n_4666)
);

AOI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_3927),
.A2(n_3948),
.B1(n_4012),
.B2(n_3981),
.Y(n_4667)
);

NOR3xp33_ASAP7_75t_SL g4668 ( 
.A(n_3626),
.B(n_3632),
.C(n_3630),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_3673),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_3927),
.B(n_3948),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_3070),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_3673),
.Y(n_4672)
);

BUFx8_ASAP7_75t_L g4673 ( 
.A(n_3784),
.Y(n_4673)
);

BUFx8_ASAP7_75t_SL g4674 ( 
.A(n_3784),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_L g4675 ( 
.A(n_3981),
.B(n_4012),
.Y(n_4675)
);

BUFx6f_ASAP7_75t_L g4676 ( 
.A(n_3078),
.Y(n_4676)
);

BUFx6f_ASAP7_75t_L g4677 ( 
.A(n_3078),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_3316),
.A2(n_3323),
.B(n_3319),
.Y(n_4678)
);

A2O1A1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_3480),
.A2(n_3483),
.B(n_3024),
.C(n_3029),
.Y(n_4679)
);

O2A1O1Ixp33_ASAP7_75t_L g4680 ( 
.A1(n_3019),
.A2(n_3029),
.B(n_3035),
.C(n_3032),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_3319),
.A2(n_3333),
.B(n_3323),
.Y(n_4681)
);

AOI22xp33_ASAP7_75t_L g4682 ( 
.A1(n_3981),
.A2(n_4056),
.B1(n_4012),
.B2(n_3035),
.Y(n_4682)
);

AOI21xp5_ASAP7_75t_L g4683 ( 
.A1(n_3333),
.A2(n_3352),
.B(n_3345),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_3298),
.B(n_3320),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_3170),
.B(n_3032),
.Y(n_4685)
);

OR2x2_ASAP7_75t_L g4686 ( 
.A(n_3128),
.B(n_3176),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_3701),
.Y(n_4687)
);

NAND3xp33_ASAP7_75t_SL g4688 ( 
.A(n_3624),
.B(n_3636),
.C(n_3632),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_3044),
.B(n_3047),
.Y(n_4689)
);

BUFx10_ASAP7_75t_L g4690 ( 
.A(n_3242),
.Y(n_4690)
);

OAI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_3947),
.A2(n_3998),
.B(n_3964),
.Y(n_4691)
);

O2A1O1Ixp33_ASAP7_75t_L g4692 ( 
.A1(n_3044),
.A2(n_3047),
.B(n_3056),
.C(n_3055),
.Y(n_4692)
);

NOR2xp33_ASAP7_75t_L g4693 ( 
.A(n_3569),
.B(n_3473),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_3701),
.Y(n_4694)
);

NOR2x1_ASAP7_75t_L g4695 ( 
.A(n_3564),
.B(n_3374),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_3714),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_3070),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_3055),
.B(n_3056),
.Y(n_4698)
);

AOI22xp33_ASAP7_75t_L g4699 ( 
.A1(n_3060),
.A2(n_3093),
.B1(n_3101),
.B2(n_3076),
.Y(n_4699)
);

BUFx3_ASAP7_75t_L g4700 ( 
.A(n_3589),
.Y(n_4700)
);

NOR2xp67_ASAP7_75t_L g4701 ( 
.A(n_2940),
.B(n_3023),
.Y(n_4701)
);

OAI22xp5_ASAP7_75t_SL g4702 ( 
.A1(n_3784),
.A2(n_3610),
.B1(n_3689),
.B2(n_3594),
.Y(n_4702)
);

AOI22xp5_ASAP7_75t_L g4703 ( 
.A1(n_3680),
.A2(n_3422),
.B1(n_3435),
.B2(n_3423),
.Y(n_4703)
);

AOI21xp5_ASAP7_75t_L g4704 ( 
.A1(n_3345),
.A2(n_3353),
.B(n_3352),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_3714),
.Y(n_4705)
);

BUFx2_ASAP7_75t_SL g4706 ( 
.A(n_3561),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_3060),
.B(n_3076),
.Y(n_4707)
);

CKINVDCx14_ASAP7_75t_R g4708 ( 
.A(n_3396),
.Y(n_4708)
);

AOI21xp5_ASAP7_75t_L g4709 ( 
.A1(n_3353),
.A2(n_3357),
.B(n_3354),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_3093),
.B(n_3101),
.Y(n_4710)
);

NOR2xp33_ASAP7_75t_L g4711 ( 
.A(n_3551),
.B(n_3595),
.Y(n_4711)
);

NOR2xp33_ASAP7_75t_L g4712 ( 
.A(n_3595),
.B(n_3552),
.Y(n_4712)
);

AOI22xp5_ASAP7_75t_L g4713 ( 
.A1(n_3680),
.A2(n_3422),
.B1(n_3435),
.B2(n_3423),
.Y(n_4713)
);

O2A1O1Ixp33_ASAP7_75t_L g4714 ( 
.A1(n_3115),
.A2(n_3124),
.B(n_3129),
.C(n_3121),
.Y(n_4714)
);

AO32x1_ASAP7_75t_L g4715 ( 
.A1(n_3229),
.A2(n_3272),
.A3(n_3191),
.B1(n_3228),
.B2(n_3199),
.Y(n_4715)
);

INVx2_ASAP7_75t_SL g4716 ( 
.A(n_3078),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_3595),
.B(n_3552),
.Y(n_4717)
);

OAI22xp5_ASAP7_75t_L g4718 ( 
.A1(n_3115),
.A2(n_3121),
.B1(n_3129),
.B2(n_3124),
.Y(n_4718)
);

NOR2xp33_ASAP7_75t_L g4719 ( 
.A(n_3148),
.B(n_3149),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_3354),
.A2(n_3360),
.B(n_3357),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_3148),
.B(n_3149),
.Y(n_4721)
);

OAI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_3151),
.A2(n_3152),
.B1(n_3160),
.B2(n_3155),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_3735),
.Y(n_4723)
);

O2A1O1Ixp33_ASAP7_75t_L g4724 ( 
.A1(n_3151),
.A2(n_3155),
.B(n_3160),
.C(n_3152),
.Y(n_4724)
);

A2O1A1Ixp33_ASAP7_75t_L g4725 ( 
.A1(n_3171),
.A2(n_3262),
.B(n_3378),
.C(n_3102),
.Y(n_4725)
);

A2O1A1Ixp33_ASAP7_75t_SL g4726 ( 
.A1(n_3378),
.A2(n_3494),
.B(n_3497),
.C(n_2998),
.Y(n_4726)
);

OAI21xp33_ASAP7_75t_SL g4727 ( 
.A1(n_3028),
.A2(n_3095),
.B(n_3355),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_SL g4728 ( 
.A(n_3401),
.B(n_3577),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_3774),
.Y(n_4729)
);

A2O1A1Ixp33_ASAP7_75t_L g4730 ( 
.A1(n_3171),
.A2(n_3102),
.B(n_3536),
.C(n_3227),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_3166),
.B(n_3001),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_3070),
.Y(n_4732)
);

AOI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_3360),
.A2(n_3367),
.B(n_3365),
.Y(n_4733)
);

AOI21xp5_ASAP7_75t_L g4734 ( 
.A1(n_3365),
.A2(n_3367),
.B(n_3536),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_SL g4735 ( 
.A(n_3577),
.B(n_3460),
.Y(n_4735)
);

A2O1A1Ixp33_ASAP7_75t_L g4736 ( 
.A1(n_3536),
.A2(n_3227),
.B(n_3432),
.C(n_3430),
.Y(n_4736)
);

BUFx6f_ASAP7_75t_L g4737 ( 
.A(n_3078),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_3166),
.B(n_3001),
.Y(n_4738)
);

AOI22xp5_ASAP7_75t_L g4739 ( 
.A1(n_3519),
.A2(n_3546),
.B1(n_3521),
.B2(n_3627),
.Y(n_4739)
);

AOI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_3536),
.A2(n_3355),
.B(n_3269),
.Y(n_4740)
);

O2A1O1Ixp33_ASAP7_75t_L g4741 ( 
.A1(n_3362),
.A2(n_3535),
.B(n_3534),
.C(n_3331),
.Y(n_4741)
);

A2O1A1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_3430),
.A2(n_3434),
.B(n_3440),
.C(n_3432),
.Y(n_4742)
);

OAI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_3394),
.A2(n_3507),
.B1(n_3166),
.B2(n_3398),
.Y(n_4743)
);

AOI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_3269),
.A2(n_3467),
.B(n_3292),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_3441),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_3001),
.B(n_3418),
.Y(n_4746)
);

NOR2xp33_ASAP7_75t_L g4747 ( 
.A(n_3388),
.B(n_3436),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_3467),
.A2(n_3292),
.B(n_3281),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_3001),
.B(n_3418),
.Y(n_4749)
);

AOI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_3281),
.A2(n_3453),
.B(n_3386),
.Y(n_4750)
);

NOR2xp33_ASAP7_75t_L g4751 ( 
.A(n_3534),
.B(n_3608),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_3386),
.A2(n_3453),
.B(n_3710),
.Y(n_4752)
);

AOI21xp5_ASAP7_75t_L g4753 ( 
.A1(n_3386),
.A2(n_3453),
.B(n_3493),
.Y(n_4753)
);

AOI22xp5_ASAP7_75t_L g4754 ( 
.A1(n_3519),
.A2(n_3546),
.B1(n_3521),
.B2(n_3627),
.Y(n_4754)
);

OR2x2_ASAP7_75t_L g4755 ( 
.A(n_3217),
.B(n_3224),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_SL g4756 ( 
.A(n_3460),
.B(n_3537),
.Y(n_4756)
);

O2A1O1Ixp33_ASAP7_75t_L g4757 ( 
.A1(n_3331),
.A2(n_3334),
.B(n_3338),
.C(n_3336),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_3418),
.B(n_3437),
.Y(n_4758)
);

BUFx3_ASAP7_75t_L g4759 ( 
.A(n_3591),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_3774),
.Y(n_4760)
);

NAND2x1p5_ASAP7_75t_L g4761 ( 
.A(n_2940),
.B(n_3023),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_R g4762 ( 
.A(n_3629),
.B(n_3539),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_3795),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_3252),
.B(n_3181),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_3795),
.Y(n_4765)
);

NOR2xp33_ASAP7_75t_L g4766 ( 
.A(n_3608),
.B(n_3591),
.Y(n_4766)
);

AOI21xp5_ASAP7_75t_L g4767 ( 
.A1(n_3386),
.A2(n_3453),
.B(n_3493),
.Y(n_4767)
);

NOR3xp33_ASAP7_75t_SL g4768 ( 
.A(n_3636),
.B(n_3623),
.C(n_3624),
.Y(n_4768)
);

AOI22xp5_ASAP7_75t_L g4769 ( 
.A1(n_3477),
.A2(n_3504),
.B1(n_3508),
.B2(n_3492),
.Y(n_4769)
);

OR2x6_ASAP7_75t_L g4770 ( 
.A(n_3222),
.B(n_3023),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_3217),
.B(n_3224),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_R g4772 ( 
.A(n_3629),
.B(n_3539),
.Y(n_4772)
);

NAND3xp33_ASAP7_75t_SL g4773 ( 
.A(n_3615),
.B(n_3622),
.C(n_3618),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_3619),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_SL g4775 ( 
.A(n_3460),
.B(n_3537),
.Y(n_4775)
);

INVx3_ASAP7_75t_L g4776 ( 
.A(n_3703),
.Y(n_4776)
);

A2O1A1Ixp33_ASAP7_75t_L g4777 ( 
.A1(n_3434),
.A2(n_3443),
.B(n_3448),
.C(n_3440),
.Y(n_4777)
);

AOI21x1_ASAP7_75t_L g4778 ( 
.A1(n_3964),
.A2(n_4014),
.B(n_3998),
.Y(n_4778)
);

AOI221xp5_ASAP7_75t_L g4779 ( 
.A1(n_3233),
.A2(n_3263),
.B1(n_3254),
.B2(n_3250),
.C(n_3215),
.Y(n_4779)
);

OAI22xp5_ASAP7_75t_L g4780 ( 
.A1(n_3394),
.A2(n_3507),
.B1(n_3336),
.B2(n_3338),
.Y(n_4780)
);

BUFx2_ASAP7_75t_L g4781 ( 
.A(n_3914),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_3252),
.B(n_3181),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_3442),
.B(n_3458),
.Y(n_4783)
);

CKINVDCx20_ASAP7_75t_R g4784 ( 
.A(n_3629),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_3807),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_SL g4786 ( 
.A(n_3460),
.B(n_3537),
.Y(n_4786)
);

AND2x6_ASAP7_75t_L g4787 ( 
.A(n_2947),
.B(n_3796),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_SL g4788 ( 
.A(n_3460),
.B(n_3537),
.Y(n_4788)
);

OR2x2_ASAP7_75t_L g4789 ( 
.A(n_3233),
.B(n_3250),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_3458),
.B(n_3472),
.Y(n_4790)
);

AOI22xp5_ASAP7_75t_L g4791 ( 
.A1(n_3573),
.A2(n_3231),
.B1(n_3537),
.B2(n_3520),
.Y(n_4791)
);

BUFx8_ASAP7_75t_SL g4792 ( 
.A(n_3633),
.Y(n_4792)
);

CKINVDCx20_ASAP7_75t_R g4793 ( 
.A(n_3629),
.Y(n_4793)
);

AOI22xp33_ASAP7_75t_L g4794 ( 
.A1(n_3252),
.A2(n_3404),
.B1(n_3481),
.B2(n_3452),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_SL g4795 ( 
.A(n_3520),
.B(n_3561),
.Y(n_4795)
);

AOI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_3386),
.A2(n_3453),
.B(n_3493),
.Y(n_4796)
);

AOI21xp5_ASAP7_75t_L g4797 ( 
.A1(n_3493),
.A2(n_3550),
.B(n_3506),
.Y(n_4797)
);

A2O1A1Ixp33_ASAP7_75t_L g4798 ( 
.A1(n_3443),
.A2(n_3451),
.B(n_3466),
.C(n_3448),
.Y(n_4798)
);

OR2x6_ASAP7_75t_SL g4799 ( 
.A(n_3130),
.B(n_3163),
.Y(n_4799)
);

NOR2xp33_ASAP7_75t_L g4800 ( 
.A(n_3397),
.B(n_3616),
.Y(n_4800)
);

BUFx3_ASAP7_75t_L g4801 ( 
.A(n_2933),
.Y(n_4801)
);

NOR2xp33_ASAP7_75t_L g4802 ( 
.A(n_3616),
.B(n_3617),
.Y(n_4802)
);

NOR3xp33_ASAP7_75t_SL g4803 ( 
.A(n_3623),
.B(n_3619),
.C(n_3618),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_3458),
.B(n_3472),
.Y(n_4804)
);

NOR2xp33_ASAP7_75t_R g4805 ( 
.A(n_3293),
.B(n_3317),
.Y(n_4805)
);

AOI21xp5_ASAP7_75t_L g4806 ( 
.A1(n_3506),
.A2(n_3550),
.B(n_3302),
.Y(n_4806)
);

INVx1_ASAP7_75t_SL g4807 ( 
.A(n_3394),
.Y(n_4807)
);

NOR2xp33_ASAP7_75t_L g4808 ( 
.A(n_3617),
.B(n_3456),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_3807),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_R g4810 ( 
.A(n_3216),
.B(n_3633),
.Y(n_4810)
);

OAI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4014),
.A2(n_4031),
.B(n_3523),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_3342),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_3814),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_3814),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_3472),
.B(n_3510),
.Y(n_4815)
);

AOI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_3506),
.A2(n_3550),
.B(n_3302),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_3228),
.B(n_3028),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_3342),
.Y(n_4818)
);

OAI22x1_ASAP7_75t_L g4819 ( 
.A1(n_3052),
.A2(n_3358),
.B1(n_3307),
.B2(n_3366),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_3510),
.B(n_3517),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_3818),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_3510),
.B(n_3517),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_3818),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_3517),
.B(n_3326),
.Y(n_4824)
);

O2A1O1Ixp33_ASAP7_75t_SL g4825 ( 
.A1(n_3628),
.A2(n_3639),
.B(n_3622),
.C(n_3615),
.Y(n_4825)
);

NOR2xp33_ASAP7_75t_L g4826 ( 
.A(n_3470),
.B(n_3555),
.Y(n_4826)
);

BUFx12f_ASAP7_75t_L g4827 ( 
.A(n_3216),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_SL g4828 ( 
.A(n_3374),
.B(n_3523),
.Y(n_4828)
);

AOI22xp5_ASAP7_75t_L g4829 ( 
.A1(n_3231),
.A2(n_3633),
.B1(n_3563),
.B2(n_3555),
.Y(n_4829)
);

INVx3_ASAP7_75t_L g4830 ( 
.A(n_3703),
.Y(n_4830)
);

OAI22x1_ASAP7_75t_L g4831 ( 
.A1(n_3307),
.A2(n_3389),
.B1(n_3366),
.B2(n_3290),
.Y(n_4831)
);

AOI22xp5_ASAP7_75t_L g4832 ( 
.A1(n_3633),
.A2(n_3563),
.B1(n_3555),
.B2(n_3594),
.Y(n_4832)
);

AOI21xp5_ASAP7_75t_L g4833 ( 
.A1(n_3506),
.A2(n_3550),
.B(n_3301),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_SL g4834 ( 
.A1(n_3494),
.A2(n_3497),
.B(n_3642),
.C(n_2998),
.Y(n_4834)
);

AOI21xp5_ASAP7_75t_L g4835 ( 
.A1(n_3506),
.A2(n_3550),
.B(n_3301),
.Y(n_4835)
);

AOI21xp5_ASAP7_75t_L g4836 ( 
.A1(n_3550),
.A2(n_3466),
.B(n_3451),
.Y(n_4836)
);

NOR3xp33_ASAP7_75t_SL g4837 ( 
.A(n_3584),
.B(n_3592),
.C(n_3607),
.Y(n_4837)
);

BUFx3_ASAP7_75t_L g4838 ( 
.A(n_2933),
.Y(n_4838)
);

O2A1O1Ixp33_ASAP7_75t_SL g4839 ( 
.A1(n_3580),
.A2(n_3585),
.B(n_3583),
.C(n_3660),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_3028),
.B(n_3095),
.Y(n_4840)
);

A2O1A1Ixp33_ASAP7_75t_L g4841 ( 
.A1(n_3468),
.A2(n_3479),
.B(n_3490),
.C(n_3475),
.Y(n_4841)
);

NOR2xp33_ASAP7_75t_R g4842 ( 
.A(n_2933),
.B(n_2943),
.Y(n_4842)
);

AOI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_3563),
.A2(n_3452),
.B1(n_3481),
.B2(n_3404),
.Y(n_4843)
);

INVxp67_ASAP7_75t_L g4844 ( 
.A(n_3404),
.Y(n_4844)
);

OR2x6_ASAP7_75t_L g4845 ( 
.A(n_3222),
.B(n_3136),
.Y(n_4845)
);

OAI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_3073),
.A2(n_3475),
.B(n_3468),
.Y(n_4846)
);

AOI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_3479),
.A2(n_3495),
.B(n_3490),
.Y(n_4847)
);

AOI21xp5_ASAP7_75t_L g4848 ( 
.A1(n_3495),
.A2(n_3501),
.B(n_3498),
.Y(n_4848)
);

O2A1O1Ixp33_ASAP7_75t_SL g4849 ( 
.A1(n_3580),
.A2(n_3585),
.B(n_3583),
.C(n_3660),
.Y(n_4849)
);

NOR2xp33_ASAP7_75t_SL g4850 ( 
.A(n_3564),
.B(n_2943),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_SL g4851 ( 
.A(n_3459),
.B(n_2943),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_3869),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_3498),
.A2(n_3513),
.B(n_3501),
.Y(n_4853)
);

CKINVDCx5p33_ASAP7_75t_R g4854 ( 
.A(n_3342),
.Y(n_4854)
);

OAI22xp5_ASAP7_75t_SL g4855 ( 
.A1(n_3222),
.A2(n_3095),
.B1(n_3389),
.B2(n_3025),
.Y(n_4855)
);

NOR2xp33_ASAP7_75t_L g4856 ( 
.A(n_3025),
.B(n_3547),
.Y(n_4856)
);

NOR2xp33_ASAP7_75t_L g4857 ( 
.A(n_3025),
.B(n_3547),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_3326),
.B(n_3328),
.Y(n_4858)
);

CKINVDCx20_ASAP7_75t_R g4859 ( 
.A(n_3010),
.Y(n_4859)
);

AOI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_3452),
.A2(n_3514),
.B1(n_3481),
.B2(n_3346),
.Y(n_4860)
);

OAI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_3507),
.A2(n_3334),
.B1(n_3347),
.B2(n_3339),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_3328),
.B(n_3346),
.Y(n_4862)
);

AOI22xp33_ASAP7_75t_L g4863 ( 
.A1(n_3514),
.A2(n_3222),
.B1(n_3370),
.B2(n_3368),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_3869),
.Y(n_4864)
);

AOI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_3513),
.A2(n_3531),
.B(n_3526),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_3368),
.B(n_3370),
.Y(n_4866)
);

AOI221xp5_ASAP7_75t_L g4867 ( 
.A1(n_3254),
.A2(n_3263),
.B1(n_3223),
.B2(n_3251),
.C(n_3237),
.Y(n_4867)
);

AOI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_3526),
.A2(n_3532),
.B(n_3531),
.Y(n_4868)
);

OAI22xp5_ASAP7_75t_L g4869 ( 
.A1(n_3339),
.A2(n_3364),
.B1(n_3369),
.B2(n_3347),
.Y(n_4869)
);

BUFx6f_ASAP7_75t_L g4870 ( 
.A(n_3106),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_SL g4871 ( 
.A(n_3459),
.B(n_3010),
.Y(n_4871)
);

OAI22xp5_ASAP7_75t_L g4872 ( 
.A1(n_3364),
.A2(n_3373),
.B1(n_3376),
.B2(n_3369),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_L g4873 ( 
.A(n_3025),
.B(n_3547),
.Y(n_4873)
);

BUFx2_ASAP7_75t_L g4874 ( 
.A(n_3305),
.Y(n_4874)
);

NOR2xp33_ASAP7_75t_L g4875 ( 
.A(n_3010),
.B(n_3063),
.Y(n_4875)
);

INVx5_ASAP7_75t_L g4876 ( 
.A(n_4062),
.Y(n_4876)
);

AOI21x1_ASAP7_75t_L g4877 ( 
.A1(n_3273),
.A2(n_3548),
.B(n_3220),
.Y(n_4877)
);

AOI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_3514),
.A2(n_3464),
.B1(n_3444),
.B2(n_3439),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_3384),
.B(n_3407),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_3384),
.B(n_3407),
.Y(n_4880)
);

NOR2xp33_ASAP7_75t_R g4881 ( 
.A(n_3063),
.B(n_3132),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_3410),
.B(n_3413),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_3410),
.B(n_3413),
.Y(n_4883)
);

INVxp67_ASAP7_75t_L g4884 ( 
.A(n_3373),
.Y(n_4884)
);

AOI21xp5_ASAP7_75t_L g4885 ( 
.A1(n_3532),
.A2(n_3533),
.B(n_3309),
.Y(n_4885)
);

NAND3xp33_ASAP7_75t_SL g4886 ( 
.A(n_3533),
.B(n_3511),
.C(n_3484),
.Y(n_4886)
);

AOI22xp5_ASAP7_75t_L g4887 ( 
.A1(n_3415),
.A2(n_3464),
.B1(n_3444),
.B2(n_3439),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_SL g4888 ( 
.A(n_3063),
.B(n_3132),
.Y(n_4888)
);

AOI21xp5_ASAP7_75t_L g4889 ( 
.A1(n_3309),
.A2(n_3545),
.B(n_3542),
.Y(n_4889)
);

A2O1A1Ixp33_ASAP7_75t_L g4890 ( 
.A1(n_3210),
.A2(n_3251),
.B(n_3223),
.C(n_3237),
.Y(n_4890)
);

O2A1O1Ixp33_ASAP7_75t_L g4891 ( 
.A1(n_3376),
.A2(n_3488),
.B(n_3399),
.C(n_3402),
.Y(n_4891)
);

NOR2xp33_ASAP7_75t_L g4892 ( 
.A(n_3132),
.B(n_3232),
.Y(n_4892)
);

NOR2xp33_ASAP7_75t_R g4893 ( 
.A(n_3232),
.B(n_3433),
.Y(n_4893)
);

AND2x4_ASAP7_75t_L g4894 ( 
.A(n_3165),
.B(n_3712),
.Y(n_4894)
);

AOI21xp5_ASAP7_75t_L g4895 ( 
.A1(n_3545),
.A2(n_3542),
.B(n_3277),
.Y(n_4895)
);

BUFx3_ASAP7_75t_L g4896 ( 
.A(n_3232),
.Y(n_4896)
);

OAI21xp33_ASAP7_75t_SL g4897 ( 
.A1(n_3318),
.A2(n_3321),
.B(n_3542),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_3885),
.B(n_3915),
.Y(n_4898)
);

AOI21xp5_ASAP7_75t_L g4899 ( 
.A1(n_3277),
.A2(n_3392),
.B(n_3111),
.Y(n_4899)
);

A2O1A1Ixp33_ASAP7_75t_L g4900 ( 
.A1(n_3607),
.A2(n_3976),
.B(n_3433),
.C(n_4047),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_3415),
.B(n_3419),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_3419),
.B(n_3491),
.Y(n_4902)
);

NOR2xp33_ASAP7_75t_L g4903 ( 
.A(n_3433),
.B(n_3657),
.Y(n_4903)
);

BUFx3_ASAP7_75t_L g4904 ( 
.A(n_3657),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_3922),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_3657),
.B(n_3671),
.Y(n_4906)
);

BUFx3_ASAP7_75t_L g4907 ( 
.A(n_3671),
.Y(n_4907)
);

OAI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_3111),
.A2(n_3548),
.B(n_3922),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_3923),
.B(n_3925),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_3923),
.B(n_3925),
.Y(n_4910)
);

AO21x2_ASAP7_75t_L g4911 ( 
.A1(n_3273),
.A2(n_3511),
.B(n_3484),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_SL g4912 ( 
.A(n_3671),
.B(n_3976),
.Y(n_4912)
);

BUFx8_ASAP7_75t_L g4913 ( 
.A(n_3429),
.Y(n_4913)
);

OAI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_3399),
.A2(n_3518),
.B1(n_3402),
.B2(n_3406),
.Y(n_4914)
);

BUFx6f_ASAP7_75t_L g4915 ( 
.A(n_3106),
.Y(n_4915)
);

AOI21xp5_ASAP7_75t_L g4916 ( 
.A1(n_3277),
.A2(n_3392),
.B(n_3111),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4033),
.Y(n_4917)
);

BUFx12f_ASAP7_75t_L g4918 ( 
.A(n_3590),
.Y(n_4918)
);

AOI22xp5_ASAP7_75t_L g4919 ( 
.A1(n_3491),
.A2(n_3530),
.B1(n_3524),
.B2(n_3503),
.Y(n_4919)
);

OAI22xp5_ASAP7_75t_L g4920 ( 
.A1(n_3406),
.A2(n_3500),
.B1(n_3409),
.B2(n_3411),
.Y(n_4920)
);

NOR3xp33_ASAP7_75t_L g4921 ( 
.A(n_3635),
.B(n_3169),
.C(n_3136),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_3503),
.B(n_3524),
.Y(n_4922)
);

INVx2_ASAP7_75t_SL g4923 ( 
.A(n_3106),
.Y(n_4923)
);

A2O1A1Ixp33_ASAP7_75t_L g4924 ( 
.A1(n_3976),
.A2(n_4047),
.B(n_3606),
.C(n_3321),
.Y(n_4924)
);

INVx3_ASAP7_75t_L g4925 ( 
.A(n_3703),
.Y(n_4925)
);

AND2x2_ASAP7_75t_L g4926 ( 
.A(n_4033),
.B(n_4043),
.Y(n_4926)
);

CKINVDCx5p33_ASAP7_75t_R g4927 ( 
.A(n_3008),
.Y(n_4927)
);

A2O1A1Ixp33_ASAP7_75t_L g4928 ( 
.A1(n_4047),
.A2(n_3606),
.B(n_3318),
.C(n_3793),
.Y(n_4928)
);

A2O1A1Ixp33_ASAP7_75t_L g4929 ( 
.A1(n_3793),
.A2(n_3409),
.B(n_3411),
.C(n_3412),
.Y(n_4929)
);

AOI22xp5_ASAP7_75t_L g4930 ( 
.A1(n_3530),
.A2(n_3541),
.B1(n_3426),
.B2(n_3488),
.Y(n_4930)
);

O2A1O1Ixp33_ASAP7_75t_L g4931 ( 
.A1(n_3412),
.A2(n_3515),
.B(n_3426),
.C(n_3427),
.Y(n_4931)
);

BUFx2_ASAP7_75t_L g4932 ( 
.A(n_3305),
.Y(n_4932)
);

O2A1O1Ixp33_ASAP7_75t_L g4933 ( 
.A1(n_3424),
.A2(n_3500),
.B(n_3427),
.C(n_3525),
.Y(n_4933)
);

NOR2xp33_ASAP7_75t_L g4934 ( 
.A(n_3424),
.B(n_3457),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_3187),
.B(n_3192),
.Y(n_4935)
);

BUFx3_ASAP7_75t_L g4936 ( 
.A(n_3106),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_3392),
.A2(n_3111),
.B(n_3462),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_3392),
.A2(n_3476),
.B(n_3462),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_SL g4939 ( 
.A(n_3572),
.B(n_3582),
.Y(n_4939)
);

O2A1O1Ixp33_ASAP7_75t_L g4940 ( 
.A1(n_3457),
.A2(n_3512),
.B(n_3461),
.C(n_3525),
.Y(n_4940)
);

INVx3_ASAP7_75t_L g4941 ( 
.A(n_3703),
.Y(n_4941)
);

A2O1A1Ixp33_ASAP7_75t_L g4942 ( 
.A1(n_3461),
.A2(n_3512),
.B(n_3515),
.C(n_3516),
.Y(n_4942)
);

NOR2x1_ASAP7_75t_R g4943 ( 
.A(n_3499),
.B(n_3008),
.Y(n_4943)
);

AOI21xp5_ASAP7_75t_L g4944 ( 
.A1(n_3408),
.A2(n_3462),
.B(n_3476),
.Y(n_4944)
);

OR2x2_ASAP7_75t_L g4945 ( 
.A(n_2938),
.B(n_3733),
.Y(n_4945)
);

AOI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_3408),
.A2(n_3462),
.B(n_3476),
.Y(n_4946)
);

O2A1O1Ixp5_ASAP7_75t_L g4947 ( 
.A1(n_3511),
.A2(n_4065),
.B(n_3136),
.C(n_3169),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_3187),
.B(n_3192),
.Y(n_4948)
);

OAI22xp5_ASAP7_75t_L g4949 ( 
.A1(n_3465),
.A2(n_3516),
.B1(n_3478),
.B2(n_3482),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_3187),
.B(n_3192),
.Y(n_4950)
);

A2O1A1Ixp33_ASAP7_75t_L g4951 ( 
.A1(n_3465),
.A2(n_3522),
.B(n_3486),
.C(n_3482),
.Y(n_4951)
);

O2A1O1Ixp33_ASAP7_75t_L g4952 ( 
.A1(n_3478),
.A2(n_3522),
.B(n_3518),
.C(n_3486),
.Y(n_4952)
);

OAI22xp5_ASAP7_75t_SL g4953 ( 
.A1(n_2938),
.A2(n_3783),
.B1(n_3733),
.B2(n_4020),
.Y(n_4953)
);

OAI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4065),
.A2(n_3757),
.B(n_4020),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_SL g4955 ( 
.A(n_3572),
.B(n_3582),
.Y(n_4955)
);

INVxp67_ASAP7_75t_L g4956 ( 
.A(n_3541),
.Y(n_4956)
);

OAI22xp5_ASAP7_75t_L g4957 ( 
.A1(n_3008),
.A2(n_3968),
.B1(n_3243),
.B2(n_3899),
.Y(n_4957)
);

AOI21xp5_ASAP7_75t_L g4958 ( 
.A1(n_3408),
.A2(n_3476),
.B(n_3417),
.Y(n_4958)
);

NOR2xp33_ASAP7_75t_L g4959 ( 
.A(n_3130),
.B(n_3163),
.Y(n_4959)
);

OAI22xp5_ASAP7_75t_SL g4960 ( 
.A1(n_3757),
.A2(n_3921),
.B1(n_3783),
.B2(n_3703),
.Y(n_4960)
);

O2A1O1Ixp5_ASAP7_75t_L g4961 ( 
.A1(n_3136),
.A2(n_3997),
.B(n_3169),
.C(n_3712),
.Y(n_4961)
);

OAI22xp5_ASAP7_75t_L g4962 ( 
.A1(n_3243),
.A2(n_3968),
.B1(n_3899),
.B2(n_3921),
.Y(n_4962)
);

OR2x2_ASAP7_75t_L g4963 ( 
.A(n_3130),
.B(n_3163),
.Y(n_4963)
);

INVx1_ASAP7_75t_SL g4964 ( 
.A(n_3604),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_3243),
.Y(n_4965)
);

A2O1A1Ixp33_ASAP7_75t_SL g4966 ( 
.A1(n_3494),
.A2(n_3497),
.B(n_2998),
.C(n_4060),
.Y(n_4966)
);

AOI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_3408),
.A2(n_3462),
.B(n_3450),
.Y(n_4967)
);

BUFx6f_ASAP7_75t_L g4968 ( 
.A(n_3106),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_SL g4969 ( 
.A(n_3572),
.B(n_3582),
.Y(n_4969)
);

BUFx6f_ASAP7_75t_L g4970 ( 
.A(n_3106),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_SL g4971 ( 
.A(n_3582),
.B(n_3564),
.Y(n_4971)
);

O2A1O1Ixp5_ASAP7_75t_L g4972 ( 
.A1(n_3997),
.A2(n_3876),
.B(n_3712),
.C(n_3940),
.Y(n_4972)
);

AOI21xp5_ASAP7_75t_L g4973 ( 
.A1(n_3408),
.A2(n_3476),
.B(n_3417),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_SL g4974 ( 
.A(n_3582),
.B(n_3564),
.Y(n_4974)
);

BUFx6f_ASAP7_75t_L g4975 ( 
.A(n_3106),
.Y(n_4975)
);

BUFx6f_ASAP7_75t_L g4976 ( 
.A(n_3182),
.Y(n_4976)
);

OAI22xp5_ASAP7_75t_L g4977 ( 
.A1(n_3899),
.A2(n_3968),
.B1(n_3004),
.B2(n_4049),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_3604),
.Y(n_4978)
);

BUFx2_ASAP7_75t_L g4979 ( 
.A(n_3876),
.Y(n_4979)
);

NOR2xp33_ASAP7_75t_L g4980 ( 
.A(n_3604),
.B(n_3876),
.Y(n_4980)
);

NOR2xp33_ASAP7_75t_L g4981 ( 
.A(n_3940),
.B(n_4049),
.Y(n_4981)
);

HB1xp67_ASAP7_75t_L g4982 ( 
.A(n_3190),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_3193),
.B(n_3202),
.Y(n_4983)
);

A2O1A1Ixp33_ASAP7_75t_L g4984 ( 
.A1(n_3190),
.A2(n_3597),
.B(n_3593),
.C(n_3635),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_3193),
.B(n_3202),
.Y(n_4985)
);

INVx3_ASAP7_75t_L g4986 ( 
.A(n_3781),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_SL g4987 ( 
.A(n_3582),
.B(n_3564),
.Y(n_4987)
);

AOI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_3408),
.A2(n_3462),
.B(n_3417),
.Y(n_4988)
);

AOI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_3408),
.A2(n_3462),
.B(n_3417),
.Y(n_4989)
);

AOI22xp5_ASAP7_75t_L g4990 ( 
.A1(n_4049),
.A2(n_3635),
.B1(n_3004),
.B2(n_3997),
.Y(n_4990)
);

AOI22xp5_ASAP7_75t_L g4991 ( 
.A1(n_4049),
.A2(n_3004),
.B1(n_3997),
.B2(n_3574),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_3417),
.A2(n_3476),
.B(n_3450),
.Y(n_4992)
);

HB1xp67_ASAP7_75t_L g4993 ( 
.A(n_3182),
.Y(n_4993)
);

OR2x6_ASAP7_75t_L g4994 ( 
.A(n_3997),
.B(n_3182),
.Y(n_4994)
);

NOR2xp33_ASAP7_75t_R g4995 ( 
.A(n_3494),
.B(n_3497),
.Y(n_4995)
);

OAI22xp5_ASAP7_75t_L g4996 ( 
.A1(n_3182),
.A2(n_3214),
.B1(n_3185),
.B2(n_3781),
.Y(n_4996)
);

O2A1O1Ixp33_ASAP7_75t_L g4997 ( 
.A1(n_3560),
.A2(n_3581),
.B(n_3567),
.C(n_3574),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_3182),
.Y(n_4998)
);

AOI21xp5_ASAP7_75t_L g4999 ( 
.A1(n_3417),
.A2(n_3476),
.B(n_3450),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_3182),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_3209),
.B(n_3240),
.Y(n_5001)
);

NOR2x1_ASAP7_75t_L g5002 ( 
.A(n_3576),
.B(n_3560),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_3240),
.B(n_3259),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_3185),
.Y(n_5004)
);

HB1xp67_ASAP7_75t_L g5005 ( 
.A(n_3185),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_3185),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_3185),
.B(n_3214),
.Y(n_5007)
);

BUFx6f_ASAP7_75t_L g5008 ( 
.A(n_3185),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_SL g5009 ( 
.A(n_3582),
.B(n_3214),
.Y(n_5009)
);

BUFx2_ASAP7_75t_L g5010 ( 
.A(n_3214),
.Y(n_5010)
);

A2O1A1Ixp33_ASAP7_75t_L g5011 ( 
.A1(n_3593),
.A2(n_3597),
.B(n_3598),
.C(n_3219),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_3214),
.B(n_3642),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_3259),
.B(n_3359),
.Y(n_5013)
);

AOI22xp5_ASAP7_75t_L g5014 ( 
.A1(n_3567),
.A2(n_3581),
.B1(n_3214),
.B2(n_3576),
.Y(n_5014)
);

BUFx2_ASAP7_75t_L g5015 ( 
.A(n_3167),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_3219),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_3417),
.A2(n_3450),
.B(n_3363),
.Y(n_5017)
);

AOI21xp5_ASAP7_75t_L g5018 ( 
.A1(n_3450),
.A2(n_3363),
.B(n_3576),
.Y(n_5018)
);

NOR2xp33_ASAP7_75t_L g5019 ( 
.A(n_2998),
.B(n_3954),
.Y(n_5019)
);

NOR2xp33_ASAP7_75t_L g5020 ( 
.A(n_3642),
.B(n_3954),
.Y(n_5020)
);

AOI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_3450),
.A2(n_3315),
.B(n_3184),
.Y(n_5021)
);

NAND2xp33_ASAP7_75t_L g5022 ( 
.A(n_3450),
.B(n_3601),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_3286),
.B(n_3372),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_SL g5024 ( 
.A(n_3598),
.B(n_2947),
.Y(n_5024)
);

AOI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_3184),
.A2(n_3315),
.B(n_3341),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_3184),
.A2(n_3315),
.B(n_3341),
.Y(n_5026)
);

AOI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_3286),
.A2(n_3372),
.B1(n_3361),
.B2(n_3359),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_L g5028 ( 
.A(n_3642),
.B(n_3717),
.Y(n_5028)
);

OAI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_3544),
.A2(n_3167),
.B(n_3781),
.Y(n_5029)
);

OAI21x1_ASAP7_75t_L g5030 ( 
.A1(n_3781),
.A2(n_3683),
.B(n_3953),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_3184),
.A2(n_3315),
.B(n_3372),
.Y(n_5031)
);

A2O1A1Ixp33_ASAP7_75t_L g5032 ( 
.A1(n_3675),
.A2(n_3700),
.B(n_3826),
.C(n_3895),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_3308),
.B(n_3329),
.Y(n_5033)
);

A2O1A1Ixp33_ASAP7_75t_L g5034 ( 
.A1(n_3675),
.A2(n_3700),
.B(n_3826),
.C(n_3895),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_3683),
.B(n_3717),
.Y(n_5035)
);

OAI22xp5_ASAP7_75t_L g5036 ( 
.A1(n_3675),
.A2(n_3700),
.B1(n_3826),
.B2(n_3895),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_3308),
.B(n_3361),
.Y(n_5037)
);

INVx4_ASAP7_75t_L g5038 ( 
.A(n_2947),
.Y(n_5038)
);

O2A1O1Ixp33_ASAP7_75t_L g5039 ( 
.A1(n_3683),
.A2(n_3717),
.B(n_3851),
.C(n_3865),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_3329),
.A2(n_3361),
.B(n_3359),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_3329),
.B(n_3341),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_3006),
.B(n_3067),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_3006),
.B(n_3067),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_3544),
.Y(n_5044)
);

AOI22xp5_ASAP7_75t_L g5045 ( 
.A1(n_4062),
.A2(n_3717),
.B1(n_3954),
.B2(n_3953),
.Y(n_5045)
);

AOI22xp33_ASAP7_75t_L g5046 ( 
.A1(n_2947),
.A2(n_3823),
.B1(n_3860),
.B2(n_3991),
.Y(n_5046)
);

CKINVDCx16_ASAP7_75t_R g5047 ( 
.A(n_3499),
.Y(n_5047)
);

OAI22xp5_ASAP7_75t_L g5048 ( 
.A1(n_3601),
.A2(n_4060),
.B1(n_3954),
.B2(n_3953),
.Y(n_5048)
);

NAND3xp33_ASAP7_75t_L g5049 ( 
.A(n_2947),
.B(n_3823),
.C(n_3860),
.Y(n_5049)
);

NOR2xp33_ASAP7_75t_L g5050 ( 
.A(n_3683),
.B(n_4060),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_3311),
.Y(n_5051)
);

AOI221xp5_ASAP7_75t_L g5052 ( 
.A1(n_3851),
.A2(n_4060),
.B1(n_3953),
.B2(n_3865),
.C(n_3796),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_3006),
.B(n_3067),
.Y(n_5053)
);

O2A1O1Ixp33_ASAP7_75t_L g5054 ( 
.A1(n_3851),
.A2(n_3865),
.B(n_3006),
.C(n_3067),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_SL g5055 ( 
.A(n_2947),
.B(n_3823),
.Y(n_5055)
);

OAI22x1_ASAP7_75t_L g5056 ( 
.A1(n_3851),
.A2(n_3865),
.B1(n_3284),
.B2(n_3135),
.Y(n_5056)
);

BUFx3_ASAP7_75t_L g5057 ( 
.A(n_4062),
.Y(n_5057)
);

NOR2xp67_ASAP7_75t_L g5058 ( 
.A(n_3135),
.B(n_3284),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_3135),
.B(n_3284),
.Y(n_5059)
);

INVx4_ASAP7_75t_L g5060 ( 
.A(n_3796),
.Y(n_5060)
);

NOR2xp67_ASAP7_75t_SL g5061 ( 
.A(n_3796),
.B(n_3823),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_3311),
.Y(n_5062)
);

AOI221xp5_ASAP7_75t_L g5063 ( 
.A1(n_3796),
.A2(n_3823),
.B1(n_3991),
.B2(n_3982),
.C(n_3956),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_3311),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_3348),
.Y(n_5065)
);

OR2x6_ASAP7_75t_SL g5066 ( 
.A(n_4062),
.B(n_3429),
.Y(n_5066)
);

BUFx4_ASAP7_75t_SL g5067 ( 
.A(n_3429),
.Y(n_5067)
);

OAI22xp5_ASAP7_75t_L g5068 ( 
.A1(n_3601),
.A2(n_3823),
.B1(n_3991),
.B2(n_3982),
.Y(n_5068)
);

HB1xp67_ASAP7_75t_L g5069 ( 
.A(n_3348),
.Y(n_5069)
);

NOR2xp33_ASAP7_75t_L g5070 ( 
.A(n_3796),
.B(n_3823),
.Y(n_5070)
);

AOI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_3348),
.A2(n_3377),
.B(n_3379),
.Y(n_5071)
);

BUFx6f_ASAP7_75t_L g5072 ( 
.A(n_3844),
.Y(n_5072)
);

AOI21xp5_ASAP7_75t_L g5073 ( 
.A1(n_3348),
.A2(n_3377),
.B(n_3379),
.Y(n_5073)
);

A2O1A1Ixp33_ASAP7_75t_L g5074 ( 
.A1(n_3844),
.A2(n_3860),
.B(n_3991),
.C(n_3982),
.Y(n_5074)
);

BUFx3_ASAP7_75t_L g5075 ( 
.A(n_4062),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_3135),
.B(n_3284),
.Y(n_5076)
);

OAI22xp5_ASAP7_75t_L g5077 ( 
.A1(n_3601),
.A2(n_3872),
.B1(n_3991),
.B2(n_3982),
.Y(n_5077)
);

AOI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_3377),
.A2(n_3379),
.B(n_3872),
.Y(n_5078)
);

AOI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_3377),
.A2(n_3379),
.B(n_3872),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_SL g5080 ( 
.A(n_3844),
.B(n_3872),
.Y(n_5080)
);

HAxp5_ASAP7_75t_L g5081 ( 
.A(n_3429),
.B(n_4062),
.CON(n_5081),
.SN(n_5081)
);

NAND2xp5_ASAP7_75t_SL g5082 ( 
.A(n_3844),
.B(n_3872),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_3377),
.B(n_3379),
.Y(n_5083)
);

AOI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_3377),
.A2(n_3379),
.B(n_3872),
.Y(n_5084)
);

AOI21xp5_ASAP7_75t_L g5085 ( 
.A1(n_3844),
.A2(n_3893),
.B(n_3860),
.Y(n_5085)
);

O2A1O1Ixp33_ASAP7_75t_L g5086 ( 
.A1(n_3429),
.A2(n_4062),
.B(n_3844),
.C(n_3860),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_4062),
.B(n_3872),
.Y(n_5087)
);

AOI21xp5_ASAP7_75t_L g5088 ( 
.A1(n_3844),
.A2(n_3956),
.B(n_3860),
.Y(n_5088)
);

O2A1O1Ixp33_ASAP7_75t_L g5089 ( 
.A1(n_3429),
.A2(n_4062),
.B(n_3860),
.C(n_3893),
.Y(n_5089)
);

NAND2xp5_ASAP7_75t_L g5090 ( 
.A(n_4336),
.B(n_3893),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_5044),
.Y(n_5091)
);

HAxp5_ASAP7_75t_L g5092 ( 
.A(n_4148),
.B(n_3429),
.CON(n_5092),
.SN(n_5092)
);

CKINVDCx6p67_ASAP7_75t_R g5093 ( 
.A(n_4330),
.Y(n_5093)
);

BUFx6f_ASAP7_75t_L g5094 ( 
.A(n_4876),
.Y(n_5094)
);

NOR2xp33_ASAP7_75t_L g5095 ( 
.A(n_4162),
.B(n_3893),
.Y(n_5095)
);

INVx3_ASAP7_75t_L g5096 ( 
.A(n_4246),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5044),
.Y(n_5097)
);

BUFx3_ASAP7_75t_L g5098 ( 
.A(n_4799),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4650),
.Y(n_5099)
);

INVx4_ASAP7_75t_L g5100 ( 
.A(n_4876),
.Y(n_5100)
);

NOR2xp33_ASAP7_75t_L g5101 ( 
.A(n_4162),
.B(n_3893),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_4246),
.Y(n_5102)
);

A2O1A1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_4210),
.A2(n_3956),
.B(n_3982),
.C(n_3991),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4336),
.B(n_3956),
.Y(n_5104)
);

INVx3_ASAP7_75t_L g5105 ( 
.A(n_4246),
.Y(n_5105)
);

BUFx3_ASAP7_75t_L g5106 ( 
.A(n_4799),
.Y(n_5106)
);

BUFx2_ASAP7_75t_L g5107 ( 
.A(n_4913),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_5081),
.B(n_3956),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4650),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_5081),
.B(n_3956),
.Y(n_5110)
);

NAND3xp33_ASAP7_75t_L g5111 ( 
.A(n_4109),
.B(n_3956),
.C(n_3982),
.Y(n_5111)
);

CKINVDCx8_ASAP7_75t_R g5112 ( 
.A(n_4876),
.Y(n_5112)
);

AO32x2_ASAP7_75t_L g5113 ( 
.A1(n_4960),
.A2(n_3590),
.A3(n_3982),
.B1(n_3991),
.B2(n_4718),
.Y(n_5113)
);

AOI22xp33_ASAP7_75t_L g5114 ( 
.A1(n_4100),
.A2(n_3590),
.B1(n_4227),
.B2(n_4197),
.Y(n_5114)
);

BUFx12f_ASAP7_75t_L g5115 ( 
.A(n_4152),
.Y(n_5115)
);

OR2x6_ASAP7_75t_L g5116 ( 
.A(n_4770),
.B(n_3590),
.Y(n_5116)
);

AOI22xp33_ASAP7_75t_L g5117 ( 
.A1(n_4100),
.A2(n_3590),
.B1(n_4227),
.B2(n_4197),
.Y(n_5117)
);

INVx3_ASAP7_75t_L g5118 ( 
.A(n_4246),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_4671),
.Y(n_5119)
);

INVxp67_ASAP7_75t_SL g5120 ( 
.A(n_4745),
.Y(n_5120)
);

NAND2x1p5_ASAP7_75t_L g5121 ( 
.A(n_4876),
.B(n_3590),
.Y(n_5121)
);

BUFx8_ASAP7_75t_SL g5122 ( 
.A(n_4091),
.Y(n_5122)
);

BUFx16f_ASAP7_75t_R g5123 ( 
.A(n_4152),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_4347),
.B(n_3590),
.Y(n_5124)
);

HB1xp67_ASAP7_75t_L g5125 ( 
.A(n_4130),
.Y(n_5125)
);

BUFx2_ASAP7_75t_L g5126 ( 
.A(n_4913),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_4347),
.B(n_4370),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_5081),
.B(n_4070),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_4671),
.Y(n_5129)
);

HB1xp67_ASAP7_75t_L g5130 ( 
.A(n_4130),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4573),
.A2(n_4865),
.B(n_4848),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4370),
.B(n_4375),
.Y(n_5132)
);

BUFx2_ASAP7_75t_L g5133 ( 
.A(n_4913),
.Y(n_5133)
);

BUFx8_ASAP7_75t_SL g5134 ( 
.A(n_4314),
.Y(n_5134)
);

NOR2xp33_ASAP7_75t_R g5135 ( 
.A(n_4333),
.B(n_4497),
.Y(n_5135)
);

BUFx12f_ASAP7_75t_L g5136 ( 
.A(n_4152),
.Y(n_5136)
);

O2A1O1Ixp33_ASAP7_75t_L g5137 ( 
.A1(n_4095),
.A2(n_4198),
.B(n_4146),
.C(n_4184),
.Y(n_5137)
);

HB1xp67_ASAP7_75t_L g5138 ( 
.A(n_4072),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4746),
.Y(n_5139)
);

OAI22xp33_ASAP7_75t_L g5140 ( 
.A1(n_4199),
.A2(n_4141),
.B1(n_4303),
.B2(n_4077),
.Y(n_5140)
);

INVx5_ASAP7_75t_L g5141 ( 
.A(n_4876),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4375),
.B(n_4379),
.Y(n_5142)
);

BUFx2_ASAP7_75t_L g5143 ( 
.A(n_4913),
.Y(n_5143)
);

BUFx6f_ASAP7_75t_L g5144 ( 
.A(n_4876),
.Y(n_5144)
);

AOI22xp33_ASAP7_75t_L g5145 ( 
.A1(n_4134),
.A2(n_4110),
.B1(n_4109),
.B2(n_4209),
.Y(n_5145)
);

BUFx3_ASAP7_75t_L g5146 ( 
.A(n_4799),
.Y(n_5146)
);

NOR2xp33_ASAP7_75t_L g5147 ( 
.A(n_4141),
.B(n_4199),
.Y(n_5147)
);

BUFx4f_ASAP7_75t_L g5148 ( 
.A(n_4155),
.Y(n_5148)
);

BUFx12f_ASAP7_75t_L g5149 ( 
.A(n_4152),
.Y(n_5149)
);

NAND2x1p5_ASAP7_75t_L g5150 ( 
.A(n_4876),
.B(n_4114),
.Y(n_5150)
);

BUFx6f_ASAP7_75t_L g5151 ( 
.A(n_4550),
.Y(n_5151)
);

BUFx6f_ASAP7_75t_L g5152 ( 
.A(n_4550),
.Y(n_5152)
);

OAI22x1_ASAP7_75t_L g5153 ( 
.A1(n_4379),
.A2(n_4384),
.B1(n_4071),
.B2(n_4450),
.Y(n_5153)
);

INVxp67_ASAP7_75t_SL g5154 ( 
.A(n_4828),
.Y(n_5154)
);

BUFx3_ASAP7_75t_L g5155 ( 
.A(n_5066),
.Y(n_5155)
);

AND2x4_ASAP7_75t_L g5156 ( 
.A(n_4321),
.B(n_4344),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4364),
.B(n_4284),
.Y(n_5157)
);

BUFx2_ASAP7_75t_L g5158 ( 
.A(n_4913),
.Y(n_5158)
);

HB1xp67_ASAP7_75t_L g5159 ( 
.A(n_4072),
.Y(n_5159)
);

OR2x6_ASAP7_75t_L g5160 ( 
.A(n_4770),
.B(n_4845),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_SL g5161 ( 
.A(n_4219),
.B(n_4184),
.Y(n_5161)
);

HB1xp67_ASAP7_75t_L g5162 ( 
.A(n_4105),
.Y(n_5162)
);

AND2x4_ASAP7_75t_L g5163 ( 
.A(n_4321),
.B(n_4344),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_4364),
.B(n_4284),
.Y(n_5164)
);

INVx4_ASAP7_75t_L g5165 ( 
.A(n_4550),
.Y(n_5165)
);

AO32x1_ASAP7_75t_L g5166 ( 
.A1(n_4580),
.A2(n_4372),
.A3(n_4260),
.B1(n_4586),
.B2(n_4392),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_4110),
.A2(n_4209),
.B1(n_4101),
.B2(n_4260),
.Y(n_5167)
);

CKINVDCx5p33_ASAP7_75t_R g5168 ( 
.A(n_4252),
.Y(n_5168)
);

INVx3_ASAP7_75t_L g5169 ( 
.A(n_4246),
.Y(n_5169)
);

AND2x6_ASAP7_75t_L g5170 ( 
.A(n_4079),
.B(n_4096),
.Y(n_5170)
);

AOI222xp33_ASAP7_75t_L g5171 ( 
.A1(n_4188),
.A2(n_4077),
.B1(n_4069),
.B2(n_4087),
.C1(n_4081),
.C2(n_4220),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4749),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_4384),
.B(n_4283),
.Y(n_5173)
);

AOI21xp5_ASAP7_75t_L g5174 ( 
.A1(n_4573),
.A2(n_4848),
.B(n_4847),
.Y(n_5174)
);

AOI22xp5_ASAP7_75t_L g5175 ( 
.A1(n_4087),
.A2(n_4069),
.B1(n_4188),
.B2(n_4081),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4283),
.B(n_4158),
.Y(n_5176)
);

BUFx4f_ASAP7_75t_L g5177 ( 
.A(n_4155),
.Y(n_5177)
);

AOI21xp33_ASAP7_75t_SL g5178 ( 
.A1(n_4210),
.A2(n_4219),
.B(n_4303),
.Y(n_5178)
);

AND2x4_ASAP7_75t_L g5179 ( 
.A(n_4321),
.B(n_4344),
.Y(n_5179)
);

AOI21xp33_ASAP7_75t_L g5180 ( 
.A1(n_4261),
.A2(n_4281),
.B(n_4230),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4158),
.B(n_4167),
.Y(n_5181)
);

AOI22xp5_ASAP7_75t_L g5182 ( 
.A1(n_4147),
.A2(n_4362),
.B1(n_4256),
.B2(n_4356),
.Y(n_5182)
);

INVx3_ASAP7_75t_L g5183 ( 
.A(n_4267),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_SL g5184 ( 
.A(n_4261),
.B(n_4193),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4715),
.Y(n_5185)
);

AOI221x1_ASAP7_75t_L g5186 ( 
.A1(n_4117),
.A2(n_4175),
.B1(n_4183),
.B2(n_4256),
.C(n_4235),
.Y(n_5186)
);

BUFx2_ASAP7_75t_L g5187 ( 
.A(n_5066),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4715),
.Y(n_5188)
);

BUFx2_ASAP7_75t_L g5189 ( 
.A(n_5066),
.Y(n_5189)
);

BUFx8_ASAP7_75t_SL g5190 ( 
.A(n_4534),
.Y(n_5190)
);

AND2x4_ASAP7_75t_L g5191 ( 
.A(n_4321),
.B(n_4344),
.Y(n_5191)
);

AND2x4_ASAP7_75t_L g5192 ( 
.A(n_4321),
.B(n_4344),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_4075),
.B(n_4125),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4715),
.Y(n_5194)
);

BUFx2_ASAP7_75t_L g5195 ( 
.A(n_4727),
.Y(n_5195)
);

AND2x4_ASAP7_75t_L g5196 ( 
.A(n_4267),
.B(n_4770),
.Y(n_5196)
);

INVx2_ASAP7_75t_L g5197 ( 
.A(n_4697),
.Y(n_5197)
);

AND2x2_ASAP7_75t_L g5198 ( 
.A(n_4075),
.B(n_4125),
.Y(n_5198)
);

CKINVDCx5p33_ASAP7_75t_R g5199 ( 
.A(n_4377),
.Y(n_5199)
);

HB1xp67_ASAP7_75t_L g5200 ( 
.A(n_4105),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_SL g5201 ( 
.A(n_4193),
.B(n_4217),
.Y(n_5201)
);

NOR2xp33_ASAP7_75t_L g5202 ( 
.A(n_4133),
.B(n_4352),
.Y(n_5202)
);

CKINVDCx5p33_ASAP7_75t_R g5203 ( 
.A(n_4180),
.Y(n_5203)
);

AOI21xp5_ASAP7_75t_SL g5204 ( 
.A1(n_4266),
.A2(n_4421),
.B(n_4327),
.Y(n_5204)
);

OR2x6_ASAP7_75t_L g5205 ( 
.A(n_4770),
.B(n_4845),
.Y(n_5205)
);

BUFx6f_ASAP7_75t_L g5206 ( 
.A(n_4550),
.Y(n_5206)
);

BUFx3_ASAP7_75t_L g5207 ( 
.A(n_4507),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_4094),
.B(n_4104),
.Y(n_5208)
);

NOR2xp33_ASAP7_75t_L g5209 ( 
.A(n_4356),
.B(n_4243),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_4847),
.A2(n_4865),
.B(n_4853),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_4094),
.B(n_4104),
.Y(n_5211)
);

NOR2xp33_ASAP7_75t_L g5212 ( 
.A(n_4329),
.B(n_4258),
.Y(n_5212)
);

OR2x6_ASAP7_75t_L g5213 ( 
.A(n_4770),
.B(n_4845),
.Y(n_5213)
);

INVx1_ASAP7_75t_SL g5214 ( 
.A(n_4731),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_4715),
.Y(n_5215)
);

INVx4_ASAP7_75t_L g5216 ( 
.A(n_4124),
.Y(n_5216)
);

BUFx12f_ASAP7_75t_L g5217 ( 
.A(n_4152),
.Y(n_5217)
);

NAND2xp5_ASAP7_75t_L g5218 ( 
.A(n_4167),
.B(n_4412),
.Y(n_5218)
);

INVx3_ASAP7_75t_L g5219 ( 
.A(n_4267),
.Y(n_5219)
);

INVx2_ASAP7_75t_L g5220 ( 
.A(n_4732),
.Y(n_5220)
);

INVx2_ASAP7_75t_SL g5221 ( 
.A(n_4770),
.Y(n_5221)
);

A2O1A1Ixp33_ASAP7_75t_L g5222 ( 
.A1(n_4266),
.A2(n_4217),
.B(n_4242),
.C(n_4230),
.Y(n_5222)
);

A2O1A1Ixp33_ASAP7_75t_L g5223 ( 
.A1(n_4242),
.A2(n_4253),
.B(n_4362),
.C(n_4207),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_4715),
.Y(n_5224)
);

OAI31xp33_ASAP7_75t_SL g5225 ( 
.A1(n_4327),
.A2(n_4175),
.A3(n_4207),
.B(n_4235),
.Y(n_5225)
);

BUFx3_ASAP7_75t_L g5226 ( 
.A(n_4507),
.Y(n_5226)
);

BUFx12f_ASAP7_75t_L g5227 ( 
.A(n_4288),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_4732),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4715),
.Y(n_5229)
);

AOI22xp5_ASAP7_75t_L g5230 ( 
.A1(n_4329),
.A2(n_4201),
.B1(n_4117),
.B2(n_4071),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4715),
.Y(n_5231)
);

NOR2xp33_ASAP7_75t_L g5232 ( 
.A(n_4409),
.B(n_4145),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_4128),
.B(n_4273),
.Y(n_5233)
);

AOI221xp5_ASAP7_75t_L g5234 ( 
.A1(n_4241),
.A2(n_4253),
.B1(n_4183),
.B2(n_4281),
.C(n_4165),
.Y(n_5234)
);

INVx3_ASAP7_75t_L g5235 ( 
.A(n_4267),
.Y(n_5235)
);

AOI22xp5_ASAP7_75t_L g5236 ( 
.A1(n_4068),
.A2(n_4078),
.B1(n_4274),
.B2(n_4247),
.Y(n_5236)
);

O2A1O1Ixp33_ASAP7_75t_L g5237 ( 
.A1(n_4236),
.A2(n_4149),
.B(n_4232),
.C(n_4416),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_4302),
.B(n_4306),
.Y(n_5238)
);

INVxp67_ASAP7_75t_L g5239 ( 
.A(n_4390),
.Y(n_5239)
);

INVx1_ASAP7_75t_SL g5240 ( 
.A(n_4738),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_4125),
.B(n_4176),
.Y(n_5241)
);

OR2x6_ASAP7_75t_L g5242 ( 
.A(n_4845),
.B(n_4607),
.Y(n_5242)
);

BUFx3_ASAP7_75t_L g5243 ( 
.A(n_4622),
.Y(n_5243)
);

AOI22xp5_ASAP7_75t_L g5244 ( 
.A1(n_4274),
.A2(n_4247),
.B1(n_4289),
.B2(n_4367),
.Y(n_5244)
);

NOR2x1_ASAP7_75t_SL g5245 ( 
.A(n_4845),
.B(n_4215),
.Y(n_5245)
);

BUFx12f_ASAP7_75t_L g5246 ( 
.A(n_4288),
.Y(n_5246)
);

BUFx12f_ASAP7_75t_L g5247 ( 
.A(n_4288),
.Y(n_5247)
);

BUFx2_ASAP7_75t_L g5248 ( 
.A(n_4727),
.Y(n_5248)
);

OR2x6_ASAP7_75t_L g5249 ( 
.A(n_4845),
.B(n_4607),
.Y(n_5249)
);

A2O1A1Ixp33_ASAP7_75t_L g5250 ( 
.A1(n_4421),
.A2(n_4165),
.B(n_4156),
.C(n_4241),
.Y(n_5250)
);

AOI21x1_ASAP7_75t_L g5251 ( 
.A1(n_4114),
.A2(n_4194),
.B(n_4138),
.Y(n_5251)
);

OAI33xp33_ASAP7_75t_L g5252 ( 
.A1(n_4289),
.A2(n_4371),
.A3(n_4328),
.B1(n_4323),
.B2(n_4465),
.B3(n_4076),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4861),
.B(n_4884),
.Y(n_5253)
);

INVxp67_ASAP7_75t_SL g5254 ( 
.A(n_4853),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_4176),
.B(n_4211),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_4176),
.B(n_4211),
.Y(n_5256)
);

OAI22xp5_ASAP7_75t_L g5257 ( 
.A1(n_4124),
.A2(n_4218),
.B1(n_4297),
.B2(n_4316),
.Y(n_5257)
);

AND2x4_ASAP7_75t_L g5258 ( 
.A(n_4267),
.B(n_4369),
.Y(n_5258)
);

NAND2x1p5_ASAP7_75t_L g5259 ( 
.A(n_4138),
.B(n_4194),
.Y(n_5259)
);

AOI22xp5_ASAP7_75t_L g5260 ( 
.A1(n_4367),
.A2(n_4297),
.B1(n_4269),
.B2(n_4245),
.Y(n_5260)
);

CKINVDCx20_ASAP7_75t_R g5261 ( 
.A(n_4332),
.Y(n_5261)
);

INVx6_ASAP7_75t_L g5262 ( 
.A(n_4122),
.Y(n_5262)
);

AOI22xp33_ASAP7_75t_L g5263 ( 
.A1(n_4301),
.A2(n_4121),
.B1(n_4170),
.B2(n_4157),
.Y(n_5263)
);

INVxp67_ASAP7_75t_L g5264 ( 
.A(n_4390),
.Y(n_5264)
);

AND2x2_ASAP7_75t_L g5265 ( 
.A(n_4211),
.B(n_4265),
.Y(n_5265)
);

BUFx3_ASAP7_75t_L g5266 ( 
.A(n_4622),
.Y(n_5266)
);

NOR2xp33_ASAP7_75t_L g5267 ( 
.A(n_4427),
.B(n_4076),
.Y(n_5267)
);

AND2x4_ASAP7_75t_L g5268 ( 
.A(n_4369),
.B(n_4391),
.Y(n_5268)
);

CKINVDCx5p33_ASAP7_75t_R g5269 ( 
.A(n_4190),
.Y(n_5269)
);

BUFx4f_ASAP7_75t_SL g5270 ( 
.A(n_4628),
.Y(n_5270)
);

AOI22xp5_ASAP7_75t_L g5271 ( 
.A1(n_4269),
.A2(n_4316),
.B1(n_4354),
.B2(n_4106),
.Y(n_5271)
);

INVx2_ASAP7_75t_SL g5272 ( 
.A(n_4994),
.Y(n_5272)
);

CKINVDCx5p33_ASAP7_75t_R g5273 ( 
.A(n_4674),
.Y(n_5273)
);

O2A1O1Ixp5_ASAP7_75t_L g5274 ( 
.A1(n_4322),
.A2(n_4189),
.B(n_4140),
.C(n_4137),
.Y(n_5274)
);

AOI22xp5_ASAP7_75t_L g5275 ( 
.A1(n_4354),
.A2(n_4106),
.B1(n_4066),
.B2(n_4086),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_4127),
.Y(n_5276)
);

AOI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_4868),
.A2(n_4552),
.B(n_4742),
.Y(n_5277)
);

A2O1A1Ixp33_ASAP7_75t_L g5278 ( 
.A1(n_4156),
.A2(n_4218),
.B(n_4124),
.C(n_4380),
.Y(n_5278)
);

NAND2x2_ASAP7_75t_L g5279 ( 
.A(n_4226),
.B(n_4361),
.Y(n_5279)
);

NOR2xp67_ASAP7_75t_L g5280 ( 
.A(n_4744),
.B(n_4604),
.Y(n_5280)
);

NOR2xp67_ASAP7_75t_L g5281 ( 
.A(n_4744),
.B(n_4604),
.Y(n_5281)
);

BUFx2_ASAP7_75t_L g5282 ( 
.A(n_4405),
.Y(n_5282)
);

OR2x6_ASAP7_75t_L g5283 ( 
.A(n_4797),
.B(n_4552),
.Y(n_5283)
);

AND2x2_ASAP7_75t_L g5284 ( 
.A(n_4265),
.B(n_4309),
.Y(n_5284)
);

HB1xp67_ASAP7_75t_L g5285 ( 
.A(n_4089),
.Y(n_5285)
);

BUFx3_ASAP7_75t_L g5286 ( 
.A(n_4622),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_4343),
.B(n_4380),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4868),
.A2(n_4798),
.B(n_4777),
.Y(n_5288)
);

INVx4_ASAP7_75t_L g5289 ( 
.A(n_4124),
.Y(n_5289)
);

INVx1_ASAP7_75t_SL g5290 ( 
.A(n_4738),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_4383),
.B(n_4387),
.Y(n_5291)
);

INVx2_ASAP7_75t_SL g5292 ( 
.A(n_4994),
.Y(n_5292)
);

BUFx2_ASAP7_75t_L g5293 ( 
.A(n_4405),
.Y(n_5293)
);

CKINVDCx20_ASAP7_75t_R g5294 ( 
.A(n_4203),
.Y(n_5294)
);

BUFx12f_ASAP7_75t_L g5295 ( 
.A(n_4288),
.Y(n_5295)
);

INVx5_ASAP7_75t_L g5296 ( 
.A(n_4080),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4383),
.B(n_4387),
.Y(n_5297)
);

NAND2xp5_ASAP7_75t_L g5298 ( 
.A(n_4399),
.B(n_4407),
.Y(n_5298)
);

AOI22xp33_ASAP7_75t_L g5299 ( 
.A1(n_4121),
.A2(n_4144),
.B1(n_4585),
.B2(n_4407),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4841),
.A2(n_4538),
.B(n_4529),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_4089),
.Y(n_5301)
);

INVx4_ASAP7_75t_L g5302 ( 
.A(n_4218),
.Y(n_5302)
);

OAI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_4189),
.A2(n_4363),
.B(n_4366),
.Y(n_5303)
);

INVx2_ASAP7_75t_SL g5304 ( 
.A(n_4994),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_4265),
.B(n_4309),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4529),
.A2(n_4539),
.B(n_4538),
.Y(n_5306)
);

CKINVDCx5p33_ASAP7_75t_R g5307 ( 
.A(n_4792),
.Y(n_5307)
);

CKINVDCx5p33_ASAP7_75t_R g5308 ( 
.A(n_4119),
.Y(n_5308)
);

AND2x4_ASAP7_75t_L g5309 ( 
.A(n_4417),
.B(n_4234),
.Y(n_5309)
);

INVx1_ASAP7_75t_SL g5310 ( 
.A(n_4807),
.Y(n_5310)
);

BUFx12f_ASAP7_75t_L g5311 ( 
.A(n_4288),
.Y(n_5311)
);

INVx4_ASAP7_75t_L g5312 ( 
.A(n_4218),
.Y(n_5312)
);

AND2x4_ASAP7_75t_L g5313 ( 
.A(n_4417),
.B(n_4234),
.Y(n_5313)
);

OAI22xp5_ASAP7_75t_L g5314 ( 
.A1(n_4324),
.A2(n_4373),
.B1(n_4410),
.B2(n_4399),
.Y(n_5314)
);

INVx4_ASAP7_75t_L g5315 ( 
.A(n_4080),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_4410),
.B(n_4411),
.Y(n_5316)
);

BUFx6f_ASAP7_75t_L g5317 ( 
.A(n_4215),
.Y(n_5317)
);

BUFx6f_ASAP7_75t_L g5318 ( 
.A(n_4215),
.Y(n_5318)
);

NOR2xp33_ASAP7_75t_L g5319 ( 
.A(n_4427),
.B(n_4195),
.Y(n_5319)
);

BUFx2_ASAP7_75t_L g5320 ( 
.A(n_4405),
.Y(n_5320)
);

BUFx8_ASAP7_75t_L g5321 ( 
.A(n_4079),
.Y(n_5321)
);

BUFx2_ASAP7_75t_L g5322 ( 
.A(n_4405),
.Y(n_5322)
);

INVx1_ASAP7_75t_SL g5323 ( 
.A(n_4807),
.Y(n_5323)
);

OR2x6_ASAP7_75t_L g5324 ( 
.A(n_4797),
.B(n_4539),
.Y(n_5324)
);

AOI22xp33_ASAP7_75t_L g5325 ( 
.A1(n_4411),
.A2(n_4373),
.B1(n_4268),
.B2(n_4625),
.Y(n_5325)
);

BUFx12f_ASAP7_75t_L g5326 ( 
.A(n_4350),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_4861),
.B(n_4137),
.Y(n_5327)
);

OR2x2_ASAP7_75t_L g5328 ( 
.A(n_4755),
.B(n_4771),
.Y(n_5328)
);

INVx1_ASAP7_75t_SL g5329 ( 
.A(n_5015),
.Y(n_5329)
);

CKINVDCx5p33_ASAP7_75t_R g5330 ( 
.A(n_4181),
.Y(n_5330)
);

BUFx12f_ASAP7_75t_L g5331 ( 
.A(n_4350),
.Y(n_5331)
);

OR2x2_ASAP7_75t_L g5332 ( 
.A(n_4755),
.B(n_4771),
.Y(n_5332)
);

AND2x4_ASAP7_75t_L g5333 ( 
.A(n_4417),
.B(n_4240),
.Y(n_5333)
);

O2A1O1Ixp33_ASAP7_75t_L g5334 ( 
.A1(n_4420),
.A2(n_4345),
.B(n_4378),
.C(n_4366),
.Y(n_5334)
);

AOI22xp33_ASAP7_75t_L g5335 ( 
.A1(n_4268),
.A2(n_4702),
.B1(n_4582),
.B2(n_4298),
.Y(n_5335)
);

OR2x6_ASAP7_75t_L g5336 ( 
.A(n_4088),
.B(n_4090),
.Y(n_5336)
);

CKINVDCx5p33_ASAP7_75t_R g5337 ( 
.A(n_4536),
.Y(n_5337)
);

CKINVDCx5p33_ASAP7_75t_R g5338 ( 
.A(n_4643),
.Y(n_5338)
);

OAI21x1_ASAP7_75t_L g5339 ( 
.A1(n_4088),
.A2(n_4098),
.B(n_4090),
.Y(n_5339)
);

BUFx2_ASAP7_75t_L g5340 ( 
.A(n_4405),
.Y(n_5340)
);

AO21x1_ASAP7_75t_L g5341 ( 
.A1(n_4415),
.A2(n_4623),
.B(n_4418),
.Y(n_5341)
);

AND2x4_ASAP7_75t_L g5342 ( 
.A(n_4417),
.B(n_4240),
.Y(n_5342)
);

AND2x4_ASAP7_75t_L g5343 ( 
.A(n_4278),
.B(n_4556),
.Y(n_5343)
);

AND2x4_ASAP7_75t_L g5344 ( 
.A(n_4278),
.B(n_4556),
.Y(n_5344)
);

NOR2xp33_ASAP7_75t_SL g5345 ( 
.A(n_4850),
.B(n_4248),
.Y(n_5345)
);

AOI22xp33_ASAP7_75t_L g5346 ( 
.A1(n_4268),
.A2(n_4702),
.B1(n_4298),
.B2(n_4186),
.Y(n_5346)
);

BUFx6f_ASAP7_75t_L g5347 ( 
.A(n_4215),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_4309),
.B(n_4313),
.Y(n_5348)
);

BUFx12f_ASAP7_75t_L g5349 ( 
.A(n_4350),
.Y(n_5349)
);

NOR2xp33_ASAP7_75t_L g5350 ( 
.A(n_4195),
.B(n_4561),
.Y(n_5350)
);

AOI22xp33_ASAP7_75t_L g5351 ( 
.A1(n_4268),
.A2(n_4186),
.B1(n_4451),
.B2(n_4115),
.Y(n_5351)
);

OR2x6_ASAP7_75t_L g5352 ( 
.A(n_4098),
.B(n_4102),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_4324),
.A2(n_4491),
.B1(n_4531),
.B2(n_4639),
.Y(n_5353)
);

INVx2_ASAP7_75t_SL g5354 ( 
.A(n_4994),
.Y(n_5354)
);

NOR2xp33_ASAP7_75t_L g5355 ( 
.A(n_4561),
.B(n_4131),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_4102),
.A2(n_4108),
.B(n_4103),
.Y(n_5356)
);

INVx4_ASAP7_75t_L g5357 ( 
.A(n_4080),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_SL g5358 ( 
.A(n_4850),
.B(n_4248),
.Y(n_5358)
);

BUFx6f_ASAP7_75t_L g5359 ( 
.A(n_4215),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_4313),
.B(n_4817),
.Y(n_5360)
);

INVx2_ASAP7_75t_SL g5361 ( 
.A(n_4994),
.Y(n_5361)
);

AOI22xp33_ASAP7_75t_L g5362 ( 
.A1(n_4451),
.A2(n_4115),
.B1(n_4208),
.B2(n_4282),
.Y(n_5362)
);

NOR2xp33_ASAP7_75t_L g5363 ( 
.A(n_4131),
.B(n_4132),
.Y(n_5363)
);

INVxp67_ASAP7_75t_SL g5364 ( 
.A(n_4997),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_L g5365 ( 
.A(n_4884),
.B(n_4934),
.Y(n_5365)
);

AND2x2_ASAP7_75t_L g5366 ( 
.A(n_4313),
.B(n_4817),
.Y(n_5366)
);

OAI22xp5_ASAP7_75t_L g5367 ( 
.A1(n_4491),
.A2(n_4531),
.B1(n_4682),
.B2(n_4555),
.Y(n_5367)
);

AOI22xp5_ASAP7_75t_L g5368 ( 
.A1(n_4066),
.A2(n_4086),
.B1(n_4208),
.B2(n_4434),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_4934),
.B(n_4634),
.Y(n_5369)
);

BUFx8_ASAP7_75t_L g5370 ( 
.A(n_4079),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_4817),
.B(n_4215),
.Y(n_5371)
);

BUFx6f_ASAP7_75t_L g5372 ( 
.A(n_4079),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_4634),
.B(n_4780),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_4780),
.B(n_4869),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_4546),
.Y(n_5375)
);

NOR2xp33_ASAP7_75t_L g5376 ( 
.A(n_4132),
.B(n_4465),
.Y(n_5376)
);

BUFx2_ASAP7_75t_L g5377 ( 
.A(n_4897),
.Y(n_5377)
);

AOI22xp33_ASAP7_75t_SL g5378 ( 
.A1(n_4611),
.A2(n_4568),
.B1(n_4655),
.B2(n_4593),
.Y(n_5378)
);

INVx2_ASAP7_75t_SL g5379 ( 
.A(n_4994),
.Y(n_5379)
);

BUFx2_ASAP7_75t_R g5380 ( 
.A(n_4248),
.Y(n_5380)
);

BUFx6f_ASAP7_75t_L g5381 ( 
.A(n_4079),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_L g5382 ( 
.A(n_4140),
.B(n_4244),
.Y(n_5382)
);

OAI22xp5_ASAP7_75t_L g5383 ( 
.A1(n_4682),
.A2(n_4541),
.B1(n_4566),
.B2(n_4555),
.Y(n_5383)
);

BUFx6f_ASAP7_75t_L g5384 ( 
.A(n_4079),
.Y(n_5384)
);

NOR2xp33_ASAP7_75t_L g5385 ( 
.A(n_4518),
.B(n_4425),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_4244),
.B(n_4103),
.Y(n_5386)
);

NAND2xp5_ASAP7_75t_L g5387 ( 
.A(n_4108),
.B(n_4113),
.Y(n_5387)
);

AOI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_4434),
.A2(n_4516),
.B1(n_4514),
.B2(n_4611),
.Y(n_5388)
);

OR2x6_ASAP7_75t_L g5389 ( 
.A(n_4113),
.B(n_4116),
.Y(n_5389)
);

NOR2xp33_ASAP7_75t_L g5390 ( 
.A(n_4425),
.B(n_4773),
.Y(n_5390)
);

BUFx2_ASAP7_75t_L g5391 ( 
.A(n_4897),
.Y(n_5391)
);

AOI21x1_ASAP7_75t_L g5392 ( 
.A1(n_4251),
.A2(n_4877),
.B(n_4111),
.Y(n_5392)
);

NAND2xp5_ASAP7_75t_L g5393 ( 
.A(n_4116),
.B(n_4123),
.Y(n_5393)
);

OAI22x1_ASAP7_75t_L g5394 ( 
.A1(n_4450),
.A2(n_4659),
.B1(n_4667),
.B2(n_4067),
.Y(n_5394)
);

INVx3_ASAP7_75t_L g5395 ( 
.A(n_4645),
.Y(n_5395)
);

AOI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_4123),
.A2(n_4163),
.B(n_4129),
.Y(n_5396)
);

OAI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_4541),
.A2(n_4566),
.B1(n_4621),
.B2(n_4540),
.Y(n_5397)
);

CKINVDCx16_ASAP7_75t_R g5398 ( 
.A(n_4842),
.Y(n_5398)
);

INVx1_ASAP7_75t_SL g5399 ( 
.A(n_5015),
.Y(n_5399)
);

BUFx4f_ASAP7_75t_L g5400 ( 
.A(n_4155),
.Y(n_5400)
);

AOI22xp33_ASAP7_75t_L g5401 ( 
.A1(n_4282),
.A2(n_4773),
.B1(n_4355),
.B2(n_4413),
.Y(n_5401)
);

BUFx6f_ASAP7_75t_L g5402 ( 
.A(n_4079),
.Y(n_5402)
);

AOI22x1_ASAP7_75t_L g5403 ( 
.A1(n_4415),
.A2(n_4126),
.B1(n_4740),
.B2(n_4163),
.Y(n_5403)
);

BUFx6f_ASAP7_75t_L g5404 ( 
.A(n_4096),
.Y(n_5404)
);

NAND2xp5_ASAP7_75t_L g5405 ( 
.A(n_4129),
.B(n_4166),
.Y(n_5405)
);

BUFx6f_ASAP7_75t_L g5406 ( 
.A(n_4096),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_4166),
.B(n_4172),
.Y(n_5407)
);

INVx6_ASAP7_75t_L g5408 ( 
.A(n_4122),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_4172),
.B(n_4177),
.Y(n_5409)
);

OR2x6_ASAP7_75t_L g5410 ( 
.A(n_4177),
.B(n_4178),
.Y(n_5410)
);

BUFx6f_ASAP7_75t_L g5411 ( 
.A(n_4096),
.Y(n_5411)
);

AOI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_4178),
.A2(n_4205),
.B(n_4204),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_4204),
.B(n_4205),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_4216),
.B(n_4221),
.Y(n_5414)
);

BUFx4f_ASAP7_75t_L g5415 ( 
.A(n_4155),
.Y(n_5415)
);

NOR2xp33_ASAP7_75t_SL g5416 ( 
.A(n_4097),
.B(n_4206),
.Y(n_5416)
);

BUFx6f_ASAP7_75t_L g5417 ( 
.A(n_4096),
.Y(n_5417)
);

OAI22xp5_ASAP7_75t_L g5418 ( 
.A1(n_4621),
.A2(n_4540),
.B1(n_4182),
.B2(n_4381),
.Y(n_5418)
);

NOR2xp33_ASAP7_75t_L g5419 ( 
.A(n_4479),
.B(n_4477),
.Y(n_5419)
);

BUFx6f_ASAP7_75t_L g5420 ( 
.A(n_4096),
.Y(n_5420)
);

AOI222xp33_ASAP7_75t_L g5421 ( 
.A1(n_4396),
.A2(n_4524),
.B1(n_4577),
.B2(n_4355),
.C1(n_4583),
.C2(n_4372),
.Y(n_5421)
);

NOR2xp33_ASAP7_75t_SL g5422 ( 
.A(n_4097),
.B(n_4206),
.Y(n_5422)
);

INVx2_ASAP7_75t_SL g5423 ( 
.A(n_5067),
.Y(n_5423)
);

NAND2xp33_ASAP7_75t_L g5424 ( 
.A(n_4762),
.B(n_4772),
.Y(n_5424)
);

NOR2x1_ASAP7_75t_L g5425 ( 
.A(n_4067),
.B(n_4695),
.Y(n_5425)
);

NAND2xp5_ASAP7_75t_L g5426 ( 
.A(n_4216),
.B(n_4221),
.Y(n_5426)
);

OAI22xp33_ASAP7_75t_L g5427 ( 
.A1(n_4299),
.A2(n_4605),
.B1(n_4774),
.B2(n_4649),
.Y(n_5427)
);

AOI21xp33_ASAP7_75t_L g5428 ( 
.A1(n_4378),
.A2(n_4406),
.B(n_4394),
.Y(n_5428)
);

NOR2x1p5_ASAP7_75t_L g5429 ( 
.A(n_4629),
.B(n_4664),
.Y(n_5429)
);

OR2x2_ASAP7_75t_L g5430 ( 
.A(n_4755),
.B(n_4771),
.Y(n_5430)
);

INVx1_ASAP7_75t_SL g5431 ( 
.A(n_4982),
.Y(n_5431)
);

O2A1O1Ixp33_ASAP7_75t_SL g5432 ( 
.A1(n_4476),
.A2(n_4900),
.B(n_4730),
.C(n_4590),
.Y(n_5432)
);

OAI22x1_ASAP7_75t_L g5433 ( 
.A1(n_4659),
.A2(n_4667),
.B1(n_4990),
.B2(n_4840),
.Y(n_5433)
);

BUFx10_ASAP7_75t_L g5434 ( 
.A(n_4484),
.Y(n_5434)
);

INVx2_ASAP7_75t_SL g5435 ( 
.A(n_5067),
.Y(n_5435)
);

AOI22xp5_ASAP7_75t_L g5436 ( 
.A1(n_4605),
.A2(n_4396),
.B1(n_4598),
.B2(n_4593),
.Y(n_5436)
);

INVx3_ASAP7_75t_SL g5437 ( 
.A(n_4568),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_4869),
.B(n_4872),
.Y(n_5438)
);

A2O1A1Ixp33_ASAP7_75t_L g5439 ( 
.A1(n_4394),
.A2(n_4406),
.B(n_4444),
.C(n_5086),
.Y(n_5439)
);

OAI22xp5_ASAP7_75t_L g5440 ( 
.A1(n_4182),
.A2(n_4381),
.B1(n_4617),
.B2(n_4513),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_4872),
.B(n_4914),
.Y(n_5441)
);

O2A1O1Ixp33_ASAP7_75t_L g5442 ( 
.A1(n_4287),
.A2(n_4349),
.B(n_4473),
.C(n_4569),
.Y(n_5442)
);

INVx1_ASAP7_75t_SL g5443 ( 
.A(n_4982),
.Y(n_5443)
);

A2O1A1Ixp33_ASAP7_75t_L g5444 ( 
.A1(n_4444),
.A2(n_5089),
.B(n_5086),
.C(n_4602),
.Y(n_5444)
);

CKINVDCx5p33_ASAP7_75t_R g5445 ( 
.A(n_4546),
.Y(n_5445)
);

AOI21xp5_ASAP7_75t_L g5446 ( 
.A1(n_4223),
.A2(n_4237),
.B(n_4231),
.Y(n_5446)
);

AND3x1_ASAP7_75t_SL g5447 ( 
.A(n_4803),
.B(n_4537),
.C(n_4779),
.Y(n_5447)
);

AOI22xp33_ASAP7_75t_L g5448 ( 
.A1(n_4688),
.A2(n_4469),
.B1(n_4478),
.B2(n_4251),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_4223),
.B(n_4231),
.Y(n_5449)
);

AOI22xp33_ASAP7_75t_L g5450 ( 
.A1(n_4688),
.A2(n_4474),
.B1(n_4598),
.B2(n_4584),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_4096),
.Y(n_5451)
);

INVx1_ASAP7_75t_SL g5452 ( 
.A(n_4619),
.Y(n_5452)
);

NAND2x1_ASAP7_75t_L g5453 ( 
.A(n_4270),
.B(n_4428),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_4914),
.B(n_4920),
.Y(n_5454)
);

INVx2_ASAP7_75t_SL g5455 ( 
.A(n_4676),
.Y(n_5455)
);

NOR2xp33_ASAP7_75t_R g5456 ( 
.A(n_5047),
.B(n_4784),
.Y(n_5456)
);

BUFx6f_ASAP7_75t_L g5457 ( 
.A(n_4120),
.Y(n_5457)
);

BUFx6f_ASAP7_75t_L g5458 ( 
.A(n_4120),
.Y(n_5458)
);

BUFx6f_ASAP7_75t_L g5459 ( 
.A(n_4120),
.Y(n_5459)
);

NAND2xp5_ASAP7_75t_L g5460 ( 
.A(n_4237),
.B(n_4249),
.Y(n_5460)
);

AOI221xp5_ASAP7_75t_L g5461 ( 
.A1(n_4287),
.A2(n_4349),
.B1(n_4448),
.B2(n_4255),
.C(n_4259),
.Y(n_5461)
);

BUFx4f_ASAP7_75t_L g5462 ( 
.A(n_4250),
.Y(n_5462)
);

AOI222xp33_ASAP7_75t_L g5463 ( 
.A1(n_4524),
.A2(n_4644),
.B1(n_4632),
.B2(n_4385),
.C1(n_4493),
.C2(n_4485),
.Y(n_5463)
);

AOI21xp5_ASAP7_75t_L g5464 ( 
.A1(n_4249),
.A2(n_4255),
.B(n_4254),
.Y(n_5464)
);

OAI22xp5_ASAP7_75t_L g5465 ( 
.A1(n_4182),
.A2(n_4381),
.B1(n_4617),
.B2(n_4513),
.Y(n_5465)
);

INVxp67_ASAP7_75t_SL g5466 ( 
.A(n_4997),
.Y(n_5466)
);

OAI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_4699),
.A2(n_4655),
.B1(n_4930),
.B2(n_4794),
.Y(n_5467)
);

AOI21x1_ASAP7_75t_L g5468 ( 
.A1(n_4877),
.A2(n_4111),
.B(n_4424),
.Y(n_5468)
);

AOI22xp33_ASAP7_75t_L g5469 ( 
.A1(n_4474),
.A2(n_4259),
.B1(n_4262),
.B2(n_4254),
.Y(n_5469)
);

INVx1_ASAP7_75t_SL g5470 ( 
.A(n_4619),
.Y(n_5470)
);

BUFx4f_ASAP7_75t_L g5471 ( 
.A(n_4250),
.Y(n_5471)
);

BUFx12f_ASAP7_75t_L g5472 ( 
.A(n_4350),
.Y(n_5472)
);

CKINVDCx5p33_ASAP7_75t_R g5473 ( 
.A(n_4708),
.Y(n_5473)
);

NAND2xp5_ASAP7_75t_L g5474 ( 
.A(n_4262),
.B(n_4277),
.Y(n_5474)
);

BUFx6f_ASAP7_75t_L g5475 ( 
.A(n_4120),
.Y(n_5475)
);

O2A1O1Ixp33_ASAP7_75t_L g5476 ( 
.A1(n_4473),
.A2(n_4311),
.B(n_4285),
.C(n_4549),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_4277),
.B(n_4280),
.Y(n_5477)
);

AOI21xp5_ASAP7_75t_SL g5478 ( 
.A1(n_4943),
.A2(n_4477),
.B(n_4736),
.Y(n_5478)
);

BUFx6f_ASAP7_75t_L g5479 ( 
.A(n_4120),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_L g5480 ( 
.A1(n_4280),
.A2(n_4295),
.B1(n_4312),
.B2(n_4291),
.Y(n_5480)
);

AO21x2_ASAP7_75t_L g5481 ( 
.A1(n_4886),
.A2(n_4295),
.B(n_4291),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_4312),
.B(n_4317),
.Y(n_5482)
);

AOI22xp33_ASAP7_75t_L g5483 ( 
.A1(n_4317),
.A2(n_4339),
.B1(n_4348),
.B2(n_4335),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_4335),
.B(n_4339),
.Y(n_5484)
);

OAI22xp5_ASAP7_75t_L g5485 ( 
.A1(n_4699),
.A2(n_4655),
.B1(n_4930),
.B2(n_4794),
.Y(n_5485)
);

OAI22xp5_ASAP7_75t_L g5486 ( 
.A1(n_4655),
.A2(n_4942),
.B1(n_4951),
.B2(n_4579),
.Y(n_5486)
);

BUFx6f_ASAP7_75t_L g5487 ( 
.A(n_4120),
.Y(n_5487)
);

CKINVDCx5p33_ASAP7_75t_R g5488 ( 
.A(n_4446),
.Y(n_5488)
);

BUFx6f_ASAP7_75t_L g5489 ( 
.A(n_4120),
.Y(n_5489)
);

INVxp67_ASAP7_75t_SL g5490 ( 
.A(n_5040),
.Y(n_5490)
);

INVx1_ASAP7_75t_SL g5491 ( 
.A(n_4789),
.Y(n_5491)
);

BUFx6f_ASAP7_75t_L g5492 ( 
.A(n_4150),
.Y(n_5492)
);

OAI22xp5_ASAP7_75t_L g5493 ( 
.A1(n_4579),
.A2(n_4311),
.B1(n_4285),
.B2(n_4843),
.Y(n_5493)
);

NOR2xp33_ASAP7_75t_L g5494 ( 
.A(n_4526),
.B(n_4685),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_4920),
.B(n_4949),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_4949),
.B(n_4603),
.Y(n_5496)
);

INVx1_ASAP7_75t_SL g5497 ( 
.A(n_4789),
.Y(n_5497)
);

CKINVDCx14_ASAP7_75t_R g5498 ( 
.A(n_4793),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_4348),
.B(n_4353),
.Y(n_5499)
);

NOR2x1_ASAP7_75t_R g5500 ( 
.A(n_4286),
.B(n_4568),
.Y(n_5500)
);

BUFx2_ASAP7_75t_SL g5501 ( 
.A(n_4122),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_4353),
.B(n_4725),
.Y(n_5502)
);

AOI22xp33_ASAP7_75t_L g5503 ( 
.A1(n_4568),
.A2(n_4496),
.B1(n_4644),
.B2(n_4632),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_4446),
.Y(n_5504)
);

CKINVDCx11_ASAP7_75t_R g5505 ( 
.A(n_4159),
.Y(n_5505)
);

INVxp67_ASAP7_75t_L g5506 ( 
.A(n_4858),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_4586),
.B(n_4685),
.Y(n_5507)
);

BUFx8_ASAP7_75t_SL g5508 ( 
.A(n_4286),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_4757),
.B(n_4891),
.Y(n_5509)
);

NAND2xp5_ASAP7_75t_L g5510 ( 
.A(n_4757),
.B(n_4891),
.Y(n_5510)
);

OAI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_4843),
.A2(n_4860),
.B1(n_4571),
.B2(n_4803),
.Y(n_5511)
);

A2O1A1Ixp33_ASAP7_75t_L g5512 ( 
.A1(n_5089),
.A2(n_4837),
.B(n_4448),
.C(n_4740),
.Y(n_5512)
);

INVx1_ASAP7_75t_SL g5513 ( 
.A(n_4789),
.Y(n_5513)
);

INVx2_ASAP7_75t_SL g5514 ( 
.A(n_4676),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_4931),
.B(n_4933),
.Y(n_5515)
);

BUFx6f_ASAP7_75t_L g5516 ( 
.A(n_4150),
.Y(n_5516)
);

OAI22xp5_ASAP7_75t_L g5517 ( 
.A1(n_4860),
.A2(n_4571),
.B1(n_4837),
.B2(n_4878),
.Y(n_5517)
);

NAND3xp33_ASAP7_75t_L g5518 ( 
.A(n_4196),
.B(n_4341),
.C(n_4304),
.Y(n_5518)
);

BUFx2_ASAP7_75t_L g5519 ( 
.A(n_4954),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_L g5520 ( 
.A1(n_4568),
.A2(n_4802),
.B1(n_4286),
.B2(n_4665),
.Y(n_5520)
);

NOR2xp33_ASAP7_75t_L g5521 ( 
.A(n_4629),
.B(n_4664),
.Y(n_5521)
);

NAND2xp5_ASAP7_75t_L g5522 ( 
.A(n_4931),
.B(n_4933),
.Y(n_5522)
);

NOR2xp67_ASAP7_75t_L g5523 ( 
.A(n_4895),
.B(n_4886),
.Y(n_5523)
);

INVx1_ASAP7_75t_SL g5524 ( 
.A(n_4136),
.Y(n_5524)
);

AOI222xp33_ASAP7_75t_L g5525 ( 
.A1(n_4385),
.A2(n_4468),
.B1(n_4456),
.B2(n_4808),
.C1(n_4673),
.C2(n_4665),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_4940),
.B(n_4952),
.Y(n_5526)
);

OAI22xp5_ASAP7_75t_L g5527 ( 
.A1(n_4571),
.A2(n_4878),
.B1(n_4919),
.B2(n_4887),
.Y(n_5527)
);

INVxp67_ASAP7_75t_L g5528 ( 
.A(n_4858),
.Y(n_5528)
);

AOI21xp5_ASAP7_75t_L g5529 ( 
.A1(n_4734),
.A2(n_4885),
.B(n_4836),
.Y(n_5529)
);

AOI22xp33_ASAP7_75t_L g5530 ( 
.A1(n_4350),
.A2(n_4673),
.B1(n_4665),
.B2(n_4505),
.Y(n_5530)
);

O2A1O1Ixp5_ASAP7_75t_L g5531 ( 
.A1(n_4304),
.A2(n_4341),
.B(n_4436),
.C(n_4422),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_4603),
.B(n_4296),
.Y(n_5532)
);

AOI22xp33_ASAP7_75t_L g5533 ( 
.A1(n_4665),
.A2(n_4673),
.B1(n_4503),
.B2(n_4299),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_4832),
.A2(n_4627),
.B1(n_4751),
.B2(n_4647),
.Y(n_5534)
);

CKINVDCx6p67_ASAP7_75t_R g5535 ( 
.A(n_4330),
.Y(n_5535)
);

BUFx12f_ASAP7_75t_L g5536 ( 
.A(n_4665),
.Y(n_5536)
);

AND2x2_ASAP7_75t_L g5537 ( 
.A(n_4840),
.B(n_4490),
.Y(n_5537)
);

AOI22xp33_ASAP7_75t_L g5538 ( 
.A1(n_4673),
.A2(n_4751),
.B1(n_4666),
.B2(n_4800),
.Y(n_5538)
);

INVx3_ASAP7_75t_SL g5539 ( 
.A(n_4168),
.Y(n_5539)
);

INVx2_ASAP7_75t_SL g5540 ( 
.A(n_4677),
.Y(n_5540)
);

BUFx2_ASAP7_75t_L g5541 ( 
.A(n_4954),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_4940),
.B(n_4952),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_4840),
.B(n_4490),
.Y(n_5543)
);

OAI22xp33_ASAP7_75t_L g5544 ( 
.A1(n_4649),
.A2(n_4517),
.B1(n_4308),
.B2(n_4408),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_4525),
.B(n_4594),
.Y(n_5545)
);

NOR2xp67_ASAP7_75t_L g5546 ( 
.A(n_4895),
.B(n_4122),
.Y(n_5546)
);

CKINVDCx16_ASAP7_75t_R g5547 ( 
.A(n_4881),
.Y(n_5547)
);

CKINVDCx20_ASAP7_75t_R g5548 ( 
.A(n_4673),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_4525),
.B(n_4594),
.Y(n_5549)
);

NOR2xp33_ASAP7_75t_L g5550 ( 
.A(n_4856),
.B(n_4857),
.Y(n_5550)
);

OAI22xp5_ASAP7_75t_L g5551 ( 
.A1(n_4887),
.A2(n_4919),
.B1(n_4679),
.B2(n_4559),
.Y(n_5551)
);

NOR2xp33_ASAP7_75t_L g5552 ( 
.A(n_4856),
.B(n_4857),
.Y(n_5552)
);

AND2x2_ASAP7_75t_L g5553 ( 
.A(n_4490),
.B(n_4502),
.Y(n_5553)
);

O2A1O1Ixp33_ASAP7_75t_L g5554 ( 
.A1(n_4549),
.A2(n_4560),
.B(n_4543),
.C(n_4825),
.Y(n_5554)
);

AOI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_4832),
.A2(n_4627),
.B1(n_4873),
.B2(n_4517),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_4502),
.B(n_4542),
.Y(n_5556)
);

INVx1_ASAP7_75t_SL g5557 ( 
.A(n_4401),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_4159),
.Y(n_5558)
);

INVxp67_ASAP7_75t_SL g5559 ( 
.A(n_5040),
.Y(n_5559)
);

O2A1O1Ixp33_ASAP7_75t_L g5560 ( 
.A1(n_4560),
.A2(n_4661),
.B(n_4535),
.C(n_4528),
.Y(n_5560)
);

AOI22xp33_ASAP7_75t_L g5561 ( 
.A1(n_4610),
.A2(n_4614),
.B1(n_4719),
.B2(n_4693),
.Y(n_5561)
);

CKINVDCx20_ASAP7_75t_R g5562 ( 
.A(n_4859),
.Y(n_5562)
);

A2O1A1Ixp33_ASAP7_75t_L g5563 ( 
.A1(n_4836),
.A2(n_4480),
.B(n_4606),
.C(n_4626),
.Y(n_5563)
);

OAI22xp5_ASAP7_75t_L g5564 ( 
.A1(n_4559),
.A2(n_4641),
.B1(n_4698),
.B2(n_4689),
.Y(n_5564)
);

AOI22xp33_ASAP7_75t_L g5565 ( 
.A1(n_4614),
.A2(n_4719),
.B1(n_4271),
.B2(n_4308),
.Y(n_5565)
);

OAI22xp5_ASAP7_75t_L g5566 ( 
.A1(n_4641),
.A2(n_4698),
.B1(n_4707),
.B2(n_4689),
.Y(n_5566)
);

OR2x6_ASAP7_75t_L g5567 ( 
.A(n_4527),
.B(n_4806),
.Y(n_5567)
);

BUFx4_ASAP7_75t_SL g5568 ( 
.A(n_4812),
.Y(n_5568)
);

NAND2xp5_ASAP7_75t_L g5569 ( 
.A(n_4779),
.B(n_4811),
.Y(n_5569)
);

NAND2xp5_ASAP7_75t_L g5570 ( 
.A(n_4811),
.B(n_4867),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_L g5571 ( 
.A(n_4867),
.B(n_4433),
.Y(n_5571)
);

CKINVDCx8_ASAP7_75t_R g5572 ( 
.A(n_5047),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_4502),
.B(n_4542),
.Y(n_5573)
);

A2O1A1Ixp33_ASAP7_75t_L g5574 ( 
.A1(n_4480),
.A2(n_4606),
.B(n_4626),
.C(n_4734),
.Y(n_5574)
);

AOI22xp5_ASAP7_75t_L g5575 ( 
.A1(n_4873),
.A2(n_4408),
.B1(n_4713),
.B2(n_4703),
.Y(n_5575)
);

A2O1A1Ixp33_ASAP7_75t_L g5576 ( 
.A1(n_4924),
.A2(n_4885),
.B(n_4748),
.C(n_4752),
.Y(n_5576)
);

AOI21xp5_ASAP7_75t_L g5577 ( 
.A1(n_4631),
.A2(n_4648),
.B(n_4638),
.Y(n_5577)
);

NAND2xp5_ASAP7_75t_L g5578 ( 
.A(n_4433),
.B(n_4441),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_SL g5579 ( 
.A(n_4741),
.B(n_4357),
.Y(n_5579)
);

AND2x2_ASAP7_75t_L g5580 ( 
.A(n_4542),
.B(n_4764),
.Y(n_5580)
);

AOI221xp5_ASAP7_75t_L g5581 ( 
.A1(n_4642),
.A2(n_4654),
.B1(n_4714),
.B2(n_4692),
.C(n_4680),
.Y(n_5581)
);

BUFx2_ASAP7_75t_SL g5582 ( 
.A(n_4122),
.Y(n_5582)
);

INVxp33_ASAP7_75t_L g5583 ( 
.A(n_4826),
.Y(n_5583)
);

BUFx12f_ASAP7_75t_L g5584 ( 
.A(n_4118),
.Y(n_5584)
);

AND2x4_ASAP7_75t_SL g5585 ( 
.A(n_4653),
.B(n_4164),
.Y(n_5585)
);

AOI22xp33_ASAP7_75t_L g5586 ( 
.A1(n_4271),
.A2(n_4722),
.B1(n_4718),
.B2(n_4728),
.Y(n_5586)
);

AND2x2_ASAP7_75t_L g5587 ( 
.A(n_4764),
.B(n_4782),
.Y(n_5587)
);

NOR2xp33_ASAP7_75t_L g5588 ( 
.A(n_4851),
.B(n_4871),
.Y(n_5588)
);

A2O1A1Ixp33_ASAP7_75t_L g5589 ( 
.A1(n_4748),
.A2(n_4752),
.B(n_4564),
.C(n_4741),
.Y(n_5589)
);

OR2x6_ASAP7_75t_L g5590 ( 
.A(n_4527),
.B(n_4806),
.Y(n_5590)
);

AOI22xp33_ASAP7_75t_SL g5591 ( 
.A1(n_4855),
.A2(n_4960),
.B1(n_4082),
.B2(n_4153),
.Y(n_5591)
);

BUFx4_ASAP7_75t_SL g5592 ( 
.A(n_4818),
.Y(n_5592)
);

AND2x6_ASAP7_75t_L g5593 ( 
.A(n_4233),
.B(n_4263),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_4686),
.Y(n_5594)
);

INVx4_ASAP7_75t_L g5595 ( 
.A(n_4233),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_4686),
.Y(n_5596)
);

AOI22xp5_ASAP7_75t_L g5597 ( 
.A1(n_4703),
.A2(n_4713),
.B1(n_4747),
.B2(n_4337),
.Y(n_5597)
);

AOI21xp5_ASAP7_75t_L g5598 ( 
.A1(n_4631),
.A2(n_4648),
.B(n_4638),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_4597),
.Y(n_5599)
);

AND2x4_ASAP7_75t_L g5600 ( 
.A(n_4894),
.B(n_4426),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_4684),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_4684),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_L g5603 ( 
.A(n_4441),
.B(n_4463),
.Y(n_5603)
);

INVx5_ASAP7_75t_L g5604 ( 
.A(n_4657),
.Y(n_5604)
);

AOI22xp33_ASAP7_75t_L g5605 ( 
.A1(n_4722),
.A2(n_4710),
.B1(n_4721),
.B2(n_4707),
.Y(n_5605)
);

O2A1O1Ixp33_ASAP7_75t_L g5606 ( 
.A1(n_4528),
.A2(n_4578),
.B(n_4574),
.C(n_4656),
.Y(n_5606)
);

AND3x1_ASAP7_75t_SL g5607 ( 
.A(n_4537),
.B(n_4118),
.C(n_4630),
.Y(n_5607)
);

INVx4_ASAP7_75t_L g5608 ( 
.A(n_4233),
.Y(n_5608)
);

AND2x6_ASAP7_75t_L g5609 ( 
.A(n_4233),
.B(n_4263),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_4463),
.B(n_4475),
.Y(n_5610)
);

INVx6_ASAP7_75t_L g5611 ( 
.A(n_4122),
.Y(n_5611)
);

BUFx8_ASAP7_75t_SL g5612 ( 
.A(n_4854),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_SL g5613 ( 
.A(n_4695),
.B(n_4595),
.Y(n_5613)
);

NOR2xp33_ASAP7_75t_L g5614 ( 
.A(n_4747),
.B(n_4608),
.Y(n_5614)
);

HB1xp67_ASAP7_75t_L g5615 ( 
.A(n_4945),
.Y(n_5615)
);

INVx5_ASAP7_75t_L g5616 ( 
.A(n_4657),
.Y(n_5616)
);

INVx2_ASAP7_75t_L g5617 ( 
.A(n_4597),
.Y(n_5617)
);

NOR2xp67_ASAP7_75t_L g5618 ( 
.A(n_4122),
.B(n_4151),
.Y(n_5618)
);

AND2x2_ASAP7_75t_L g5619 ( 
.A(n_4764),
.B(n_4782),
.Y(n_5619)
);

BUFx10_ASAP7_75t_L g5620 ( 
.A(n_4484),
.Y(n_5620)
);

CKINVDCx6p67_ASAP7_75t_R g5621 ( 
.A(n_4330),
.Y(n_5621)
);

OR2x2_ASAP7_75t_L g5622 ( 
.A(n_4911),
.B(n_4945),
.Y(n_5622)
);

A2O1A1Ixp33_ASAP7_75t_L g5623 ( 
.A1(n_4564),
.A2(n_4595),
.B(n_4511),
.C(n_4816),
.Y(n_5623)
);

OAI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_4710),
.A2(n_4721),
.B1(n_4481),
.B2(n_4515),
.Y(n_5624)
);

CKINVDCx5p33_ASAP7_75t_R g5625 ( 
.A(n_4159),
.Y(n_5625)
);

AOI22xp5_ASAP7_75t_L g5626 ( 
.A1(n_4337),
.A2(n_4515),
.B1(n_4475),
.B2(n_4481),
.Y(n_5626)
);

AOI22xp33_ASAP7_75t_L g5627 ( 
.A1(n_4530),
.A2(n_4112),
.B1(n_4464),
.B2(n_4107),
.Y(n_5627)
);

AOI21xp5_ASAP7_75t_L g5628 ( 
.A1(n_4658),
.A2(n_4662),
.B(n_4660),
.Y(n_5628)
);

OAI22xp33_ASAP7_75t_SL g5629 ( 
.A1(n_4651),
.A2(n_4392),
.B1(n_4795),
.B2(n_4082),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_4824),
.B(n_4635),
.Y(n_5630)
);

NAND2xp5_ASAP7_75t_L g5631 ( 
.A(n_4824),
.B(n_4635),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_4615),
.Y(n_5632)
);

AOI22xp33_ASAP7_75t_L g5633 ( 
.A1(n_4107),
.A2(n_4464),
.B1(n_4112),
.B2(n_4168),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_5029),
.Y(n_5634)
);

AND2x4_ASAP7_75t_L g5635 ( 
.A(n_4894),
.B(n_4426),
.Y(n_5635)
);

BUFx6f_ASAP7_75t_L g5636 ( 
.A(n_4263),
.Y(n_5636)
);

INVx2_ASAP7_75t_L g5637 ( 
.A(n_4615),
.Y(n_5637)
);

OAI22xp33_ASAP7_75t_L g5638 ( 
.A1(n_4739),
.A2(n_4754),
.B1(n_4791),
.B2(n_4829),
.Y(n_5638)
);

INVx5_ASAP7_75t_L g5639 ( 
.A(n_4657),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_4620),
.Y(n_5640)
);

INVx2_ASAP7_75t_L g5641 ( 
.A(n_4620),
.Y(n_5641)
);

OR2x2_ASAP7_75t_L g5642 ( 
.A(n_4911),
.B(n_4395),
.Y(n_5642)
);

AOI22xp33_ASAP7_75t_L g5643 ( 
.A1(n_4168),
.A2(n_4953),
.B1(n_4126),
.B2(n_4855),
.Y(n_5643)
);

AND2x2_ASAP7_75t_SL g5644 ( 
.A(n_4863),
.B(n_5022),
.Y(n_5644)
);

OR2x2_ASAP7_75t_L g5645 ( 
.A(n_4911),
.B(n_4395),
.Y(n_5645)
);

AOI22xp5_ASAP7_75t_L g5646 ( 
.A1(n_4739),
.A2(n_4754),
.B1(n_4766),
.B2(n_4630),
.Y(n_5646)
);

AOI22xp33_ASAP7_75t_L g5647 ( 
.A1(n_4168),
.A2(n_4953),
.B1(n_4126),
.B2(n_4766),
.Y(n_5647)
);

NAND2x1_ASAP7_75t_L g5648 ( 
.A(n_5061),
.B(n_4657),
.Y(n_5648)
);

INVx2_ASAP7_75t_L g5649 ( 
.A(n_4636),
.Y(n_5649)
);

OAI22xp5_ASAP7_75t_L g5650 ( 
.A1(n_5063),
.A2(n_4844),
.B1(n_4142),
.B2(n_4154),
.Y(n_5650)
);

CKINVDCx5p33_ASAP7_75t_R g5651 ( 
.A(n_4927),
.Y(n_5651)
);

INVx1_ASAP7_75t_SL g5652 ( 
.A(n_5069),
.Y(n_5652)
);

BUFx8_ASAP7_75t_L g5653 ( 
.A(n_4293),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_4636),
.Y(n_5654)
);

NOR2xp67_ASAP7_75t_L g5655 ( 
.A(n_4151),
.B(n_4276),
.Y(n_5655)
);

AND2x4_ASAP7_75t_L g5656 ( 
.A(n_4894),
.B(n_4426),
.Y(n_5656)
);

INVxp67_ASAP7_75t_L g5657 ( 
.A(n_4651),
.Y(n_5657)
);

CKINVDCx8_ASAP7_75t_R g5658 ( 
.A(n_4151),
.Y(n_5658)
);

AO22x1_ASAP7_75t_L g5659 ( 
.A1(n_4334),
.A2(n_4437),
.B1(n_4921),
.B2(n_4361),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_4669),
.Y(n_5660)
);

INVx1_ASAP7_75t_SL g5661 ( 
.A(n_5069),
.Y(n_5661)
);

AOI22xp5_ASAP7_75t_L g5662 ( 
.A1(n_4791),
.A2(n_4829),
.B1(n_4962),
.B2(n_4768),
.Y(n_5662)
);

AOI221xp5_ASAP7_75t_L g5663 ( 
.A1(n_4642),
.A2(n_4692),
.B1(n_4714),
.B2(n_4680),
.C(n_4654),
.Y(n_5663)
);

INVx2_ASAP7_75t_L g5664 ( 
.A(n_4669),
.Y(n_5664)
);

BUFx12f_ASAP7_75t_L g5665 ( 
.A(n_4690),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_4672),
.Y(n_5666)
);

INVxp67_ASAP7_75t_L g5667 ( 
.A(n_4651),
.Y(n_5667)
);

AOI21x1_ASAP7_75t_L g5668 ( 
.A1(n_4424),
.A2(n_4430),
.B(n_4238),
.Y(n_5668)
);

BUFx2_ASAP7_75t_L g5669 ( 
.A(n_5029),
.Y(n_5669)
);

OR2x6_ASAP7_75t_SL g5670 ( 
.A(n_4403),
.B(n_4443),
.Y(n_5670)
);

OAI221xp5_ASAP7_75t_L g5671 ( 
.A1(n_4668),
.A2(n_4768),
.B1(n_4511),
.B2(n_4488),
.C(n_4984),
.Y(n_5671)
);

AOI22xp33_ASAP7_75t_L g5672 ( 
.A1(n_4962),
.A2(n_4805),
.B1(n_4293),
.B2(n_4393),
.Y(n_5672)
);

AOI22xp5_ASAP7_75t_L g5673 ( 
.A1(n_4711),
.A2(n_4712),
.B1(n_4717),
.B2(n_4735),
.Y(n_5673)
);

AOI22xp33_ASAP7_75t_L g5674 ( 
.A1(n_4293),
.A2(n_4319),
.B1(n_4400),
.B2(n_4393),
.Y(n_5674)
);

CKINVDCx5p33_ASAP7_75t_R g5675 ( 
.A(n_4965),
.Y(n_5675)
);

OAI22xp5_ASAP7_75t_L g5676 ( 
.A1(n_5063),
.A2(n_4844),
.B1(n_4142),
.B2(n_4154),
.Y(n_5676)
);

INVx4_ASAP7_75t_L g5677 ( 
.A(n_4293),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_4691),
.B(n_4596),
.Y(n_5678)
);

AND2x6_ASAP7_75t_L g5679 ( 
.A(n_4293),
.B(n_4319),
.Y(n_5679)
);

INVx1_ASAP7_75t_SL g5680 ( 
.A(n_5016),
.Y(n_5680)
);

CKINVDCx20_ASAP7_75t_R g5681 ( 
.A(n_4978),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_L g5682 ( 
.A(n_4691),
.B(n_4899),
.Y(n_5682)
);

AOI22xp33_ASAP7_75t_L g5683 ( 
.A1(n_4293),
.A2(n_4319),
.B1(n_4400),
.B2(n_4393),
.Y(n_5683)
);

OAI22xp5_ASAP7_75t_L g5684 ( 
.A1(n_4139),
.A2(n_4161),
.B1(n_4169),
.B2(n_4160),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_4672),
.Y(n_5685)
);

OAI22xp5_ASAP7_75t_L g5686 ( 
.A1(n_4139),
.A2(n_4161),
.B1(n_4169),
.B2(n_4160),
.Y(n_5686)
);

AOI22xp5_ASAP7_75t_L g5687 ( 
.A1(n_4711),
.A2(n_4712),
.B1(n_4717),
.B2(n_4668),
.Y(n_5687)
);

AOI22xp5_ASAP7_75t_L g5688 ( 
.A1(n_4171),
.A2(n_4174),
.B1(n_4179),
.B2(n_4173),
.Y(n_5688)
);

NAND2xp5_ASAP7_75t_L g5689 ( 
.A(n_4899),
.B(n_4916),
.Y(n_5689)
);

AOI22xp5_ASAP7_75t_L g5690 ( 
.A1(n_4171),
.A2(n_4174),
.B1(n_4179),
.B2(n_4173),
.Y(n_5690)
);

INVx5_ASAP7_75t_L g5691 ( 
.A(n_4657),
.Y(n_5691)
);

OAI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_4769),
.A2(n_4082),
.B1(n_4153),
.B2(n_4092),
.Y(n_5692)
);

BUFx2_ASAP7_75t_L g5693 ( 
.A(n_4908),
.Y(n_5693)
);

AOI22xp33_ASAP7_75t_L g5694 ( 
.A1(n_4319),
.A2(n_4400),
.B1(n_4423),
.B2(n_4393),
.Y(n_5694)
);

OR2x6_ASAP7_75t_L g5695 ( 
.A(n_4816),
.B(n_4833),
.Y(n_5695)
);

OAI22xp33_ASAP7_75t_L g5696 ( 
.A1(n_4769),
.A2(n_4092),
.B1(n_4153),
.B2(n_4319),
.Y(n_5696)
);

AND2x6_ASAP7_75t_L g5697 ( 
.A(n_4319),
.B(n_4393),
.Y(n_5697)
);

AOI22xp33_ASAP7_75t_L g5698 ( 
.A1(n_4393),
.A2(n_4423),
.B1(n_4429),
.B2(n_4400),
.Y(n_5698)
);

NOR2xp33_ASAP7_75t_L g5699 ( 
.A(n_4608),
.B(n_4959),
.Y(n_5699)
);

INVx4_ASAP7_75t_L g5700 ( 
.A(n_4400),
.Y(n_5700)
);

NAND2xp5_ASAP7_75t_L g5701 ( 
.A(n_4916),
.B(n_4436),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_4687),
.Y(n_5702)
);

OR2x6_ASAP7_75t_L g5703 ( 
.A(n_4833),
.B(n_4835),
.Y(n_5703)
);

OR2x6_ASAP7_75t_SL g5704 ( 
.A(n_4403),
.B(n_4443),
.Y(n_5704)
);

INVx2_ASAP7_75t_L g5705 ( 
.A(n_4687),
.Y(n_5705)
);

AOI22xp33_ASAP7_75t_L g5706 ( 
.A1(n_4400),
.A2(n_4429),
.B1(n_4452),
.B2(n_4423),
.Y(n_5706)
);

INVx4_ASAP7_75t_L g5707 ( 
.A(n_4423),
.Y(n_5707)
);

CKINVDCx16_ASAP7_75t_R g5708 ( 
.A(n_4893),
.Y(n_5708)
);

OAI22xp5_ASAP7_75t_L g5709 ( 
.A1(n_4185),
.A2(n_4187),
.B1(n_4192),
.B2(n_4191),
.Y(n_5709)
);

CKINVDCx5p33_ASAP7_75t_R g5710 ( 
.A(n_4810),
.Y(n_5710)
);

NOR2xp33_ASAP7_75t_SL g5711 ( 
.A(n_4943),
.B(n_4575),
.Y(n_5711)
);

NAND2xp5_ASAP7_75t_L g5712 ( 
.A(n_4432),
.B(n_4898),
.Y(n_5712)
);

INVx1_ASAP7_75t_SL g5713 ( 
.A(n_5016),
.Y(n_5713)
);

OAI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_4092),
.A2(n_4429),
.B1(n_4452),
.B2(n_4423),
.Y(n_5714)
);

INVx1_ASAP7_75t_SL g5715 ( 
.A(n_5056),
.Y(n_5715)
);

OAI222xp33_ASAP7_75t_L g5716 ( 
.A1(n_4616),
.A2(n_4624),
.B1(n_4640),
.B2(n_4670),
.C1(n_4652),
.C2(n_4618),
.Y(n_5716)
);

NAND2xp5_ASAP7_75t_L g5717 ( 
.A(n_4432),
.B(n_4898),
.Y(n_5717)
);

OR2x2_ASAP7_75t_L g5718 ( 
.A(n_4470),
.B(n_4472),
.Y(n_5718)
);

CKINVDCx8_ASAP7_75t_R g5719 ( 
.A(n_4151),
.Y(n_5719)
);

OR2x6_ASAP7_75t_L g5720 ( 
.A(n_4835),
.B(n_4575),
.Y(n_5720)
);

BUFx2_ASAP7_75t_L g5721 ( 
.A(n_4908),
.Y(n_5721)
);

AOI22xp33_ASAP7_75t_L g5722 ( 
.A1(n_4429),
.A2(n_4467),
.B1(n_4545),
.B2(n_4452),
.Y(n_5722)
);

NAND2xp5_ASAP7_75t_L g5723 ( 
.A(n_4358),
.B(n_4956),
.Y(n_5723)
);

AOI22xp5_ASAP7_75t_L g5724 ( 
.A1(n_4185),
.A2(n_4191),
.B1(n_4192),
.B2(n_4187),
.Y(n_5724)
);

CKINVDCx20_ASAP7_75t_R g5725 ( 
.A(n_4957),
.Y(n_5725)
);

AOI21xp5_ASAP7_75t_SL g5726 ( 
.A1(n_5011),
.A2(n_4957),
.B(n_5074),
.Y(n_5726)
);

INVx1_ASAP7_75t_SL g5727 ( 
.A(n_5056),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_4694),
.Y(n_5728)
);

AOI22xp5_ASAP7_75t_L g5729 ( 
.A1(n_4200),
.A2(n_4212),
.B1(n_4213),
.B2(n_4202),
.Y(n_5729)
);

BUFx12f_ASAP7_75t_L g5730 ( 
.A(n_4690),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_SL g5731 ( 
.A(n_4929),
.B(n_4995),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_4694),
.Y(n_5732)
);

INVx2_ASAP7_75t_L g5733 ( 
.A(n_4696),
.Y(n_5733)
);

AO22x1_ASAP7_75t_L g5734 ( 
.A1(n_4334),
.A2(n_4437),
.B1(n_4921),
.B2(n_4226),
.Y(n_5734)
);

INVx4_ASAP7_75t_L g5735 ( 
.A(n_4452),
.Y(n_5735)
);

NAND2xp33_ASAP7_75t_SL g5736 ( 
.A(n_4334),
.B(n_4437),
.Y(n_5736)
);

OAI22xp5_ASAP7_75t_L g5737 ( 
.A1(n_4200),
.A2(n_4212),
.B1(n_4213),
.B2(n_4202),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_4696),
.Y(n_5738)
);

INVx4_ASAP7_75t_L g5739 ( 
.A(n_4467),
.Y(n_5739)
);

BUFx6f_ASAP7_75t_SL g5740 ( 
.A(n_4690),
.Y(n_5740)
);

AND2x2_ASAP7_75t_SL g5741 ( 
.A(n_4863),
.B(n_4979),
.Y(n_5741)
);

CKINVDCx8_ASAP7_75t_R g5742 ( 
.A(n_4151),
.Y(n_5742)
);

AOI22xp5_ASAP7_75t_L g5743 ( 
.A1(n_4222),
.A2(n_4228),
.B1(n_4229),
.B2(n_4225),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_4898),
.B(n_4909),
.Y(n_5744)
);

INVx2_ASAP7_75t_L g5745 ( 
.A(n_4705),
.Y(n_5745)
);

NAND2xp5_ASAP7_75t_SL g5746 ( 
.A(n_4750),
.B(n_5052),
.Y(n_5746)
);

NOR2xp33_ASAP7_75t_L g5747 ( 
.A(n_4959),
.B(n_4222),
.Y(n_5747)
);

CKINVDCx11_ASAP7_75t_R g5748 ( 
.A(n_4827),
.Y(n_5748)
);

BUFx8_ASAP7_75t_SL g5749 ( 
.A(n_4376),
.Y(n_5749)
);

O2A1O1Ixp33_ASAP7_75t_L g5750 ( 
.A1(n_4521),
.A2(n_4488),
.B(n_4726),
.C(n_4509),
.Y(n_5750)
);

AND2x2_ASAP7_75t_L g5751 ( 
.A(n_5007),
.B(n_4910),
.Y(n_5751)
);

INVx1_ASAP7_75t_SL g5752 ( 
.A(n_5056),
.Y(n_5752)
);

AOI22xp5_ASAP7_75t_L g5753 ( 
.A1(n_4225),
.A2(n_4228),
.B1(n_4257),
.B2(n_4229),
.Y(n_5753)
);

NOR2xp33_ASAP7_75t_L g5754 ( 
.A(n_4257),
.B(n_4264),
.Y(n_5754)
);

AOI22xp5_ASAP7_75t_L g5755 ( 
.A1(n_4264),
.A2(n_4275),
.B1(n_4279),
.B2(n_4272),
.Y(n_5755)
);

BUFx4f_ASAP7_75t_SL g5756 ( 
.A(n_4827),
.Y(n_5756)
);

NAND2xp5_ASAP7_75t_L g5757 ( 
.A(n_4926),
.B(n_4501),
.Y(n_5757)
);

AOI21xp5_ASAP7_75t_L g5758 ( 
.A1(n_4658),
.A2(n_4662),
.B(n_4660),
.Y(n_5758)
);

AOI22xp33_ASAP7_75t_L g5759 ( 
.A1(n_4467),
.A2(n_4588),
.B1(n_4612),
.B2(n_4545),
.Y(n_5759)
);

OR2x2_ASAP7_75t_L g5760 ( 
.A(n_4470),
.B(n_4472),
.Y(n_5760)
);

OR2x2_ASAP7_75t_L g5761 ( 
.A(n_4482),
.B(n_4483),
.Y(n_5761)
);

INVx5_ASAP7_75t_L g5762 ( 
.A(n_4657),
.Y(n_5762)
);

NOR2xp33_ASAP7_75t_L g5763 ( 
.A(n_4272),
.B(n_4275),
.Y(n_5763)
);

O2A1O1Ixp33_ASAP7_75t_SL g5764 ( 
.A1(n_4834),
.A2(n_4966),
.B(n_4928),
.C(n_5032),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_L g5765 ( 
.A(n_4956),
.B(n_4279),
.Y(n_5765)
);

NAND2xp5_ASAP7_75t_L g5766 ( 
.A(n_4290),
.B(n_4292),
.Y(n_5766)
);

BUFx6f_ASAP7_75t_L g5767 ( 
.A(n_4467),
.Y(n_5767)
);

INVx5_ASAP7_75t_L g5768 ( 
.A(n_4657),
.Y(n_5768)
);

INVx1_ASAP7_75t_SL g5769 ( 
.A(n_4963),
.Y(n_5769)
);

AOI222xp33_ASAP7_75t_L g5770 ( 
.A1(n_4290),
.A2(n_4305),
.B1(n_4292),
.B2(n_4315),
.C1(n_4307),
.C2(n_4294),
.Y(n_5770)
);

INVxp67_ASAP7_75t_L g5771 ( 
.A(n_4862),
.Y(n_5771)
);

OAI22xp5_ASAP7_75t_L g5772 ( 
.A1(n_4294),
.A2(n_4307),
.B1(n_4315),
.B2(n_4305),
.Y(n_5772)
);

O2A1O1Ixp5_ASAP7_75t_L g5773 ( 
.A1(n_4532),
.A2(n_4947),
.B(n_4637),
.C(n_5024),
.Y(n_5773)
);

BUFx6f_ASAP7_75t_L g5774 ( 
.A(n_4467),
.Y(n_5774)
);

BUFx6f_ASAP7_75t_L g5775 ( 
.A(n_4545),
.Y(n_5775)
);

AOI22xp33_ASAP7_75t_L g5776 ( 
.A1(n_4545),
.A2(n_4612),
.B1(n_4588),
.B2(n_4361),
.Y(n_5776)
);

OR2x6_ASAP7_75t_SL g5777 ( 
.A(n_4482),
.B(n_4483),
.Y(n_5777)
);

AOI22xp5_ASAP7_75t_L g5778 ( 
.A1(n_4318),
.A2(n_4325),
.B1(n_4340),
.B2(n_4326),
.Y(n_5778)
);

OAI21xp5_ASAP7_75t_L g5779 ( 
.A1(n_4196),
.A2(n_4532),
.B(n_4637),
.Y(n_5779)
);

AOI221xp5_ASAP7_75t_L g5780 ( 
.A1(n_4724),
.A2(n_4501),
.B1(n_4743),
.B2(n_4508),
.C(n_4500),
.Y(n_5780)
);

CKINVDCx8_ASAP7_75t_R g5781 ( 
.A(n_4276),
.Y(n_5781)
);

AOI22xp5_ASAP7_75t_L g5782 ( 
.A1(n_4318),
.A2(n_4325),
.B1(n_4340),
.B2(n_4326),
.Y(n_5782)
);

BUFx12f_ASAP7_75t_L g5783 ( 
.A(n_4690),
.Y(n_5783)
);

AOI21xp5_ASAP7_75t_L g5784 ( 
.A1(n_5288),
.A2(n_4430),
.B(n_4678),
.Y(n_5784)
);

BUFx2_ASAP7_75t_L g5785 ( 
.A(n_5113),
.Y(n_5785)
);

CKINVDCx5p33_ASAP7_75t_R g5786 ( 
.A(n_5122),
.Y(n_5786)
);

NAND2xp5_ASAP7_75t_L g5787 ( 
.A(n_5176),
.B(n_4724),
.Y(n_5787)
);

AOI22xp5_ASAP7_75t_L g5788 ( 
.A1(n_5147),
.A2(n_4977),
.B1(n_4775),
.B2(n_4786),
.Y(n_5788)
);

NAND3xp33_ASAP7_75t_L g5789 ( 
.A(n_5137),
.B(n_4438),
.C(n_4435),
.Y(n_5789)
);

INVx3_ASAP7_75t_L g5790 ( 
.A(n_5099),
.Y(n_5790)
);

INVx2_ASAP7_75t_SL g5791 ( 
.A(n_5262),
.Y(n_5791)
);

NOR2xp33_ASAP7_75t_L g5792 ( 
.A(n_5181),
.B(n_4998),
.Y(n_5792)
);

O2A1O1Ixp33_ASAP7_75t_SL g5793 ( 
.A1(n_5250),
.A2(n_4888),
.B(n_4912),
.C(n_4906),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_5099),
.Y(n_5794)
);

HB1xp67_ASAP7_75t_L g5795 ( 
.A(n_5431),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_5099),
.Y(n_5796)
);

INVx1_ASAP7_75t_L g5797 ( 
.A(n_5599),
.Y(n_5797)
);

INVx8_ASAP7_75t_L g5798 ( 
.A(n_5170),
.Y(n_5798)
);

NAND2xp5_ASAP7_75t_L g5799 ( 
.A(n_5176),
.B(n_4374),
.Y(n_5799)
);

BUFx3_ASAP7_75t_L g5800 ( 
.A(n_5648),
.Y(n_5800)
);

OAI22xp5_ASAP7_75t_L g5801 ( 
.A1(n_5230),
.A2(n_4616),
.B1(n_4624),
.B2(n_4618),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5599),
.Y(n_5802)
);

BUFx10_ASAP7_75t_L g5803 ( 
.A(n_5740),
.Y(n_5803)
);

BUFx3_ASAP7_75t_L g5804 ( 
.A(n_5648),
.Y(n_5804)
);

INVx4_ASAP7_75t_L g5805 ( 
.A(n_5115),
.Y(n_5805)
);

OAI21xp33_ASAP7_75t_L g5806 ( 
.A1(n_5225),
.A2(n_4438),
.B(n_4435),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5599),
.Y(n_5807)
);

INVx2_ASAP7_75t_L g5808 ( 
.A(n_5099),
.Y(n_5808)
);

BUFx12f_ASAP7_75t_L g5809 ( 
.A(n_5273),
.Y(n_5809)
);

INVx1_ASAP7_75t_SL g5810 ( 
.A(n_5452),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5599),
.Y(n_5811)
);

INVx5_ASAP7_75t_L g5812 ( 
.A(n_5262),
.Y(n_5812)
);

NAND2xp5_ASAP7_75t_L g5813 ( 
.A(n_5176),
.B(n_4374),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5109),
.Y(n_5814)
);

NAND2xp5_ASAP7_75t_L g5815 ( 
.A(n_5181),
.B(n_4389),
.Y(n_5815)
);

AND2x4_ASAP7_75t_L g5816 ( 
.A(n_5196),
.B(n_4581),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5617),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5617),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_5122),
.Y(n_5819)
);

INVx2_ASAP7_75t_SL g5820 ( 
.A(n_5262),
.Y(n_5820)
);

AND2x4_ASAP7_75t_L g5821 ( 
.A(n_5196),
.B(n_4581),
.Y(n_5821)
);

BUFx2_ASAP7_75t_L g5822 ( 
.A(n_5113),
.Y(n_5822)
);

HB1xp67_ASAP7_75t_L g5823 ( 
.A(n_5431),
.Y(n_5823)
);

AOI21xp5_ASAP7_75t_L g5824 ( 
.A1(n_5288),
.A2(n_4681),
.B(n_4678),
.Y(n_5824)
);

OA21x2_ASAP7_75t_L g5825 ( 
.A1(n_5531),
.A2(n_4846),
.B(n_4890),
.Y(n_5825)
);

NAND2xp5_ASAP7_75t_SL g5826 ( 
.A(n_5140),
.B(n_4972),
.Y(n_5826)
);

NAND2xp5_ASAP7_75t_L g5827 ( 
.A(n_5181),
.B(n_4389),
.Y(n_5827)
);

CKINVDCx8_ASAP7_75t_R g5828 ( 
.A(n_5398),
.Y(n_5828)
);

INVx3_ASAP7_75t_L g5829 ( 
.A(n_5109),
.Y(n_5829)
);

BUFx6f_ASAP7_75t_L g5830 ( 
.A(n_5094),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_5617),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5617),
.Y(n_5832)
);

OAI22xp5_ASAP7_75t_L g5833 ( 
.A1(n_5230),
.A2(n_4652),
.B1(n_4670),
.B2(n_4640),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5632),
.Y(n_5834)
);

BUFx3_ASAP7_75t_L g5835 ( 
.A(n_5648),
.Y(n_5835)
);

HB1xp67_ASAP7_75t_L g5836 ( 
.A(n_5431),
.Y(n_5836)
);

AOI21xp5_ASAP7_75t_SL g5837 ( 
.A1(n_5137),
.A2(n_4398),
.B(n_4226),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5632),
.Y(n_5838)
);

OAI21xp33_ASAP7_75t_L g5839 ( 
.A1(n_5225),
.A2(n_5147),
.B(n_5230),
.Y(n_5839)
);

BUFx12f_ASAP7_75t_L g5840 ( 
.A(n_5273),
.Y(n_5840)
);

AOI222xp33_ASAP7_75t_L g5841 ( 
.A1(n_5184),
.A2(n_5201),
.B1(n_5234),
.B2(n_5140),
.C1(n_5161),
.C2(n_5353),
.Y(n_5841)
);

INVx2_ASAP7_75t_SL g5842 ( 
.A(n_5262),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5632),
.Y(n_5843)
);

BUFx3_ASAP7_75t_L g5844 ( 
.A(n_5749),
.Y(n_5844)
);

AOI21xp5_ASAP7_75t_L g5845 ( 
.A1(n_5277),
.A2(n_4683),
.B(n_4681),
.Y(n_5845)
);

BUFx8_ASAP7_75t_L g5846 ( 
.A(n_5115),
.Y(n_5846)
);

OAI21xp5_ASAP7_75t_L g5847 ( 
.A1(n_5186),
.A2(n_4458),
.B(n_4442),
.Y(n_5847)
);

INVx4_ASAP7_75t_L g5848 ( 
.A(n_5115),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5632),
.Y(n_5849)
);

AO21x1_ASAP7_75t_L g5850 ( 
.A1(n_5551),
.A2(n_4580),
.B(n_4500),
.Y(n_5850)
);

NAND2xp5_ASAP7_75t_L g5851 ( 
.A(n_5545),
.B(n_4459),
.Y(n_5851)
);

BUFx3_ASAP7_75t_L g5852 ( 
.A(n_5749),
.Y(n_5852)
);

BUFx6f_ASAP7_75t_L g5853 ( 
.A(n_5094),
.Y(n_5853)
);

AOI21xp5_ASAP7_75t_L g5854 ( 
.A1(n_5277),
.A2(n_4704),
.B(n_4683),
.Y(n_5854)
);

NAND2xp5_ASAP7_75t_L g5855 ( 
.A(n_5545),
.B(n_4459),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_L g5856 ( 
.A(n_5545),
.B(n_4504),
.Y(n_5856)
);

OAI22xp5_ASAP7_75t_L g5857 ( 
.A1(n_5275),
.A2(n_4675),
.B1(n_4633),
.B2(n_4565),
.Y(n_5857)
);

INVx2_ASAP7_75t_L g5858 ( 
.A(n_5109),
.Y(n_5858)
);

AOI22xp5_ASAP7_75t_L g5859 ( 
.A1(n_5171),
.A2(n_4977),
.B1(n_4788),
.B2(n_4756),
.Y(n_5859)
);

NOR2xp33_ASAP7_75t_L g5860 ( 
.A(n_5419),
.B(n_4998),
.Y(n_5860)
);

NAND2x1p5_ASAP7_75t_L g5861 ( 
.A(n_5141),
.B(n_4276),
.Y(n_5861)
);

BUFx3_ASAP7_75t_L g5862 ( 
.A(n_5098),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5637),
.Y(n_5863)
);

NAND2xp5_ASAP7_75t_L g5864 ( 
.A(n_5549),
.B(n_4504),
.Y(n_5864)
);

INVx4_ASAP7_75t_L g5865 ( 
.A(n_5115),
.Y(n_5865)
);

BUFx6f_ASAP7_75t_L g5866 ( 
.A(n_5094),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5637),
.Y(n_5867)
);

OAI21xp5_ASAP7_75t_L g5868 ( 
.A1(n_5186),
.A2(n_4458),
.B(n_4442),
.Y(n_5868)
);

INVx2_ASAP7_75t_SL g5869 ( 
.A(n_5262),
.Y(n_5869)
);

CKINVDCx5p33_ASAP7_75t_R g5870 ( 
.A(n_5135),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_5549),
.B(n_4519),
.Y(n_5871)
);

AOI21xp5_ASAP7_75t_L g5872 ( 
.A1(n_5300),
.A2(n_5210),
.B(n_5174),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5637),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5109),
.Y(n_5874)
);

INVx2_ASAP7_75t_L g5875 ( 
.A(n_5119),
.Y(n_5875)
);

NAND2xp5_ASAP7_75t_L g5876 ( 
.A(n_5549),
.B(n_4519),
.Y(n_5876)
);

CKINVDCx8_ASAP7_75t_R g5877 ( 
.A(n_5398),
.Y(n_5877)
);

AND2x4_ASAP7_75t_L g5878 ( 
.A(n_5196),
.B(n_4701),
.Y(n_5878)
);

AOI21xp5_ASAP7_75t_L g5879 ( 
.A1(n_5300),
.A2(n_4709),
.B(n_4704),
.Y(n_5879)
);

BUFx6f_ASAP7_75t_L g5880 ( 
.A(n_5094),
.Y(n_5880)
);

O2A1O1Ixp5_ASAP7_75t_L g5881 ( 
.A1(n_5161),
.A2(n_4460),
.B(n_4489),
.C(n_4487),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5637),
.Y(n_5882)
);

BUFx3_ASAP7_75t_L g5883 ( 
.A(n_5098),
.Y(n_5883)
);

NAND2x1p5_ASAP7_75t_L g5884 ( 
.A(n_5141),
.B(n_4276),
.Y(n_5884)
);

INVx1_ASAP7_75t_SL g5885 ( 
.A(n_5452),
.Y(n_5885)
);

CKINVDCx5p33_ASAP7_75t_R g5886 ( 
.A(n_5135),
.Y(n_5886)
);

INVx5_ASAP7_75t_L g5887 ( 
.A(n_5262),
.Y(n_5887)
);

INVx3_ASAP7_75t_L g5888 ( 
.A(n_5119),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_SL g5889 ( 
.A(n_5225),
.B(n_4972),
.Y(n_5889)
);

AOI221xp5_ASAP7_75t_L g5890 ( 
.A1(n_5178),
.A2(n_4508),
.B1(n_4495),
.B2(n_4743),
.C(n_4831),
.Y(n_5890)
);

NOR2xp33_ASAP7_75t_L g5891 ( 
.A(n_5419),
.B(n_5000),
.Y(n_5891)
);

OR2x2_ASAP7_75t_L g5892 ( 
.A(n_5712),
.B(n_4495),
.Y(n_5892)
);

NAND3xp33_ASAP7_75t_L g5893 ( 
.A(n_5186),
.B(n_4487),
.C(n_4460),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5640),
.Y(n_5894)
);

A2O1A1Ixp33_ASAP7_75t_L g5895 ( 
.A1(n_5178),
.A2(n_4494),
.B(n_4498),
.C(n_4489),
.Y(n_5895)
);

AOI21xp33_ASAP7_75t_SL g5896 ( 
.A1(n_5209),
.A2(n_4351),
.B(n_4250),
.Y(n_5896)
);

NOR2xp33_ASAP7_75t_L g5897 ( 
.A(n_5232),
.B(n_5000),
.Y(n_5897)
);

A2O1A1Ixp33_ASAP7_75t_L g5898 ( 
.A1(n_5178),
.A2(n_4498),
.B(n_4499),
.C(n_4494),
.Y(n_5898)
);

BUFx10_ASAP7_75t_L g5899 ( 
.A(n_5740),
.Y(n_5899)
);

NAND2x1p5_ASAP7_75t_L g5900 ( 
.A(n_5141),
.B(n_4276),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5640),
.Y(n_5901)
);

AOI22xp33_ASAP7_75t_L g5902 ( 
.A1(n_5171),
.A2(n_4831),
.B1(n_4588),
.B2(n_4612),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5640),
.Y(n_5903)
);

INVx2_ASAP7_75t_L g5904 ( 
.A(n_5119),
.Y(n_5904)
);

CKINVDCx5p33_ASAP7_75t_R g5905 ( 
.A(n_5134),
.Y(n_5905)
);

OA21x2_ASAP7_75t_L g5906 ( 
.A1(n_5531),
.A2(n_4846),
.B(n_4523),
.Y(n_5906)
);

NAND2xp5_ASAP7_75t_SL g5907 ( 
.A(n_5581),
.B(n_4690),
.Y(n_5907)
);

BUFx2_ASAP7_75t_L g5908 ( 
.A(n_5113),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5640),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5641),
.Y(n_5910)
);

INVx3_ASAP7_75t_SL g5911 ( 
.A(n_5731),
.Y(n_5911)
);

O2A1O1Ixp33_ASAP7_75t_L g5912 ( 
.A1(n_5250),
.A2(n_4849),
.B(n_4839),
.C(n_4523),
.Y(n_5912)
);

A2O1A1Ixp33_ASAP7_75t_SL g5913 ( 
.A1(n_5521),
.A2(n_4990),
.B(n_4875),
.C(n_4903),
.Y(n_5913)
);

NAND2xp5_ASAP7_75t_L g5914 ( 
.A(n_5218),
.B(n_4723),
.Y(n_5914)
);

CKINVDCx16_ASAP7_75t_R g5915 ( 
.A(n_5456),
.Y(n_5915)
);

NAND2xp5_ASAP7_75t_L g5916 ( 
.A(n_5218),
.B(n_4723),
.Y(n_5916)
);

AOI21xp5_ASAP7_75t_L g5917 ( 
.A1(n_5210),
.A2(n_4720),
.B(n_4709),
.Y(n_5917)
);

CKINVDCx5p33_ASAP7_75t_R g5918 ( 
.A(n_5134),
.Y(n_5918)
);

INVx4_ASAP7_75t_L g5919 ( 
.A(n_5136),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5641),
.Y(n_5920)
);

A2O1A1Ixp33_ASAP7_75t_L g5921 ( 
.A1(n_5581),
.A2(n_4499),
.B(n_4750),
.C(n_4889),
.Y(n_5921)
);

INVx1_ASAP7_75t_L g5922 ( 
.A(n_5641),
.Y(n_5922)
);

AND2x2_ASAP7_75t_SL g5923 ( 
.A(n_5377),
.B(n_4979),
.Y(n_5923)
);

BUFx3_ASAP7_75t_L g5924 ( 
.A(n_5098),
.Y(n_5924)
);

HB1xp67_ASAP7_75t_L g5925 ( 
.A(n_5443),
.Y(n_5925)
);

NAND2xp5_ASAP7_75t_L g5926 ( 
.A(n_5218),
.B(n_4729),
.Y(n_5926)
);

AOI21xp5_ASAP7_75t_L g5927 ( 
.A1(n_5131),
.A2(n_4733),
.B(n_4720),
.Y(n_5927)
);

NAND2xp5_ASAP7_75t_L g5928 ( 
.A(n_5506),
.B(n_4729),
.Y(n_5928)
);

INVxp67_ASAP7_75t_SL g5929 ( 
.A(n_5364),
.Y(n_5929)
);

OR2x2_ASAP7_75t_L g5930 ( 
.A(n_5712),
.B(n_4963),
.Y(n_5930)
);

INVx5_ASAP7_75t_L g5931 ( 
.A(n_5262),
.Y(n_5931)
);

NOR2xp33_ASAP7_75t_L g5932 ( 
.A(n_5232),
.B(n_5004),
.Y(n_5932)
);

BUFx6f_ASAP7_75t_L g5933 ( 
.A(n_5094),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5641),
.Y(n_5934)
);

AOI21xp5_ASAP7_75t_L g5935 ( 
.A1(n_5131),
.A2(n_4733),
.B(n_4889),
.Y(n_5935)
);

AOI21xp5_ASAP7_75t_L g5936 ( 
.A1(n_5174),
.A2(n_4767),
.B(n_4753),
.Y(n_5936)
);

INVx2_ASAP7_75t_SL g5937 ( 
.A(n_5262),
.Y(n_5937)
);

INVx1_ASAP7_75t_SL g5938 ( 
.A(n_5452),
.Y(n_5938)
);

BUFx12f_ASAP7_75t_L g5939 ( 
.A(n_5168),
.Y(n_5939)
);

INVx1_ASAP7_75t_SL g5940 ( 
.A(n_5470),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5649),
.Y(n_5941)
);

NAND2xp5_ASAP7_75t_L g5942 ( 
.A(n_5506),
.B(n_4760),
.Y(n_5942)
);

NAND2x1p5_ASAP7_75t_L g5943 ( 
.A(n_5141),
.B(n_4276),
.Y(n_5943)
);

NAND2xp5_ASAP7_75t_L g5944 ( 
.A(n_5528),
.B(n_4760),
.Y(n_5944)
);

BUFx3_ASAP7_75t_L g5945 ( 
.A(n_5098),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5649),
.Y(n_5946)
);

INVx1_ASAP7_75t_SL g5947 ( 
.A(n_5470),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5649),
.Y(n_5948)
);

INVx1_ASAP7_75t_L g5949 ( 
.A(n_5649),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_L g5950 ( 
.A(n_5528),
.B(n_4763),
.Y(n_5950)
);

OA21x2_ASAP7_75t_L g5951 ( 
.A1(n_5529),
.A2(n_4947),
.B(n_4601),
.Y(n_5951)
);

INVx1_ASAP7_75t_SL g5952 ( 
.A(n_5470),
.Y(n_5952)
);

BUFx8_ASAP7_75t_L g5953 ( 
.A(n_5136),
.Y(n_5953)
);

AOI22xp5_ASAP7_75t_L g5954 ( 
.A1(n_5171),
.A2(n_4588),
.B1(n_4612),
.B2(n_4545),
.Y(n_5954)
);

INVx2_ASAP7_75t_L g5955 ( 
.A(n_5119),
.Y(n_5955)
);

OR2x2_ASAP7_75t_L g5956 ( 
.A(n_5712),
.B(n_4963),
.Y(n_5956)
);

AOI21xp5_ASAP7_75t_L g5957 ( 
.A1(n_5529),
.A2(n_4767),
.B(n_4753),
.Y(n_5957)
);

INVx2_ASAP7_75t_SL g5958 ( 
.A(n_5408),
.Y(n_5958)
);

AND2x4_ASAP7_75t_L g5959 ( 
.A(n_5604),
.B(n_4567),
.Y(n_5959)
);

OAI22xp5_ASAP7_75t_SL g5960 ( 
.A1(n_5335),
.A2(n_4675),
.B1(n_4831),
.B2(n_4875),
.Y(n_5960)
);

HB1xp67_ASAP7_75t_L g5961 ( 
.A(n_5443),
.Y(n_5961)
);

BUFx3_ASAP7_75t_L g5962 ( 
.A(n_5106),
.Y(n_5962)
);

INVx3_ASAP7_75t_L g5963 ( 
.A(n_5129),
.Y(n_5963)
);

AOI21xp5_ASAP7_75t_L g5964 ( 
.A1(n_5254),
.A2(n_4796),
.B(n_5071),
.Y(n_5964)
);

NAND2xp5_ASAP7_75t_L g5965 ( 
.A(n_5253),
.B(n_4763),
.Y(n_5965)
);

OAI22xp5_ASAP7_75t_L g5966 ( 
.A1(n_5275),
.A2(n_5182),
.B1(n_5175),
.B2(n_5167),
.Y(n_5966)
);

INVx1_ASAP7_75t_SL g5967 ( 
.A(n_5329),
.Y(n_5967)
);

OAI21xp5_ASAP7_75t_L g5968 ( 
.A1(n_5390),
.A2(n_5204),
.B(n_5476),
.Y(n_5968)
);

AOI22xp33_ASAP7_75t_L g5969 ( 
.A1(n_5201),
.A2(n_4588),
.B1(n_4612),
.B2(n_4545),
.Y(n_5969)
);

INVx1_ASAP7_75t_SL g5970 ( 
.A(n_5329),
.Y(n_5970)
);

CKINVDCx6p67_ASAP7_75t_R g5971 ( 
.A(n_5505),
.Y(n_5971)
);

BUFx3_ASAP7_75t_L g5972 ( 
.A(n_5106),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5253),
.B(n_4765),
.Y(n_5973)
);

INVx3_ASAP7_75t_L g5974 ( 
.A(n_5129),
.Y(n_5974)
);

OAI22xp5_ASAP7_75t_L g5975 ( 
.A1(n_5275),
.A2(n_4633),
.B1(n_4565),
.B2(n_4342),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5496),
.B(n_4765),
.Y(n_5976)
);

INVx2_ASAP7_75t_SL g5977 ( 
.A(n_5408),
.Y(n_5977)
);

AOI21xp5_ASAP7_75t_L g5978 ( 
.A1(n_5254),
.A2(n_5306),
.B(n_5577),
.Y(n_5978)
);

HB1xp67_ASAP7_75t_L g5979 ( 
.A(n_5443),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5654),
.Y(n_5980)
);

O2A1O1Ixp33_ASAP7_75t_L g5981 ( 
.A1(n_5237),
.A2(n_4974),
.B(n_4987),
.C(n_4971),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5654),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_5496),
.B(n_4785),
.Y(n_5983)
);

AND3x1_ASAP7_75t_SL g5984 ( 
.A(n_5429),
.B(n_5006),
.C(n_5004),
.Y(n_5984)
);

INVx4_ASAP7_75t_L g5985 ( 
.A(n_5136),
.Y(n_5985)
);

AOI22xp5_ASAP7_75t_L g5986 ( 
.A1(n_5209),
.A2(n_4588),
.B1(n_4612),
.B2(n_4545),
.Y(n_5986)
);

HB1xp67_ASAP7_75t_L g5987 ( 
.A(n_5680),
.Y(n_5987)
);

NAND2xp5_ASAP7_75t_L g5988 ( 
.A(n_5373),
.B(n_4785),
.Y(n_5988)
);

NAND2xp5_ASAP7_75t_SL g5989 ( 
.A(n_5663),
.B(n_5014),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5373),
.B(n_4809),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5654),
.Y(n_5991)
);

OR2x2_ASAP7_75t_L g5992 ( 
.A(n_5717),
.B(n_4310),
.Y(n_5992)
);

BUFx6f_ASAP7_75t_L g5993 ( 
.A(n_5094),
.Y(n_5993)
);

BUFx6f_ASAP7_75t_L g5994 ( 
.A(n_5094),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5654),
.Y(n_5995)
);

AOI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_5306),
.A2(n_5073),
.B(n_5071),
.Y(n_5996)
);

BUFx3_ASAP7_75t_L g5997 ( 
.A(n_5106),
.Y(n_5997)
);

AOI22xp5_ASAP7_75t_L g5998 ( 
.A1(n_5212),
.A2(n_5182),
.B1(n_5353),
.B2(n_5175),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5660),
.Y(n_5999)
);

BUFx2_ASAP7_75t_L g6000 ( 
.A(n_5113),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5660),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5747),
.B(n_5365),
.Y(n_6002)
);

NAND2xp5_ASAP7_75t_L g6003 ( 
.A(n_5747),
.B(n_4809),
.Y(n_6003)
);

AND2x6_ASAP7_75t_L g6004 ( 
.A(n_5151),
.B(n_5057),
.Y(n_6004)
);

AOI21xp5_ASAP7_75t_L g6005 ( 
.A1(n_5577),
.A2(n_5073),
.B(n_4946),
.Y(n_6005)
);

INVx1_ASAP7_75t_SL g6006 ( 
.A(n_5329),
.Y(n_6006)
);

BUFx6f_ASAP7_75t_L g6007 ( 
.A(n_5094),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5660),
.Y(n_6008)
);

A2O1A1Ixp33_ASAP7_75t_L g6009 ( 
.A1(n_5663),
.A2(n_4587),
.B(n_4991),
.C(n_5052),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5660),
.Y(n_6010)
);

OR2x2_ASAP7_75t_L g6011 ( 
.A(n_5717),
.B(n_4310),
.Y(n_6011)
);

OAI22xp5_ASAP7_75t_L g6012 ( 
.A1(n_5182),
.A2(n_4633),
.B1(n_4565),
.B2(n_4342),
.Y(n_6012)
);

HB1xp67_ASAP7_75t_L g6013 ( 
.A(n_5680),
.Y(n_6013)
);

AOI22xp33_ASAP7_75t_L g6014 ( 
.A1(n_5212),
.A2(n_4612),
.B1(n_4588),
.B2(n_4874),
.Y(n_6014)
);

BUFx3_ASAP7_75t_L g6015 ( 
.A(n_5106),
.Y(n_6015)
);

OAI31xp33_ASAP7_75t_L g6016 ( 
.A1(n_5427),
.A2(n_4351),
.A3(n_4520),
.B(n_4250),
.Y(n_6016)
);

OAI21x1_ASAP7_75t_L g6017 ( 
.A1(n_5668),
.A2(n_4778),
.B(n_4961),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5751),
.B(n_5128),
.Y(n_6018)
);

AOI22xp5_ASAP7_75t_L g6019 ( 
.A1(n_5353),
.A2(n_4346),
.B1(n_4365),
.B2(n_4360),
.Y(n_6019)
);

AOI22xp33_ASAP7_75t_L g6020 ( 
.A1(n_5184),
.A2(n_4932),
.B1(n_4874),
.B2(n_4414),
.Y(n_6020)
);

NAND2xp5_ASAP7_75t_L g6021 ( 
.A(n_5365),
.B(n_4813),
.Y(n_6021)
);

INVx2_ASAP7_75t_SL g6022 ( 
.A(n_5408),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5664),
.Y(n_6023)
);

BUFx6f_ASAP7_75t_L g6024 ( 
.A(n_5094),
.Y(n_6024)
);

OAI22xp5_ASAP7_75t_L g6025 ( 
.A1(n_5175),
.A2(n_4360),
.B1(n_4365),
.B2(n_4346),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_L g6026 ( 
.A(n_5438),
.B(n_4814),
.Y(n_6026)
);

A2O1A1Ixp33_ASAP7_75t_L g6027 ( 
.A1(n_5560),
.A2(n_4587),
.B(n_4991),
.C(n_5049),
.Y(n_6027)
);

AOI21xp5_ASAP7_75t_L g6028 ( 
.A1(n_5598),
.A2(n_4946),
.B(n_4944),
.Y(n_6028)
);

O2A1O1Ixp5_ASAP7_75t_L g6029 ( 
.A1(n_5579),
.A2(n_5009),
.B(n_4996),
.C(n_4939),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5664),
.Y(n_6030)
);

AO32x2_ASAP7_75t_L g6031 ( 
.A1(n_5624),
.A2(n_4996),
.A3(n_4923),
.B1(n_4455),
.B2(n_4084),
.Y(n_6031)
);

INVxp67_ASAP7_75t_L g6032 ( 
.A(n_5154),
.Y(n_6032)
);

INVx6_ASAP7_75t_SL g6033 ( 
.A(n_5160),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5664),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5438),
.B(n_4821),
.Y(n_6035)
);

HB1xp67_ASAP7_75t_L g6036 ( 
.A(n_5680),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5664),
.Y(n_6037)
);

NAND2xp5_ASAP7_75t_L g6038 ( 
.A(n_5441),
.B(n_5454),
.Y(n_6038)
);

AOI21xp5_ASAP7_75t_L g6039 ( 
.A1(n_5598),
.A2(n_4958),
.B(n_4944),
.Y(n_6039)
);

AOI22xp5_ASAP7_75t_L g6040 ( 
.A1(n_5145),
.A2(n_4382),
.B1(n_4388),
.B2(n_4386),
.Y(n_6040)
);

AO21x1_ASAP7_75t_L g6041 ( 
.A1(n_5551),
.A2(n_4823),
.B(n_4821),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5666),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5666),
.Y(n_6043)
);

NAND2xp5_ASAP7_75t_L g6044 ( 
.A(n_5441),
.B(n_4823),
.Y(n_6044)
);

NAND2xp5_ASAP7_75t_L g6045 ( 
.A(n_5454),
.B(n_4852),
.Y(n_6045)
);

OAI22xp5_ASAP7_75t_L g6046 ( 
.A1(n_5167),
.A2(n_4382),
.B1(n_4388),
.B2(n_4386),
.Y(n_6046)
);

INVx5_ASAP7_75t_L g6047 ( 
.A(n_5408),
.Y(n_6047)
);

NOR2xp33_ASAP7_75t_L g6048 ( 
.A(n_5350),
.B(n_5006),
.Y(n_6048)
);

INVx1_ASAP7_75t_SL g6049 ( 
.A(n_5399),
.Y(n_6049)
);

A2O1A1Ixp33_ASAP7_75t_L g6050 ( 
.A1(n_5560),
.A2(n_5049),
.B(n_5075),
.C(n_5057),
.Y(n_6050)
);

AOI21xp5_ASAP7_75t_L g6051 ( 
.A1(n_5628),
.A2(n_4967),
.B(n_4958),
.Y(n_6051)
);

BUFx3_ASAP7_75t_L g6052 ( 
.A(n_5146),
.Y(n_6052)
);

AOI21xp5_ASAP7_75t_L g6053 ( 
.A1(n_5628),
.A2(n_4973),
.B(n_4967),
.Y(n_6053)
);

NAND2x1_ASAP7_75t_L g6054 ( 
.A(n_5726),
.B(n_5478),
.Y(n_6054)
);

AOI21xp5_ASAP7_75t_L g6055 ( 
.A1(n_5758),
.A2(n_4988),
.B(n_4973),
.Y(n_6055)
);

AO22x1_ASAP7_75t_L g6056 ( 
.A1(n_5385),
.A2(n_5551),
.B1(n_5267),
.B2(n_5319),
.Y(n_6056)
);

O2A1O1Ixp5_ASAP7_75t_L g6057 ( 
.A1(n_5579),
.A2(n_4955),
.B(n_4969),
.C(n_4937),
.Y(n_6057)
);

O2A1O1Ixp33_ASAP7_75t_L g6058 ( 
.A1(n_5237),
.A2(n_5034),
.B(n_5048),
.C(n_4520),
.Y(n_6058)
);

BUFx2_ASAP7_75t_L g6059 ( 
.A(n_5113),
.Y(n_6059)
);

INVx2_ASAP7_75t_SL g6060 ( 
.A(n_5408),
.Y(n_6060)
);

A2O1A1Ixp33_ASAP7_75t_L g6061 ( 
.A1(n_5476),
.A2(n_5057),
.B(n_5075),
.C(n_5014),
.Y(n_6061)
);

BUFx6f_ASAP7_75t_L g6062 ( 
.A(n_5094),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5495),
.B(n_4852),
.Y(n_6063)
);

BUFx3_ASAP7_75t_L g6064 ( 
.A(n_5146),
.Y(n_6064)
);

AOI21xp5_ASAP7_75t_L g6065 ( 
.A1(n_5758),
.A2(n_4989),
.B(n_4988),
.Y(n_6065)
);

AND2x4_ASAP7_75t_SL g6066 ( 
.A(n_5216),
.B(n_4737),
.Y(n_6066)
);

BUFx3_ASAP7_75t_L g6067 ( 
.A(n_5146),
.Y(n_6067)
);

A2O1A1Ixp33_ASAP7_75t_SL g6068 ( 
.A1(n_5521),
.A2(n_5390),
.B(n_5303),
.C(n_5334),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5666),
.Y(n_6069)
);

O2A1O1Ixp5_ASAP7_75t_L g6070 ( 
.A1(n_5257),
.A2(n_5061),
.B(n_5021),
.C(n_5068),
.Y(n_6070)
);

BUFx2_ASAP7_75t_L g6071 ( 
.A(n_5113),
.Y(n_6071)
);

INVx6_ASAP7_75t_L g6072 ( 
.A(n_5279),
.Y(n_6072)
);

OR2x2_ASAP7_75t_L g6073 ( 
.A(n_5717),
.B(n_4331),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5666),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_5495),
.B(n_4864),
.Y(n_6075)
);

A2O1A1Ixp33_ASAP7_75t_L g6076 ( 
.A1(n_5606),
.A2(n_5075),
.B(n_4992),
.C(n_4999),
.Y(n_6076)
);

O2A1O1Ixp5_ASAP7_75t_L g6077 ( 
.A1(n_5257),
.A2(n_5021),
.B(n_5077),
.C(n_5068),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5491),
.B(n_5497),
.Y(n_6078)
);

BUFx4f_ASAP7_75t_SL g6079 ( 
.A(n_5294),
.Y(n_6079)
);

OAI21xp5_ASAP7_75t_L g6080 ( 
.A1(n_5368),
.A2(n_4600),
.B(n_4492),
.Y(n_6080)
);

INVx3_ASAP7_75t_L g6081 ( 
.A(n_5197),
.Y(n_6081)
);

AOI21xp5_ASAP7_75t_L g6082 ( 
.A1(n_5356),
.A2(n_4992),
.B(n_4989),
.Y(n_6082)
);

NOR2xp33_ASAP7_75t_L g6083 ( 
.A(n_5350),
.B(n_4980),
.Y(n_6083)
);

AND2x6_ASAP7_75t_L g6084 ( 
.A(n_5151),
.B(n_5045),
.Y(n_6084)
);

INVx2_ASAP7_75t_SL g6085 ( 
.A(n_5408),
.Y(n_6085)
);

INVx1_ASAP7_75t_SL g6086 ( 
.A(n_5399),
.Y(n_6086)
);

BUFx2_ASAP7_75t_L g6087 ( 
.A(n_5113),
.Y(n_6087)
);

AOI22xp5_ASAP7_75t_L g6088 ( 
.A1(n_5145),
.A2(n_4440),
.B1(n_4449),
.B2(n_4402),
.Y(n_6088)
);

NOR3xp33_ASAP7_75t_L g6089 ( 
.A(n_5234),
.B(n_5048),
.C(n_5077),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5685),
.Y(n_6090)
);

AOI21xp5_ASAP7_75t_L g6091 ( 
.A1(n_5396),
.A2(n_4999),
.B(n_5078),
.Y(n_6091)
);

INVx2_ASAP7_75t_SL g6092 ( 
.A(n_5408),
.Y(n_6092)
);

O2A1O1Ixp5_ASAP7_75t_SL g6093 ( 
.A1(n_5314),
.A2(n_5036),
.B(n_4905),
.C(n_4917),
.Y(n_6093)
);

CKINVDCx5p33_ASAP7_75t_R g6094 ( 
.A(n_5190),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5685),
.Y(n_6095)
);

AOI22xp33_ASAP7_75t_L g6096 ( 
.A1(n_5385),
.A2(n_4932),
.B1(n_4414),
.B2(n_4563),
.Y(n_6096)
);

INVx8_ASAP7_75t_L g6097 ( 
.A(n_5170),
.Y(n_6097)
);

BUFx3_ASAP7_75t_L g6098 ( 
.A(n_5146),
.Y(n_6098)
);

AOI22xp5_ASAP7_75t_L g6099 ( 
.A1(n_5368),
.A2(n_4440),
.B1(n_4449),
.B2(n_4402),
.Y(n_6099)
);

AND2x4_ASAP7_75t_L g6100 ( 
.A(n_5616),
.B(n_5639),
.Y(n_6100)
);

BUFx12f_ASAP7_75t_L g6101 ( 
.A(n_5168),
.Y(n_6101)
);

BUFx3_ASAP7_75t_L g6102 ( 
.A(n_5136),
.Y(n_6102)
);

AOI21xp5_ASAP7_75t_L g6103 ( 
.A1(n_5396),
.A2(n_5079),
.B(n_5078),
.Y(n_6103)
);

CKINVDCx5p33_ASAP7_75t_R g6104 ( 
.A(n_5190),
.Y(n_6104)
);

OAI22xp5_ASAP7_75t_L g6105 ( 
.A1(n_5263),
.A2(n_4453),
.B1(n_4457),
.B2(n_4454),
.Y(n_6105)
);

BUFx4_ASAP7_75t_SL g6106 ( 
.A(n_5294),
.Y(n_6106)
);

AOI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_5412),
.A2(n_5084),
.B(n_5079),
.Y(n_6107)
);

A2O1A1Ixp33_ASAP7_75t_SL g6108 ( 
.A1(n_5303),
.A2(n_4903),
.B(n_4892),
.C(n_5012),
.Y(n_6108)
);

AOI221xp5_ASAP7_75t_L g6109 ( 
.A1(n_5428),
.A2(n_4819),
.B1(n_4663),
.B2(n_4471),
.C(n_4462),
.Y(n_6109)
);

AOI21xp5_ASAP7_75t_L g6110 ( 
.A1(n_5412),
.A2(n_5084),
.B(n_4938),
.Y(n_6110)
);

CKINVDCx6p67_ASAP7_75t_R g6111 ( 
.A(n_5505),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_5685),
.Y(n_6112)
);

NOR2xp33_ASAP7_75t_SL g6113 ( 
.A(n_5252),
.B(n_4827),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5685),
.Y(n_6114)
);

AOI22xp33_ASAP7_75t_L g6115 ( 
.A1(n_5355),
.A2(n_5252),
.B1(n_5263),
.B2(n_5376),
.Y(n_6115)
);

OAI22xp5_ASAP7_75t_L g6116 ( 
.A1(n_5335),
.A2(n_4466),
.B1(n_4453),
.B2(n_4454),
.Y(n_6116)
);

AOI22xp33_ASAP7_75t_L g6117 ( 
.A1(n_5355),
.A2(n_4551),
.B1(n_4563),
.B2(n_4599),
.Y(n_6117)
);

NAND2xp5_ASAP7_75t_SL g6118 ( 
.A(n_5486),
.B(n_5554),
.Y(n_6118)
);

INVx1_ASAP7_75t_SL g6119 ( 
.A(n_5399),
.Y(n_6119)
);

BUFx2_ASAP7_75t_L g6120 ( 
.A(n_5113),
.Y(n_6120)
);

O2A1O1Ixp5_ASAP7_75t_L g6121 ( 
.A1(n_5257),
.A2(n_5017),
.B(n_5031),
.C(n_5026),
.Y(n_6121)
);

NAND2xp5_ASAP7_75t_L g6122 ( 
.A(n_5513),
.B(n_4492),
.Y(n_6122)
);

O2A1O1Ixp5_ASAP7_75t_L g6123 ( 
.A1(n_5314),
.A2(n_5017),
.B(n_5031),
.C(n_5026),
.Y(n_6123)
);

AOI21xp5_ASAP7_75t_L g6124 ( 
.A1(n_5446),
.A2(n_4938),
.B(n_5025),
.Y(n_6124)
);

OAI21x1_ASAP7_75t_L g6125 ( 
.A1(n_5668),
.A2(n_4600),
.B(n_5054),
.Y(n_6125)
);

AOI21xp5_ASAP7_75t_L g6126 ( 
.A1(n_5446),
.A2(n_5025),
.B(n_5085),
.Y(n_6126)
);

BUFx2_ASAP7_75t_L g6127 ( 
.A(n_5113),
.Y(n_6127)
);

AOI22xp5_ASAP7_75t_L g6128 ( 
.A1(n_5368),
.A2(n_4570),
.B1(n_4462),
.B2(n_4466),
.Y(n_6128)
);

AOI21xp5_ASAP7_75t_L g6129 ( 
.A1(n_5464),
.A2(n_5088),
.B(n_5085),
.Y(n_6129)
);

INVx2_ASAP7_75t_SL g6130 ( 
.A(n_5408),
.Y(n_6130)
);

AOI22xp33_ASAP7_75t_L g6131 ( 
.A1(n_5376),
.A2(n_4599),
.B1(n_4613),
.B2(n_4781),
.Y(n_6131)
);

OR2x6_ASAP7_75t_L g6132 ( 
.A(n_5160),
.B(n_5205),
.Y(n_6132)
);

AOI22xp33_ASAP7_75t_L g6133 ( 
.A1(n_5428),
.A2(n_4609),
.B1(n_4613),
.B2(n_4781),
.Y(n_6133)
);

CKINVDCx20_ASAP7_75t_R g6134 ( 
.A(n_5261),
.Y(n_6134)
);

AOI22xp33_ASAP7_75t_L g6135 ( 
.A1(n_5428),
.A2(n_4609),
.B1(n_4457),
.B2(n_4570),
.Y(n_6135)
);

NAND3xp33_ASAP7_75t_L g6136 ( 
.A(n_5401),
.B(n_5002),
.C(n_5018),
.Y(n_6136)
);

HB1xp67_ASAP7_75t_L g6137 ( 
.A(n_5713),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5702),
.Y(n_6138)
);

AOI21xp5_ASAP7_75t_L g6139 ( 
.A1(n_5464),
.A2(n_5088),
.B(n_5054),
.Y(n_6139)
);

CKINVDCx11_ASAP7_75t_R g6140 ( 
.A(n_5261),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5702),
.Y(n_6141)
);

CKINVDCx20_ASAP7_75t_R g6142 ( 
.A(n_5270),
.Y(n_6142)
);

AND2x4_ASAP7_75t_SL g6143 ( 
.A(n_5216),
.B(n_5289),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5702),
.Y(n_6144)
);

CKINVDCx20_ASAP7_75t_R g6145 ( 
.A(n_5270),
.Y(n_6145)
);

INVxp67_ASAP7_75t_L g6146 ( 
.A(n_5154),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_5770),
.B(n_4073),
.Y(n_6147)
);

NOR2xp33_ASAP7_75t_L g6148 ( 
.A(n_5267),
.B(n_4993),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5702),
.Y(n_6149)
);

INVx1_ASAP7_75t_L g6150 ( 
.A(n_5705),
.Y(n_6150)
);

NAND2xp5_ASAP7_75t_L g6151 ( 
.A(n_5770),
.B(n_4074),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5705),
.Y(n_6152)
);

AOI22xp5_ASAP7_75t_L g6153 ( 
.A1(n_5427),
.A2(n_4554),
.B1(n_4486),
.B2(n_4506),
.Y(n_6153)
);

OR2x2_ASAP7_75t_L g6154 ( 
.A(n_5622),
.B(n_4074),
.Y(n_6154)
);

BUFx6f_ASAP7_75t_L g6155 ( 
.A(n_5144),
.Y(n_6155)
);

NOR2xp33_ASAP7_75t_SL g6156 ( 
.A(n_5380),
.B(n_4398),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5705),
.Y(n_6157)
);

INVx2_ASAP7_75t_SL g6158 ( 
.A(n_5611),
.Y(n_6158)
);

NAND2xp5_ASAP7_75t_SL g6159 ( 
.A(n_5486),
.B(n_4737),
.Y(n_6159)
);

AOI21xp5_ASAP7_75t_L g6160 ( 
.A1(n_5576),
.A2(n_5502),
.B(n_5509),
.Y(n_6160)
);

AND2x6_ASAP7_75t_L g6161 ( 
.A(n_5151),
.B(n_4398),
.Y(n_6161)
);

NAND2xp5_ASAP7_75t_SL g6162 ( 
.A(n_5486),
.B(n_4737),
.Y(n_6162)
);

INVxp67_ASAP7_75t_L g6163 ( 
.A(n_5364),
.Y(n_6163)
);

AOI21xp5_ASAP7_75t_L g6164 ( 
.A1(n_5576),
.A2(n_5039),
.B(n_5055),
.Y(n_6164)
);

INVx1_ASAP7_75t_L g6165 ( 
.A(n_5705),
.Y(n_6165)
);

AND2x4_ASAP7_75t_L g6166 ( 
.A(n_5616),
.B(n_5639),
.Y(n_6166)
);

NAND2xp5_ASAP7_75t_L g6167 ( 
.A(n_5770),
.B(n_4083),
.Y(n_6167)
);

AOI21xp5_ASAP7_75t_L g6168 ( 
.A1(n_5502),
.A2(n_5039),
.B(n_5080),
.Y(n_6168)
);

BUFx3_ASAP7_75t_L g6169 ( 
.A(n_5149),
.Y(n_6169)
);

CKINVDCx6p67_ASAP7_75t_R g6170 ( 
.A(n_5149),
.Y(n_6170)
);

INVx2_ASAP7_75t_SL g6171 ( 
.A(n_5611),
.Y(n_6171)
);

AOI21xp33_ASAP7_75t_L g6172 ( 
.A1(n_5334),
.A2(n_4663),
.B(n_4083),
.Y(n_6172)
);

AOI21xp5_ASAP7_75t_L g6173 ( 
.A1(n_5502),
.A2(n_5082),
.B(n_5046),
.Y(n_6173)
);

NAND2xp5_ASAP7_75t_SL g6174 ( 
.A(n_5554),
.B(n_4870),
.Y(n_6174)
);

OAI22xp5_ASAP7_75t_L g6175 ( 
.A1(n_5244),
.A2(n_4592),
.B1(n_4506),
.B2(n_4544),
.Y(n_6175)
);

OR2x2_ASAP7_75t_L g6176 ( 
.A(n_5622),
.B(n_4085),
.Y(n_6176)
);

INVx1_ASAP7_75t_SL g6177 ( 
.A(n_5652),
.Y(n_6177)
);

A2O1A1Ixp33_ASAP7_75t_L g6178 ( 
.A1(n_5606),
.A2(n_4892),
.B(n_4461),
.C(n_4557),
.Y(n_6178)
);

NAND2xp5_ASAP7_75t_L g6179 ( 
.A(n_5630),
.B(n_4093),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_5728),
.Y(n_6180)
);

INVx3_ASAP7_75t_L g6181 ( 
.A(n_5220),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5728),
.Y(n_6182)
);

OAI22xp5_ASAP7_75t_L g6183 ( 
.A1(n_5244),
.A2(n_4592),
.B1(n_4544),
.B2(n_4548),
.Y(n_6183)
);

NAND2xp5_ASAP7_75t_L g6184 ( 
.A(n_5630),
.B(n_4093),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_5728),
.Y(n_6185)
);

NAND2xp5_ASAP7_75t_L g6186 ( 
.A(n_5631),
.B(n_4099),
.Y(n_6186)
);

BUFx2_ASAP7_75t_L g6187 ( 
.A(n_5113),
.Y(n_6187)
);

OAI22xp5_ASAP7_75t_L g6188 ( 
.A1(n_5244),
.A2(n_4576),
.B1(n_4548),
.B2(n_4553),
.Y(n_6188)
);

NAND2xp5_ASAP7_75t_L g6189 ( 
.A(n_5631),
.B(n_4099),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5728),
.Y(n_6190)
);

AOI22xp5_ASAP7_75t_L g6191 ( 
.A1(n_5319),
.A2(n_4554),
.B1(n_4576),
.B2(n_4562),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_5732),
.Y(n_6192)
);

HB1xp67_ASAP7_75t_L g6193 ( 
.A(n_5713),
.Y(n_6193)
);

AOI21xp5_ASAP7_75t_L g6194 ( 
.A1(n_5509),
.A2(n_5046),
.B(n_5058),
.Y(n_6194)
);

INVx2_ASAP7_75t_SL g6195 ( 
.A(n_5611),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_L g6196 ( 
.A(n_5699),
.B(n_4135),
.Y(n_6196)
);

BUFx12f_ASAP7_75t_L g6197 ( 
.A(n_5199),
.Y(n_6197)
);

A2O1A1Ixp33_ASAP7_75t_L g6198 ( 
.A1(n_5750),
.A2(n_4461),
.B(n_4557),
.C(n_4706),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_5732),
.Y(n_6199)
);

BUFx2_ASAP7_75t_L g6200 ( 
.A(n_5160),
.Y(n_6200)
);

NAND2xp5_ASAP7_75t_L g6201 ( 
.A(n_5699),
.B(n_4135),
.Y(n_6201)
);

AOI21xp5_ASAP7_75t_L g6202 ( 
.A1(n_5509),
.A2(n_5058),
.B(n_4866),
.Y(n_6202)
);

BUFx6f_ASAP7_75t_L g6203 ( 
.A(n_5144),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_L g6204 ( 
.A(n_5507),
.B(n_4143),
.Y(n_6204)
);

AOI21x1_ASAP7_75t_L g6205 ( 
.A1(n_5392),
.A2(n_4663),
.B(n_5002),
.Y(n_6205)
);

INVx3_ASAP7_75t_L g6206 ( 
.A(n_5220),
.Y(n_6206)
);

AOI22xp5_ASAP7_75t_L g6207 ( 
.A1(n_5271),
.A2(n_4572),
.B1(n_4486),
.B2(n_4553),
.Y(n_6207)
);

BUFx12f_ASAP7_75t_L g6208 ( 
.A(n_5199),
.Y(n_6208)
);

AOI22xp33_ASAP7_75t_L g6209 ( 
.A1(n_5421),
.A2(n_4562),
.B1(n_4572),
.B2(n_4557),
.Y(n_6209)
);

A2O1A1Ixp33_ASAP7_75t_L g6210 ( 
.A1(n_5750),
.A2(n_4461),
.B(n_4706),
.C(n_4896),
.Y(n_6210)
);

INVx1_ASAP7_75t_SL g6211 ( 
.A(n_5652),
.Y(n_6211)
);

NOR2xp67_ASAP7_75t_SL g6212 ( 
.A(n_5584),
.B(n_4918),
.Y(n_6212)
);

OAI22xp5_ASAP7_75t_L g6213 ( 
.A1(n_5271),
.A2(n_4520),
.B1(n_4351),
.B2(n_4224),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_5732),
.Y(n_6214)
);

NAND2xp5_ASAP7_75t_SL g6215 ( 
.A(n_5463),
.B(n_4870),
.Y(n_6215)
);

NAND2xp5_ASAP7_75t_SL g6216 ( 
.A(n_5463),
.B(n_4870),
.Y(n_6216)
);

INVxp67_ASAP7_75t_L g6217 ( 
.A(n_5466),
.Y(n_6217)
);

AOI21xp5_ASAP7_75t_L g6218 ( 
.A1(n_5510),
.A2(n_4902),
.B(n_4862),
.Y(n_6218)
);

AOI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_5510),
.A2(n_4902),
.B(n_4866),
.Y(n_6219)
);

HB1xp67_ASAP7_75t_L g6220 ( 
.A(n_5713),
.Y(n_6220)
);

BUFx2_ASAP7_75t_L g6221 ( 
.A(n_5160),
.Y(n_6221)
);

INVx3_ASAP7_75t_L g6222 ( 
.A(n_5228),
.Y(n_6222)
);

NAND3xp33_ASAP7_75t_L g6223 ( 
.A(n_5401),
.B(n_4880),
.C(n_4922),
.Y(n_6223)
);

AOI21xp5_ASAP7_75t_L g6224 ( 
.A1(n_5510),
.A2(n_4901),
.B(n_4922),
.Y(n_6224)
);

AOI21xp5_ASAP7_75t_L g6225 ( 
.A1(n_5515),
.A2(n_5526),
.B(n_5522),
.Y(n_6225)
);

INVx2_ASAP7_75t_SL g6226 ( 
.A(n_5611),
.Y(n_6226)
);

INVx2_ASAP7_75t_SL g6227 ( 
.A(n_5611),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_5507),
.B(n_4143),
.Y(n_6228)
);

OAI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_5271),
.A2(n_4351),
.B1(n_4520),
.B2(n_4239),
.Y(n_6229)
);

INVx4_ASAP7_75t_L g6230 ( 
.A(n_5149),
.Y(n_6230)
);

INVx4_ASAP7_75t_L g6231 ( 
.A(n_5149),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_5732),
.Y(n_6232)
);

CKINVDCx5p33_ASAP7_75t_R g6233 ( 
.A(n_5612),
.Y(n_6233)
);

CKINVDCx11_ASAP7_75t_R g6234 ( 
.A(n_5562),
.Y(n_6234)
);

AOI21xp5_ASAP7_75t_L g6235 ( 
.A1(n_5515),
.A2(n_4883),
.B(n_4901),
.Y(n_6235)
);

INVx2_ASAP7_75t_SL g6236 ( 
.A(n_5611),
.Y(n_6236)
);

NOR2xp33_ASAP7_75t_L g6237 ( 
.A(n_5236),
.B(n_4993),
.Y(n_6237)
);

NOR2xp33_ASAP7_75t_L g6238 ( 
.A(n_5236),
.B(n_5005),
.Y(n_6238)
);

AO21x2_ASAP7_75t_L g6239 ( 
.A1(n_5523),
.A2(n_5083),
.B(n_5064),
.Y(n_6239)
);

NAND2xp33_ASAP7_75t_L g6240 ( 
.A(n_5278),
.B(n_4657),
.Y(n_6240)
);

NAND2xp5_ASAP7_75t_L g6241 ( 
.A(n_5507),
.B(n_4300),
.Y(n_6241)
);

O2A1O1Ixp33_ASAP7_75t_L g6242 ( 
.A1(n_5432),
.A2(n_4883),
.B(n_4882),
.C(n_4880),
.Y(n_6242)
);

INVx3_ASAP7_75t_SL g6243 ( 
.A(n_5731),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_5733),
.Y(n_6244)
);

BUFx3_ASAP7_75t_L g6245 ( 
.A(n_5217),
.Y(n_6245)
);

AOI21xp5_ASAP7_75t_L g6246 ( 
.A1(n_5515),
.A2(n_4879),
.B(n_4882),
.Y(n_6246)
);

BUFx3_ASAP7_75t_L g6247 ( 
.A(n_5217),
.Y(n_6247)
);

OAI22xp5_ASAP7_75t_L g6248 ( 
.A1(n_5346),
.A2(n_4214),
.B1(n_4224),
.B2(n_4239),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_5733),
.Y(n_6249)
);

NOR2x1_ASAP7_75t_SL g6250 ( 
.A(n_5746),
.B(n_4870),
.Y(n_6250)
);

O2A1O1Ixp5_ASAP7_75t_L g6251 ( 
.A1(n_5314),
.A2(n_4925),
.B(n_4776),
.C(n_4830),
.Y(n_6251)
);

NAND2xp33_ASAP7_75t_L g6252 ( 
.A(n_5278),
.B(n_4787),
.Y(n_6252)
);

AOI21xp5_ASAP7_75t_L g6253 ( 
.A1(n_5522),
.A2(n_4879),
.B(n_4558),
.Y(n_6253)
);

AOI22xp33_ASAP7_75t_L g6254 ( 
.A1(n_5421),
.A2(n_5180),
.B1(n_5584),
.B2(n_5299),
.Y(n_6254)
);

AOI22xp33_ASAP7_75t_SL g6255 ( 
.A1(n_5397),
.A2(n_4776),
.B1(n_4925),
.B2(n_4830),
.Y(n_6255)
);

AOI22xp5_ASAP7_75t_L g6256 ( 
.A1(n_5260),
.A2(n_4376),
.B1(n_4981),
.B2(n_4964),
.Y(n_6256)
);

INVx5_ASAP7_75t_L g6257 ( 
.A(n_5611),
.Y(n_6257)
);

INVx5_ASAP7_75t_L g6258 ( 
.A(n_5611),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_5771),
.B(n_4320),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_SL g6260 ( 
.A(n_5463),
.B(n_5780),
.Y(n_6260)
);

NOR2xp33_ASAP7_75t_L g6261 ( 
.A(n_5236),
.B(n_5202),
.Y(n_6261)
);

CKINVDCx5p33_ASAP7_75t_R g6262 ( 
.A(n_5612),
.Y(n_6262)
);

BUFx12f_ASAP7_75t_L g6263 ( 
.A(n_5307),
.Y(n_6263)
);

INVx1_ASAP7_75t_SL g6264 ( 
.A(n_5652),
.Y(n_6264)
);

BUFx2_ASAP7_75t_L g6265 ( 
.A(n_5160),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5733),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_5771),
.B(n_4320),
.Y(n_6267)
);

NOR2xp67_ASAP7_75t_L g6268 ( 
.A(n_5239),
.B(n_5264),
.Y(n_6268)
);

O2A1O1Ixp5_ASAP7_75t_L g6269 ( 
.A1(n_5303),
.A2(n_4925),
.B(n_4646),
.C(n_4776),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5733),
.Y(n_6270)
);

BUFx6f_ASAP7_75t_L g6271 ( 
.A(n_5144),
.Y(n_6271)
);

AND2x2_ASAP7_75t_L g6272 ( 
.A(n_5282),
.B(n_5293),
.Y(n_6272)
);

AOI21xp5_ASAP7_75t_L g6273 ( 
.A1(n_5522),
.A2(n_4716),
.B(n_4923),
.Y(n_6273)
);

INVx3_ASAP7_75t_SL g6274 ( 
.A(n_5375),
.Y(n_6274)
);

BUFx12f_ASAP7_75t_L g6275 ( 
.A(n_5307),
.Y(n_6275)
);

NAND3xp33_ASAP7_75t_L g6276 ( 
.A(n_5299),
.B(n_5051),
.C(n_5062),
.Y(n_6276)
);

INVx2_ASAP7_75t_SL g6277 ( 
.A(n_5639),
.Y(n_6277)
);

AOI22xp33_ASAP7_75t_L g6278 ( 
.A1(n_5421),
.A2(n_4376),
.B1(n_4759),
.B2(n_4700),
.Y(n_6278)
);

OAI22xp5_ASAP7_75t_L g6279 ( 
.A1(n_5346),
.A2(n_4338),
.B1(n_4359),
.B2(n_4368),
.Y(n_6279)
);

BUFx6f_ASAP7_75t_L g6280 ( 
.A(n_5144),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_5738),
.Y(n_6281)
);

BUFx6f_ASAP7_75t_L g6282 ( 
.A(n_5144),
.Y(n_6282)
);

OAI21xp5_ASAP7_75t_L g6283 ( 
.A1(n_5574),
.A2(n_5030),
.B(n_5012),
.Y(n_6283)
);

AOI22xp5_ASAP7_75t_L g6284 ( 
.A1(n_5260),
.A2(n_4376),
.B1(n_4964),
.B2(n_4941),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_5738),
.Y(n_6285)
);

INVx2_ASAP7_75t_SL g6286 ( 
.A(n_5639),
.Y(n_6286)
);

O2A1O1Ixp33_ASAP7_75t_L g6287 ( 
.A1(n_5432),
.A2(n_5005),
.B(n_5051),
.C(n_5062),
.Y(n_6287)
);

BUFx3_ASAP7_75t_L g6288 ( 
.A(n_5217),
.Y(n_6288)
);

BUFx3_ASAP7_75t_L g6289 ( 
.A(n_5217),
.Y(n_6289)
);

NAND2x1p5_ASAP7_75t_L g6290 ( 
.A(n_5141),
.B(n_4646),
.Y(n_6290)
);

NOR2xp33_ASAP7_75t_R g6291 ( 
.A(n_5473),
.B(n_4801),
.Y(n_6291)
);

BUFx3_ASAP7_75t_L g6292 ( 
.A(n_5227),
.Y(n_6292)
);

AOI222xp33_ASAP7_75t_L g6293 ( 
.A1(n_5367),
.A2(n_4397),
.B1(n_4404),
.B2(n_4419),
.C1(n_4431),
.C2(n_4439),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5738),
.Y(n_6294)
);

OAI21xp5_ASAP7_75t_L g6295 ( 
.A1(n_5574),
.A2(n_5030),
.B(n_4761),
.Y(n_6295)
);

A2O1A1Ixp33_ASAP7_75t_SL g6296 ( 
.A1(n_5671),
.A2(n_4986),
.B(n_5070),
.C(n_4830),
.Y(n_6296)
);

NOR2xp33_ASAP7_75t_R g6297 ( 
.A(n_5473),
.B(n_4801),
.Y(n_6297)
);

AOI22xp5_ASAP7_75t_L g6298 ( 
.A1(n_5260),
.A2(n_4941),
.B1(n_4830),
.B2(n_4925),
.Y(n_6298)
);

AOI21xp5_ASAP7_75t_L g6299 ( 
.A1(n_5526),
.A2(n_5087),
.B(n_5083),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5738),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5745),
.Y(n_6301)
);

NOR2xp33_ASAP7_75t_L g6302 ( 
.A(n_5202),
.B(n_4700),
.Y(n_6302)
);

BUFx6f_ASAP7_75t_L g6303 ( 
.A(n_5144),
.Y(n_6303)
);

AOI21xp5_ASAP7_75t_L g6304 ( 
.A1(n_5526),
.A2(n_5087),
.B(n_4804),
.Y(n_6304)
);

AOI22xp5_ASAP7_75t_L g6305 ( 
.A1(n_5397),
.A2(n_4533),
.B1(n_4512),
.B2(n_5010),
.Y(n_6305)
);

OAI22xp5_ASAP7_75t_L g6306 ( 
.A1(n_5114),
.A2(n_4397),
.B1(n_4404),
.B2(n_4419),
.Y(n_6306)
);

AOI21xp5_ASAP7_75t_L g6307 ( 
.A1(n_5542),
.A2(n_4783),
.B(n_4815),
.Y(n_6307)
);

A2O1A1Ixp33_ASAP7_75t_L g6308 ( 
.A1(n_5444),
.A2(n_4838),
.B(n_4896),
.C(n_4904),
.Y(n_6308)
);

AOI21xp5_ASAP7_75t_L g6309 ( 
.A1(n_5542),
.A2(n_5238),
.B(n_5387),
.Y(n_6309)
);

A2O1A1Ixp33_ASAP7_75t_L g6310 ( 
.A1(n_5444),
.A2(n_4838),
.B(n_4896),
.C(n_4904),
.Y(n_6310)
);

BUFx6f_ASAP7_75t_L g6311 ( 
.A(n_5144),
.Y(n_6311)
);

NAND2x1p5_ASAP7_75t_L g6312 ( 
.A(n_5141),
.B(n_4986),
.Y(n_6312)
);

AOI22xp5_ASAP7_75t_L g6313 ( 
.A1(n_5397),
.A2(n_5010),
.B1(n_4591),
.B2(n_4700),
.Y(n_6313)
);

AOI21xp5_ASAP7_75t_L g6314 ( 
.A1(n_5542),
.A2(n_4820),
.B(n_4822),
.Y(n_6314)
);

INVx2_ASAP7_75t_SL g6315 ( 
.A(n_5691),
.Y(n_6315)
);

AOI21xp5_ASAP7_75t_L g6316 ( 
.A1(n_5238),
.A2(n_4820),
.B(n_4822),
.Y(n_6316)
);

AO21x1_ASAP7_75t_L g6317 ( 
.A1(n_5466),
.A2(n_4445),
.B(n_4447),
.Y(n_6317)
);

CKINVDCx5p33_ASAP7_75t_R g6318 ( 
.A(n_5568),
.Y(n_6318)
);

INVxp67_ASAP7_75t_L g6319 ( 
.A(n_5377),
.Y(n_6319)
);

BUFx3_ASAP7_75t_L g6320 ( 
.A(n_5227),
.Y(n_6320)
);

INVx5_ASAP7_75t_L g6321 ( 
.A(n_5144),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5745),
.Y(n_6322)
);

BUFx3_ASAP7_75t_L g6323 ( 
.A(n_5227),
.Y(n_6323)
);

INVx5_ASAP7_75t_L g6324 ( 
.A(n_5144),
.Y(n_6324)
);

NAND2xp5_ASAP7_75t_L g6325 ( 
.A(n_5214),
.B(n_5240),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_5745),
.Y(n_6326)
);

AOI21xp5_ASAP7_75t_L g6327 ( 
.A1(n_5238),
.A2(n_4790),
.B(n_4815),
.Y(n_6327)
);

BUFx6f_ASAP7_75t_L g6328 ( 
.A(n_5144),
.Y(n_6328)
);

AND2x2_ASAP7_75t_L g6329 ( 
.A(n_5320),
.B(n_5064),
.Y(n_6329)
);

NOR2xp33_ASAP7_75t_SL g6330 ( 
.A(n_5380),
.B(n_4801),
.Y(n_6330)
);

INVx1_ASAP7_75t_SL g6331 ( 
.A(n_5661),
.Y(n_6331)
);

OAI22xp5_ASAP7_75t_L g6332 ( 
.A1(n_5114),
.A2(n_4510),
.B1(n_4522),
.B2(n_4547),
.Y(n_6332)
);

INVx1_ASAP7_75t_SL g6333 ( 
.A(n_5661),
.Y(n_6333)
);

HB1xp67_ASAP7_75t_L g6334 ( 
.A(n_5138),
.Y(n_6334)
);

INVx3_ASAP7_75t_SL g6335 ( 
.A(n_5375),
.Y(n_6335)
);

AND2x2_ASAP7_75t_L g6336 ( 
.A(n_5320),
.B(n_5065),
.Y(n_6336)
);

INVx1_ASAP7_75t_SL g6337 ( 
.A(n_5661),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_5290),
.B(n_5233),
.Y(n_6338)
);

INVx2_ASAP7_75t_SL g6339 ( 
.A(n_5691),
.Y(n_6339)
);

AND2x2_ASAP7_75t_L g6340 ( 
.A(n_5322),
.B(n_5065),
.Y(n_6340)
);

CKINVDCx8_ASAP7_75t_R g6341 ( 
.A(n_5398),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_L g6342 ( 
.A(n_5290),
.B(n_5233),
.Y(n_6342)
);

AOI22xp5_ASAP7_75t_L g6343 ( 
.A1(n_5388),
.A2(n_4591),
.B1(n_4759),
.B2(n_4589),
.Y(n_6343)
);

CKINVDCx5p33_ASAP7_75t_R g6344 ( 
.A(n_5568),
.Y(n_6344)
);

CKINVDCx20_ASAP7_75t_R g6345 ( 
.A(n_5562),
.Y(n_6345)
);

NOR2xp33_ASAP7_75t_R g6346 ( 
.A(n_5203),
.B(n_4907),
.Y(n_6346)
);

OR2x2_ASAP7_75t_L g6347 ( 
.A(n_5322),
.B(n_4915),
.Y(n_6347)
);

HB1xp67_ASAP7_75t_SL g6348 ( 
.A(n_5572),
.Y(n_6348)
);

NOR2xp33_ASAP7_75t_SL g6349 ( 
.A(n_5671),
.B(n_4907),
.Y(n_6349)
);

CKINVDCx5p33_ASAP7_75t_R g6350 ( 
.A(n_5592),
.Y(n_6350)
);

CKINVDCx20_ASAP7_75t_R g6351 ( 
.A(n_5498),
.Y(n_6351)
);

A2O1A1Ixp33_ASAP7_75t_L g6352 ( 
.A1(n_5439),
.A2(n_4907),
.B(n_4838),
.C(n_4904),
.Y(n_6352)
);

NAND2xp5_ASAP7_75t_L g6353 ( 
.A(n_5233),
.B(n_5139),
.Y(n_6353)
);

OAI22xp5_ASAP7_75t_L g6354 ( 
.A1(n_5117),
.A2(n_4759),
.B1(n_5027),
.B2(n_4758),
.Y(n_6354)
);

INVx2_ASAP7_75t_SL g6355 ( 
.A(n_5691),
.Y(n_6355)
);

CKINVDCx5p33_ASAP7_75t_R g6356 ( 
.A(n_5592),
.Y(n_6356)
);

AND2x2_ASAP7_75t_L g6357 ( 
.A(n_5340),
.B(n_4968),
.Y(n_6357)
);

CKINVDCx20_ASAP7_75t_R g6358 ( 
.A(n_5498),
.Y(n_6358)
);

OR2x2_ASAP7_75t_L g6359 ( 
.A(n_5340),
.B(n_4976),
.Y(n_6359)
);

INVx6_ASAP7_75t_L g6360 ( 
.A(n_5279),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_5340),
.B(n_4976),
.Y(n_6361)
);

NOR2xp33_ASAP7_75t_L g6362 ( 
.A(n_5494),
.B(n_4976),
.Y(n_6362)
);

AOI21xp33_ASAP7_75t_L g6363 ( 
.A1(n_5442),
.A2(n_5076),
.B(n_5059),
.Y(n_6363)
);

INVxp67_ASAP7_75t_SL g6364 ( 
.A(n_5120),
.Y(n_6364)
);

AOI21xp5_ASAP7_75t_L g6365 ( 
.A1(n_5393),
.A2(n_4968),
.B(n_4970),
.Y(n_6365)
);

NOR2xp33_ASAP7_75t_L g6366 ( 
.A(n_5494),
.B(n_4968),
.Y(n_6366)
);

CKINVDCx5p33_ASAP7_75t_R g6367 ( 
.A(n_5276),
.Y(n_6367)
);

CKINVDCx5p33_ASAP7_75t_R g6368 ( 
.A(n_5276),
.Y(n_6368)
);

A2O1A1Ixp33_ASAP7_75t_L g6369 ( 
.A1(n_5439),
.A2(n_5070),
.B(n_4591),
.C(n_4936),
.Y(n_6369)
);

AND2x4_ASAP7_75t_L g6370 ( 
.A(n_5691),
.B(n_5762),
.Y(n_6370)
);

BUFx3_ASAP7_75t_L g6371 ( 
.A(n_5227),
.Y(n_6371)
);

AOI21xp5_ASAP7_75t_L g6372 ( 
.A1(n_5393),
.A2(n_5407),
.B(n_5405),
.Y(n_6372)
);

CKINVDCx5p33_ASAP7_75t_R g6373 ( 
.A(n_5269),
.Y(n_6373)
);

A2O1A1Ixp33_ASAP7_75t_SL g6374 ( 
.A1(n_5442),
.A2(n_4986),
.B(n_5019),
.C(n_5050),
.Y(n_6374)
);

NAND2xp5_ASAP7_75t_SL g6375 ( 
.A(n_5780),
.B(n_5008),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_L g6376 ( 
.A(n_5172),
.B(n_4975),
.Y(n_6376)
);

INVx5_ASAP7_75t_L g6377 ( 
.A(n_5567),
.Y(n_6377)
);

INVxp67_ASAP7_75t_L g6378 ( 
.A(n_5377),
.Y(n_6378)
);

NAND2xp5_ASAP7_75t_L g6379 ( 
.A(n_5127),
.B(n_4975),
.Y(n_6379)
);

AOI21xp5_ASAP7_75t_L g6380 ( 
.A1(n_5405),
.A2(n_4975),
.B(n_4870),
.Y(n_6380)
);

INVxp67_ASAP7_75t_SL g6381 ( 
.A(n_5120),
.Y(n_6381)
);

A2O1A1Ixp33_ASAP7_75t_L g6382 ( 
.A1(n_5512),
.A2(n_4936),
.B(n_4915),
.C(n_4976),
.Y(n_6382)
);

BUFx8_ASAP7_75t_L g6383 ( 
.A(n_5246),
.Y(n_6383)
);

OR2x6_ASAP7_75t_SL g6384 ( 
.A(n_5467),
.B(n_5485),
.Y(n_6384)
);

NAND2xp5_ASAP7_75t_L g6385 ( 
.A(n_5127),
.B(n_4975),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_5127),
.B(n_4970),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_5374),
.B(n_4970),
.Y(n_6387)
);

AOI21xp5_ASAP7_75t_L g6388 ( 
.A1(n_5405),
.A2(n_4976),
.B(n_4915),
.Y(n_6388)
);

NAND2x1p5_ASAP7_75t_L g6389 ( 
.A(n_5141),
.B(n_5008),
.Y(n_6389)
);

HB1xp67_ASAP7_75t_L g6390 ( 
.A(n_5138),
.Y(n_6390)
);

AO21x1_ASAP7_75t_L g6391 ( 
.A1(n_5467),
.A2(n_5020),
.B(n_5050),
.Y(n_6391)
);

INVx2_ASAP7_75t_SL g6392 ( 
.A(n_5762),
.Y(n_6392)
);

O2A1O1Ixp33_ASAP7_75t_L g6393 ( 
.A1(n_5563),
.A2(n_5076),
.B(n_5059),
.C(n_5053),
.Y(n_6393)
);

INVxp67_ASAP7_75t_SL g6394 ( 
.A(n_5490),
.Y(n_6394)
);

HB1xp67_ASAP7_75t_L g6395 ( 
.A(n_5159),
.Y(n_6395)
);

NAND2xp5_ASAP7_75t_L g6396 ( 
.A(n_5374),
.B(n_5754),
.Y(n_6396)
);

NOR2xp33_ASAP7_75t_SL g6397 ( 
.A(n_5345),
.B(n_4918),
.Y(n_6397)
);

NAND3xp33_ASAP7_75t_L g6398 ( 
.A(n_5461),
.B(n_5351),
.C(n_5325),
.Y(n_6398)
);

AOI22xp33_ASAP7_75t_L g6399 ( 
.A1(n_5180),
.A2(n_4970),
.B1(n_4915),
.B2(n_5008),
.Y(n_6399)
);

AOI21xp5_ASAP7_75t_L g6400 ( 
.A1(n_5407),
.A2(n_4915),
.B(n_5008),
.Y(n_6400)
);

BUFx12f_ASAP7_75t_L g6401 ( 
.A(n_5337),
.Y(n_6401)
);

AO21x1_ASAP7_75t_L g6402 ( 
.A1(n_5467),
.A2(n_5019),
.B(n_5028),
.Y(n_6402)
);

INVx4_ASAP7_75t_L g6403 ( 
.A(n_5246),
.Y(n_6403)
);

NAND2xp33_ASAP7_75t_L g6404 ( 
.A(n_5222),
.B(n_4787),
.Y(n_6404)
);

AOI22xp33_ASAP7_75t_SL g6405 ( 
.A1(n_5440),
.A2(n_5465),
.B1(n_5485),
.B2(n_5418),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_5754),
.B(n_4915),
.Y(n_6406)
);

INVx4_ASAP7_75t_L g6407 ( 
.A(n_5246),
.Y(n_6407)
);

AO21x1_ASAP7_75t_L g6408 ( 
.A1(n_5485),
.A2(n_5020),
.B(n_5035),
.Y(n_6408)
);

NOR2xp33_ASAP7_75t_L g6409 ( 
.A(n_5363),
.B(n_4976),
.Y(n_6409)
);

AOI21xp5_ASAP7_75t_L g6410 ( 
.A1(n_5407),
.A2(n_5027),
.B(n_5072),
.Y(n_6410)
);

CKINVDCx20_ASAP7_75t_R g6411 ( 
.A(n_5681),
.Y(n_6411)
);

OR2x2_ASAP7_75t_L g6412 ( 
.A(n_5391),
.B(n_4936),
.Y(n_6412)
);

AOI21xp5_ASAP7_75t_L g6413 ( 
.A1(n_5409),
.A2(n_5072),
.B(n_5023),
.Y(n_6413)
);

AOI221x1_ASAP7_75t_L g6414 ( 
.A1(n_5153),
.A2(n_5028),
.B1(n_5035),
.B2(n_5053),
.C(n_5043),
.Y(n_6414)
);

AOI21xp5_ASAP7_75t_L g6415 ( 
.A1(n_5409),
.A2(n_5072),
.B(n_5013),
.Y(n_6415)
);

NAND2xp5_ASAP7_75t_L g6416 ( 
.A(n_5763),
.B(n_5624),
.Y(n_6416)
);

NAND2xp5_ASAP7_75t_L g6417 ( 
.A(n_5763),
.B(n_5042),
.Y(n_6417)
);

AOI22xp33_ASAP7_75t_L g6418 ( 
.A1(n_5180),
.A2(n_4787),
.B1(n_5043),
.B2(n_5042),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_5624),
.B(n_5003),
.Y(n_6419)
);

CKINVDCx20_ASAP7_75t_R g6420 ( 
.A(n_5681),
.Y(n_6420)
);

BUFx12f_ASAP7_75t_L g6421 ( 
.A(n_5337),
.Y(n_6421)
);

AOI21xp5_ASAP7_75t_L g6422 ( 
.A1(n_5409),
.A2(n_5072),
.B(n_5003),
.Y(n_6422)
);

NAND2x1p5_ASAP7_75t_L g6423 ( 
.A(n_5425),
.B(n_5060),
.Y(n_6423)
);

AND2x4_ASAP7_75t_SL g6424 ( 
.A(n_5216),
.B(n_5060),
.Y(n_6424)
);

BUFx3_ASAP7_75t_L g6425 ( 
.A(n_5246),
.Y(n_6425)
);

AOI21xp5_ASAP7_75t_L g6426 ( 
.A1(n_5413),
.A2(n_5072),
.B(n_5001),
.Y(n_6426)
);

INVxp67_ASAP7_75t_L g6427 ( 
.A(n_5391),
.Y(n_6427)
);

A2O1A1Ixp33_ASAP7_75t_L g6428 ( 
.A1(n_5512),
.A2(n_5001),
.B(n_5041),
.C(n_4935),
.Y(n_6428)
);

HB1xp67_ASAP7_75t_L g6429 ( 
.A(n_5159),
.Y(n_6429)
);

BUFx12f_ASAP7_75t_L g6430 ( 
.A(n_5338),
.Y(n_6430)
);

OAI22xp5_ASAP7_75t_L g6431 ( 
.A1(n_5117),
.A2(n_4918),
.B1(n_4985),
.B2(n_4935),
.Y(n_6431)
);

OR2x2_ASAP7_75t_L g6432 ( 
.A(n_5391),
.B(n_5013),
.Y(n_6432)
);

AND2x6_ASAP7_75t_L g6433 ( 
.A(n_5151),
.B(n_4985),
.Y(n_6433)
);

INVx2_ASAP7_75t_SL g6434 ( 
.A(n_5762),
.Y(n_6434)
);

OAI22xp5_ASAP7_75t_L g6435 ( 
.A1(n_5388),
.A2(n_5041),
.B1(n_4948),
.B2(n_4950),
.Y(n_6435)
);

NOR2xp33_ASAP7_75t_L g6436 ( 
.A(n_5363),
.B(n_5038),
.Y(n_6436)
);

O2A1O1Ixp33_ASAP7_75t_L g6437 ( 
.A1(n_5563),
.A2(n_4983),
.B(n_5033),
.C(n_5037),
.Y(n_6437)
);

AND2x6_ASAP7_75t_L g6438 ( 
.A(n_5151),
.B(n_4983),
.Y(n_6438)
);

INVx4_ASAP7_75t_L g6439 ( 
.A(n_5247),
.Y(n_6439)
);

NAND2x1p5_ASAP7_75t_L g6440 ( 
.A(n_5425),
.B(n_5038),
.Y(n_6440)
);

HB1xp67_ASAP7_75t_L g6441 ( 
.A(n_5162),
.Y(n_6441)
);

BUFx3_ASAP7_75t_L g6442 ( 
.A(n_5247),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_L g6443 ( 
.A(n_5765),
.B(n_5033),
.Y(n_6443)
);

AOI21xp5_ASAP7_75t_L g6444 ( 
.A1(n_5414),
.A2(n_5037),
.B(n_5038),
.Y(n_6444)
);

AOI21xp5_ASAP7_75t_L g6445 ( 
.A1(n_5414),
.A2(n_4787),
.B(n_5426),
.Y(n_6445)
);

NOR2xp33_ASAP7_75t_L g6446 ( 
.A(n_5571),
.B(n_5369),
.Y(n_6446)
);

AOI21xp5_ASAP7_75t_L g6447 ( 
.A1(n_5414),
.A2(n_4787),
.B(n_5426),
.Y(n_6447)
);

AOI22xp5_ASAP7_75t_L g6448 ( 
.A1(n_5388),
.A2(n_4787),
.B1(n_5367),
.B2(n_5383),
.Y(n_6448)
);

NOR2xp67_ASAP7_75t_L g6449 ( 
.A(n_5239),
.B(n_4787),
.Y(n_6449)
);

INVx5_ASAP7_75t_L g6450 ( 
.A(n_5567),
.Y(n_6450)
);

OAI22xp5_ASAP7_75t_L g6451 ( 
.A1(n_5704),
.A2(n_4787),
.B1(n_5777),
.B2(n_5670),
.Y(n_6451)
);

OR2x2_ASAP7_75t_SL g6452 ( 
.A(n_5173),
.B(n_5142),
.Y(n_6452)
);

BUFx12f_ASAP7_75t_L g6453 ( 
.A(n_5338),
.Y(n_6453)
);

BUFx10_ASAP7_75t_L g6454 ( 
.A(n_5740),
.Y(n_6454)
);

OR2x6_ASAP7_75t_L g6455 ( 
.A(n_5213),
.B(n_5242),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_5768),
.B(n_5213),
.Y(n_6456)
);

CKINVDCx5p33_ASAP7_75t_R g6457 ( 
.A(n_5269),
.Y(n_6457)
);

NAND2xp5_ASAP7_75t_SL g6458 ( 
.A(n_5629),
.B(n_5351),
.Y(n_6458)
);

NOR2xp67_ASAP7_75t_L g6459 ( 
.A(n_5264),
.B(n_5768),
.Y(n_6459)
);

INVx2_ASAP7_75t_SL g6460 ( 
.A(n_5768),
.Y(n_6460)
);

AOI21xp5_ASAP7_75t_L g6461 ( 
.A1(n_5426),
.A2(n_5460),
.B(n_5449),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_5285),
.Y(n_6462)
);

AOI21xp5_ASAP7_75t_L g6463 ( 
.A1(n_5449),
.A2(n_5474),
.B(n_5460),
.Y(n_6463)
);

AOI22xp33_ASAP7_75t_L g6464 ( 
.A1(n_5584),
.A2(n_5367),
.B1(n_5383),
.B2(n_5493),
.Y(n_6464)
);

AND2x4_ASAP7_75t_L g6465 ( 
.A(n_5768),
.B(n_5213),
.Y(n_6465)
);

INVx2_ASAP7_75t_SL g6466 ( 
.A(n_5768),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_5285),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_5301),
.Y(n_6468)
);

AND2x2_ASAP7_75t_L g6469 ( 
.A(n_5360),
.B(n_5366),
.Y(n_6469)
);

BUFx6f_ASAP7_75t_L g6470 ( 
.A(n_5781),
.Y(n_6470)
);

OAI22xp5_ASAP7_75t_L g6471 ( 
.A1(n_5670),
.A2(n_5777),
.B1(n_5704),
.B2(n_5465),
.Y(n_6471)
);

AOI22xp33_ASAP7_75t_SL g6472 ( 
.A1(n_5440),
.A2(n_5465),
.B1(n_5418),
.B2(n_5584),
.Y(n_6472)
);

OAI22xp5_ASAP7_75t_L g6473 ( 
.A1(n_5670),
.A2(n_5704),
.B1(n_5777),
.B2(n_5440),
.Y(n_6473)
);

OR2x2_ASAP7_75t_SL g6474 ( 
.A(n_5173),
.B(n_5142),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_5765),
.B(n_5532),
.Y(n_6475)
);

A2O1A1Ixp33_ASAP7_75t_L g6476 ( 
.A1(n_5222),
.A2(n_5223),
.B(n_5589),
.C(n_5274),
.Y(n_6476)
);

NOR2xp33_ASAP7_75t_L g6477 ( 
.A(n_5571),
.B(n_5369),
.Y(n_6477)
);

NOR2xp33_ASAP7_75t_SL g6478 ( 
.A(n_5345),
.B(n_5358),
.Y(n_6478)
);

INVx2_ASAP7_75t_SL g6479 ( 
.A(n_5768),
.Y(n_6479)
);

BUFx6f_ASAP7_75t_L g6480 ( 
.A(n_5781),
.Y(n_6480)
);

AOI21xp5_ASAP7_75t_L g6481 ( 
.A1(n_5449),
.A2(n_5474),
.B(n_5460),
.Y(n_6481)
);

NAND2x1p5_ASAP7_75t_L g6482 ( 
.A(n_5425),
.B(n_5296),
.Y(n_6482)
);

A2O1A1Ixp33_ASAP7_75t_L g6483 ( 
.A1(n_5223),
.A2(n_5589),
.B(n_5274),
.C(n_5623),
.Y(n_6483)
);

AOI21xp5_ASAP7_75t_L g6484 ( 
.A1(n_5474),
.A2(n_5482),
.B(n_5477),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_5532),
.B(n_5594),
.Y(n_6485)
);

NOR2xp33_ASAP7_75t_SL g6486 ( 
.A(n_5345),
.B(n_5358),
.Y(n_6486)
);

AOI22xp33_ASAP7_75t_L g6487 ( 
.A1(n_5383),
.A2(n_5493),
.B1(n_5325),
.B2(n_5436),
.Y(n_6487)
);

BUFx3_ASAP7_75t_L g6488 ( 
.A(n_5247),
.Y(n_6488)
);

AOI22xp33_ASAP7_75t_L g6489 ( 
.A1(n_5493),
.A2(n_5436),
.B1(n_5418),
.B2(n_5153),
.Y(n_6489)
);

BUFx12f_ASAP7_75t_L g6490 ( 
.A(n_5558),
.Y(n_6490)
);

NOR2xp67_ASAP7_75t_SL g6491 ( 
.A(n_5247),
.B(n_5295),
.Y(n_6491)
);

A2O1A1Ixp33_ASAP7_75t_L g6492 ( 
.A1(n_5623),
.A2(n_5503),
.B(n_5527),
.C(n_5534),
.Y(n_6492)
);

BUFx12f_ASAP7_75t_L g6493 ( 
.A(n_5558),
.Y(n_6493)
);

OAI22xp5_ASAP7_75t_L g6494 ( 
.A1(n_5670),
.A2(n_5704),
.B1(n_5777),
.B2(n_5378),
.Y(n_6494)
);

AOI22xp5_ASAP7_75t_L g6495 ( 
.A1(n_5447),
.A2(n_5503),
.B1(n_5534),
.B2(n_5436),
.Y(n_6495)
);

AND2x2_ASAP7_75t_L g6496 ( 
.A(n_5360),
.B(n_5366),
.Y(n_6496)
);

A2O1A1Ixp33_ASAP7_75t_SL g6497 ( 
.A1(n_5362),
.A2(n_5448),
.B(n_5450),
.C(n_5779),
.Y(n_6497)
);

OA21x2_ASAP7_75t_L g6498 ( 
.A1(n_5339),
.A2(n_5132),
.B(n_5773),
.Y(n_6498)
);

AND2x4_ASAP7_75t_L g6499 ( 
.A(n_5768),
.B(n_5213),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_SL g6500 ( 
.A(n_5629),
.B(n_5544),
.Y(n_6500)
);

AOI21xp5_ASAP7_75t_L g6501 ( 
.A1(n_5477),
.A2(n_5484),
.B(n_5482),
.Y(n_6501)
);

INVxp67_ASAP7_75t_SL g6502 ( 
.A(n_5490),
.Y(n_6502)
);

AO32x2_ASAP7_75t_L g6503 ( 
.A1(n_5566),
.A2(n_5527),
.A3(n_5650),
.B1(n_5676),
.B2(n_5684),
.Y(n_6503)
);

CKINVDCx11_ASAP7_75t_R g6504 ( 
.A(n_5123),
.Y(n_6504)
);

NAND2xp5_ASAP7_75t_L g6505 ( 
.A(n_5596),
.B(n_5327),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_5327),
.B(n_5757),
.Y(n_6506)
);

AND2x2_ASAP7_75t_SL g6507 ( 
.A(n_5644),
.B(n_5741),
.Y(n_6507)
);

OAI22xp33_ASAP7_75t_L g6508 ( 
.A1(n_5534),
.A2(n_5571),
.B1(n_5646),
.B2(n_5358),
.Y(n_6508)
);

AOI21xp5_ASAP7_75t_L g6509 ( 
.A1(n_5477),
.A2(n_5484),
.B(n_5482),
.Y(n_6509)
);

AOI21xp5_ASAP7_75t_L g6510 ( 
.A1(n_5484),
.A2(n_5499),
.B(n_5567),
.Y(n_6510)
);

AOI22xp33_ASAP7_75t_L g6511 ( 
.A1(n_5153),
.A2(n_5173),
.B1(n_5394),
.B2(n_5429),
.Y(n_6511)
);

INVx2_ASAP7_75t_SL g6512 ( 
.A(n_5768),
.Y(n_6512)
);

AOI21xp5_ASAP7_75t_L g6513 ( 
.A1(n_5499),
.A2(n_5590),
.B(n_5567),
.Y(n_6513)
);

NAND2xp5_ASAP7_75t_L g6514 ( 
.A(n_5327),
.B(n_5757),
.Y(n_6514)
);

AND2x2_ASAP7_75t_L g6515 ( 
.A(n_5360),
.B(n_5366),
.Y(n_6515)
);

CKINVDCx11_ASAP7_75t_R g6516 ( 
.A(n_5123),
.Y(n_6516)
);

NAND2xp5_ASAP7_75t_L g6517 ( 
.A(n_5757),
.B(n_5208),
.Y(n_6517)
);

BUFx6f_ASAP7_75t_L g6518 ( 
.A(n_5658),
.Y(n_6518)
);

NOR2xp33_ASAP7_75t_L g6519 ( 
.A(n_5550),
.B(n_5552),
.Y(n_6519)
);

OAI22xp5_ASAP7_75t_L g6520 ( 
.A1(n_5378),
.A2(n_5561),
.B1(n_5718),
.B2(n_5760),
.Y(n_6520)
);

BUFx6f_ASAP7_75t_L g6521 ( 
.A(n_5781),
.Y(n_6521)
);

AND2x2_ASAP7_75t_SL g6522 ( 
.A(n_5644),
.B(n_5741),
.Y(n_6522)
);

AND2x4_ASAP7_75t_L g6523 ( 
.A(n_5768),
.B(n_5213),
.Y(n_6523)
);

BUFx10_ASAP7_75t_L g6524 ( 
.A(n_5740),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_L g6525 ( 
.A(n_5208),
.B(n_5211),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_L g6526 ( 
.A(n_5211),
.B(n_5291),
.Y(n_6526)
);

A2O1A1Ixp33_ASAP7_75t_L g6527 ( 
.A1(n_5527),
.A2(n_5646),
.B(n_5103),
.C(n_5517),
.Y(n_6527)
);

AOI21xp5_ASAP7_75t_L g6528 ( 
.A1(n_5499),
.A2(n_5590),
.B(n_5567),
.Y(n_6528)
);

OAI22xp5_ASAP7_75t_L g6529 ( 
.A1(n_5561),
.A2(n_5760),
.B1(n_5761),
.B2(n_5718),
.Y(n_6529)
);

AND2x4_ASAP7_75t_L g6530 ( 
.A(n_5207),
.B(n_5226),
.Y(n_6530)
);

AOI21xp5_ASAP7_75t_L g6531 ( 
.A1(n_5567),
.A2(n_5590),
.B(n_5352),
.Y(n_6531)
);

OAI21xp5_ASAP7_75t_L g6532 ( 
.A1(n_5362),
.A2(n_5450),
.B(n_5448),
.Y(n_6532)
);

BUFx3_ASAP7_75t_L g6533 ( 
.A(n_5295),
.Y(n_6533)
);

BUFx2_ASAP7_75t_L g6534 ( 
.A(n_5116),
.Y(n_6534)
);

AND2x4_ASAP7_75t_L g6535 ( 
.A(n_5207),
.B(n_5226),
.Y(n_6535)
);

AND2x2_ASAP7_75t_L g6536 ( 
.A(n_5360),
.B(n_5366),
.Y(n_6536)
);

NAND2xp5_ASAP7_75t_L g6537 ( 
.A(n_5291),
.B(n_5297),
.Y(n_6537)
);

CKINVDCx11_ASAP7_75t_R g6538 ( 
.A(n_5123),
.Y(n_6538)
);

NAND2xp33_ASAP7_75t_L g6539 ( 
.A(n_5456),
.B(n_5710),
.Y(n_6539)
);

OA21x2_ASAP7_75t_L g6540 ( 
.A1(n_5132),
.A2(n_5773),
.B(n_5142),
.Y(n_6540)
);

OR2x2_ASAP7_75t_L g6541 ( 
.A(n_5642),
.B(n_5645),
.Y(n_6541)
);

OR2x2_ASAP7_75t_L g6542 ( 
.A(n_5642),
.B(n_5645),
.Y(n_6542)
);

OAI21x1_ASAP7_75t_L g6543 ( 
.A1(n_5468),
.A2(n_5392),
.B(n_5251),
.Y(n_6543)
);

AND2x2_ASAP7_75t_L g6544 ( 
.A(n_5580),
.B(n_5108),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_5580),
.B(n_5108),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_5291),
.B(n_5297),
.Y(n_6546)
);

AOI21xp33_ASAP7_75t_SL g6547 ( 
.A1(n_5547),
.A2(n_5708),
.B(n_5203),
.Y(n_6547)
);

BUFx6f_ASAP7_75t_L g6548 ( 
.A(n_5781),
.Y(n_6548)
);

AND2x4_ASAP7_75t_L g6549 ( 
.A(n_5207),
.B(n_5226),
.Y(n_6549)
);

AOI21xp5_ASAP7_75t_L g6550 ( 
.A1(n_5567),
.A2(n_5590),
.B(n_5352),
.Y(n_6550)
);

NAND2xp5_ASAP7_75t_L g6551 ( 
.A(n_5297),
.B(n_5298),
.Y(n_6551)
);

CKINVDCx5p33_ASAP7_75t_R g6552 ( 
.A(n_5308),
.Y(n_6552)
);

NOR3xp33_ASAP7_75t_L g6553 ( 
.A(n_5461),
.B(n_5287),
.C(n_5164),
.Y(n_6553)
);

BUFx2_ASAP7_75t_L g6554 ( 
.A(n_5116),
.Y(n_6554)
);

HB1xp67_ASAP7_75t_L g6555 ( 
.A(n_5162),
.Y(n_6555)
);

NOR2xp33_ASAP7_75t_L g6556 ( 
.A(n_5550),
.B(n_5552),
.Y(n_6556)
);

NOR2xp33_ASAP7_75t_L g6557 ( 
.A(n_5583),
.B(n_5588),
.Y(n_6557)
);

AOI21xp5_ASAP7_75t_L g6558 ( 
.A1(n_5567),
.A2(n_5590),
.B(n_5352),
.Y(n_6558)
);

AOI22xp33_ASAP7_75t_L g6559 ( 
.A1(n_5153),
.A2(n_5394),
.B1(n_5429),
.B2(n_5544),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_5091),
.Y(n_6560)
);

BUFx2_ASAP7_75t_L g6561 ( 
.A(n_5116),
.Y(n_6561)
);

NAND2xp5_ASAP7_75t_L g6562 ( 
.A(n_5298),
.B(n_5316),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_5091),
.Y(n_6563)
);

NOR2xp67_ASAP7_75t_SL g6564 ( 
.A(n_5295),
.B(n_5311),
.Y(n_6564)
);

AOI21xp5_ASAP7_75t_L g6565 ( 
.A1(n_5590),
.A2(n_5352),
.B(n_5336),
.Y(n_6565)
);

AOI21xp5_ASAP7_75t_L g6566 ( 
.A1(n_5590),
.A2(n_5352),
.B(n_5336),
.Y(n_6566)
);

OR2x2_ASAP7_75t_L g6567 ( 
.A(n_5642),
.B(n_5645),
.Y(n_6567)
);

AND2x4_ASAP7_75t_L g6568 ( 
.A(n_5207),
.B(n_5226),
.Y(n_6568)
);

INVx5_ASAP7_75t_L g6569 ( 
.A(n_5590),
.Y(n_6569)
);

BUFx2_ASAP7_75t_L g6570 ( 
.A(n_5116),
.Y(n_6570)
);

OAI22xp5_ASAP7_75t_L g6571 ( 
.A1(n_5718),
.A2(n_5760),
.B1(n_5761),
.B2(n_5586),
.Y(n_6571)
);

NAND2x1_ASAP7_75t_L g6572 ( 
.A(n_5242),
.B(n_5249),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_5091),
.Y(n_6573)
);

AOI21xp5_ASAP7_75t_L g6574 ( 
.A1(n_5336),
.A2(n_5389),
.B(n_5352),
.Y(n_6574)
);

AOI21x1_ASAP7_75t_L g6575 ( 
.A1(n_5392),
.A2(n_5468),
.B(n_5251),
.Y(n_6575)
);

O2A1O1Ixp33_ASAP7_75t_L g6576 ( 
.A1(n_5517),
.A2(n_5569),
.B(n_5629),
.C(n_5570),
.Y(n_6576)
);

OR2x2_ASAP7_75t_L g6577 ( 
.A(n_5645),
.B(n_5769),
.Y(n_6577)
);

CKINVDCx5p33_ASAP7_75t_R g6578 ( 
.A(n_5308),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5097),
.Y(n_6579)
);

AOI21xp33_ASAP7_75t_SL g6580 ( 
.A1(n_5547),
.A2(n_5708),
.B(n_5445),
.Y(n_6580)
);

BUFx2_ASAP7_75t_L g6581 ( 
.A(n_5116),
.Y(n_6581)
);

AOI21xp5_ASAP7_75t_L g6582 ( 
.A1(n_5336),
.A2(n_5389),
.B(n_5352),
.Y(n_6582)
);

CKINVDCx20_ASAP7_75t_R g6583 ( 
.A(n_5508),
.Y(n_6583)
);

OAI22xp5_ASAP7_75t_L g6584 ( 
.A1(n_5718),
.A2(n_5760),
.B1(n_5761),
.B2(n_5586),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_5097),
.Y(n_6585)
);

OAI31xp33_ASAP7_75t_SL g6586 ( 
.A1(n_5517),
.A2(n_5511),
.A3(n_5638),
.B(n_5692),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_5097),
.Y(n_6587)
);

HB1xp67_ASAP7_75t_L g6588 ( 
.A(n_5200),
.Y(n_6588)
);

AND2x4_ASAP7_75t_L g6589 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6589)
);

OAI22xp33_ASAP7_75t_L g6590 ( 
.A1(n_5646),
.A2(n_5626),
.B1(n_5761),
.B2(n_5394),
.Y(n_6590)
);

NOR2xp33_ASAP7_75t_L g6591 ( 
.A(n_5583),
.B(n_5588),
.Y(n_6591)
);

BUFx6f_ASAP7_75t_L g6592 ( 
.A(n_5658),
.Y(n_6592)
);

AOI21xp5_ASAP7_75t_L g6593 ( 
.A1(n_5336),
.A2(n_5389),
.B(n_5352),
.Y(n_6593)
);

NAND2xp5_ASAP7_75t_L g6594 ( 
.A(n_5298),
.B(n_5316),
.Y(n_6594)
);

INVx6_ASAP7_75t_SL g6595 ( 
.A(n_5242),
.Y(n_6595)
);

BUFx12f_ASAP7_75t_L g6596 ( 
.A(n_5625),
.Y(n_6596)
);

BUFx6f_ASAP7_75t_L g6597 ( 
.A(n_5658),
.Y(n_6597)
);

AND2x4_ASAP7_75t_L g6598 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6598)
);

OAI22xp5_ASAP7_75t_L g6599 ( 
.A1(n_5647),
.A2(n_5643),
.B1(n_5591),
.B2(n_5626),
.Y(n_6599)
);

AND2x2_ASAP7_75t_L g6600 ( 
.A(n_5580),
.B(n_5108),
.Y(n_6600)
);

INVx3_ASAP7_75t_SL g6601 ( 
.A(n_5445),
.Y(n_6601)
);

AND2x4_ASAP7_75t_L g6602 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6602)
);

CKINVDCx5p33_ASAP7_75t_R g6603 ( 
.A(n_5330),
.Y(n_6603)
);

AOI22xp33_ASAP7_75t_L g6604 ( 
.A1(n_5394),
.A2(n_5511),
.B1(n_5569),
.B2(n_5164),
.Y(n_6604)
);

INVx1_ASAP7_75t_SL g6605 ( 
.A(n_5310),
.Y(n_6605)
);

BUFx3_ASAP7_75t_L g6606 ( 
.A(n_5295),
.Y(n_6606)
);

AOI21xp5_ASAP7_75t_L g6607 ( 
.A1(n_5336),
.A2(n_5410),
.B(n_5389),
.Y(n_6607)
);

OR2x2_ASAP7_75t_L g6608 ( 
.A(n_5769),
.B(n_5328),
.Y(n_6608)
);

NAND2xp5_ASAP7_75t_L g6609 ( 
.A(n_5316),
.B(n_5684),
.Y(n_6609)
);

A2O1A1Ixp33_ASAP7_75t_L g6610 ( 
.A1(n_5103),
.A2(n_5511),
.B(n_5569),
.C(n_5570),
.Y(n_6610)
);

BUFx12f_ASAP7_75t_L g6611 ( 
.A(n_5625),
.Y(n_6611)
);

AOI22xp5_ASAP7_75t_L g6612 ( 
.A1(n_5447),
.A2(n_5638),
.B1(n_5626),
.B2(n_5692),
.Y(n_6612)
);

AOI21xp5_ASAP7_75t_L g6613 ( 
.A1(n_5336),
.A2(n_5410),
.B(n_5389),
.Y(n_6613)
);

AND2x4_ASAP7_75t_L g6614 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_5615),
.Y(n_6615)
);

AOI21xp5_ASAP7_75t_L g6616 ( 
.A1(n_5336),
.A2(n_5410),
.B(n_5389),
.Y(n_6616)
);

OAI22xp5_ASAP7_75t_L g6617 ( 
.A1(n_5647),
.A2(n_5643),
.B1(n_5591),
.B2(n_5673),
.Y(n_6617)
);

OAI22xp5_ASAP7_75t_L g6618 ( 
.A1(n_5673),
.A2(n_5570),
.B1(n_5565),
.B2(n_5687),
.Y(n_6618)
);

NAND2xp5_ASAP7_75t_L g6619 ( 
.A(n_5684),
.B(n_5686),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_SL g6620 ( 
.A(n_5525),
.B(n_5696),
.Y(n_6620)
);

OAI21xp5_ASAP7_75t_L g6621 ( 
.A1(n_5287),
.A2(n_5164),
.B(n_5157),
.Y(n_6621)
);

OR2x2_ASAP7_75t_L g6622 ( 
.A(n_5769),
.B(n_5328),
.Y(n_6622)
);

AND2x4_ASAP7_75t_L g6623 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6623)
);

INVx4_ASAP7_75t_L g6624 ( 
.A(n_5311),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_5615),
.Y(n_6625)
);

NOR3xp33_ASAP7_75t_L g6626 ( 
.A(n_5287),
.B(n_5157),
.C(n_5382),
.Y(n_6626)
);

AOI22xp33_ASAP7_75t_SL g6627 ( 
.A1(n_5644),
.A2(n_5403),
.B1(n_5741),
.B2(n_5541),
.Y(n_6627)
);

INVx6_ASAP7_75t_L g6628 ( 
.A(n_5279),
.Y(n_6628)
);

NAND3xp33_ASAP7_75t_L g6629 ( 
.A(n_5157),
.B(n_5469),
.C(n_5403),
.Y(n_6629)
);

AND2x2_ASAP7_75t_L g6630 ( 
.A(n_5580),
.B(n_5108),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_5110),
.B(n_5553),
.Y(n_6631)
);

AND2x2_ASAP7_75t_L g6632 ( 
.A(n_5110),
.B(n_5553),
.Y(n_6632)
);

AND2x4_ASAP7_75t_L g6633 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6633)
);

OR2x2_ASAP7_75t_L g6634 ( 
.A(n_5328),
.B(n_5332),
.Y(n_6634)
);

AOI21xp5_ASAP7_75t_L g6635 ( 
.A1(n_5389),
.A2(n_5410),
.B(n_5764),
.Y(n_6635)
);

AOI22xp5_ASAP7_75t_L g6636 ( 
.A1(n_5597),
.A2(n_5564),
.B1(n_5607),
.B2(n_5095),
.Y(n_6636)
);

AND2x2_ASAP7_75t_L g6637 ( 
.A(n_5110),
.B(n_5553),
.Y(n_6637)
);

BUFx6f_ASAP7_75t_L g6638 ( 
.A(n_5658),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_5156),
.B(n_5163),
.Y(n_6639)
);

NOR2xp33_ASAP7_75t_L g6640 ( 
.A(n_5614),
.B(n_5578),
.Y(n_6640)
);

OAI321xp33_ASAP7_75t_L g6641 ( 
.A1(n_5779),
.A2(n_5518),
.A3(n_5469),
.B1(n_5564),
.B2(n_5382),
.C(n_5678),
.Y(n_6641)
);

INVx6_ASAP7_75t_L g6642 ( 
.A(n_5279),
.Y(n_6642)
);

NAND2xp5_ASAP7_75t_L g6643 ( 
.A(n_5686),
.B(n_5709),
.Y(n_6643)
);

NAND2xp5_ASAP7_75t_L g6644 ( 
.A(n_5686),
.B(n_5709),
.Y(n_6644)
);

O2A1O1Ixp33_ASAP7_75t_L g6645 ( 
.A1(n_5564),
.A2(n_5779),
.B(n_5746),
.C(n_5092),
.Y(n_6645)
);

NOR2xp67_ASAP7_75t_L g6646 ( 
.A(n_5111),
.B(n_5395),
.Y(n_6646)
);

AND2x2_ASAP7_75t_L g6647 ( 
.A(n_5110),
.B(n_5553),
.Y(n_6647)
);

NAND2xp33_ASAP7_75t_L g6648 ( 
.A(n_5710),
.B(n_5488),
.Y(n_6648)
);

NOR2xp67_ASAP7_75t_L g6649 ( 
.A(n_5111),
.B(n_5689),
.Y(n_6649)
);

O2A1O1Ixp33_ASAP7_75t_L g6650 ( 
.A1(n_5092),
.A2(n_5764),
.B(n_5678),
.C(n_5566),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_5556),
.B(n_5573),
.Y(n_6651)
);

INVxp67_ASAP7_75t_L g6652 ( 
.A(n_5634),
.Y(n_6652)
);

OAI22xp5_ASAP7_75t_L g6653 ( 
.A1(n_5673),
.A2(n_5565),
.B1(n_5687),
.B2(n_5605),
.Y(n_6653)
);

INVxp67_ASAP7_75t_SL g6654 ( 
.A(n_5559),
.Y(n_6654)
);

NAND2xp5_ASAP7_75t_L g6655 ( 
.A(n_5709),
.B(n_5737),
.Y(n_6655)
);

AO32x2_ASAP7_75t_L g6656 ( 
.A1(n_5566),
.A2(n_5676),
.A3(n_5650),
.B1(n_5772),
.B2(n_5737),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_5737),
.B(n_5772),
.Y(n_6657)
);

OAI21xp33_ASAP7_75t_L g6658 ( 
.A1(n_5382),
.A2(n_5403),
.B(n_5386),
.Y(n_6658)
);

CKINVDCx5p33_ASAP7_75t_R g6659 ( 
.A(n_5330),
.Y(n_6659)
);

NOR2xp33_ASAP7_75t_L g6660 ( 
.A(n_5614),
.B(n_5578),
.Y(n_6660)
);

AOI21xp5_ASAP7_75t_L g6661 ( 
.A1(n_5389),
.A2(n_5410),
.B(n_5132),
.Y(n_6661)
);

BUFx3_ASAP7_75t_L g6662 ( 
.A(n_5311),
.Y(n_6662)
);

AOI22xp33_ASAP7_75t_L g6663 ( 
.A1(n_5538),
.A2(n_5525),
.B1(n_5644),
.B2(n_5095),
.Y(n_6663)
);

NOR2xp33_ASAP7_75t_L g6664 ( 
.A(n_5578),
.B(n_5603),
.Y(n_6664)
);

INVx4_ASAP7_75t_L g6665 ( 
.A(n_5311),
.Y(n_6665)
);

NAND2xp5_ASAP7_75t_L g6666 ( 
.A(n_5772),
.B(n_5688),
.Y(n_6666)
);

BUFx3_ASAP7_75t_L g6667 ( 
.A(n_5326),
.Y(n_6667)
);

INVx3_ASAP7_75t_SL g6668 ( 
.A(n_5434),
.Y(n_6668)
);

NAND2xp5_ASAP7_75t_L g6669 ( 
.A(n_5688),
.B(n_5690),
.Y(n_6669)
);

AND2x2_ASAP7_75t_SL g6670 ( 
.A(n_5644),
.B(n_5741),
.Y(n_6670)
);

NOR2xp33_ASAP7_75t_L g6671 ( 
.A(n_5603),
.B(n_5610),
.Y(n_6671)
);

AND2x4_ASAP7_75t_L g6672 ( 
.A(n_5179),
.B(n_5191),
.Y(n_6672)
);

NAND2xp5_ASAP7_75t_L g6673 ( 
.A(n_5688),
.B(n_5690),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_5601),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6560),
.Y(n_6675)
);

INVx6_ASAP7_75t_L g6676 ( 
.A(n_5846),
.Y(n_6676)
);

BUFx10_ASAP7_75t_L g6677 ( 
.A(n_6318),
.Y(n_6677)
);

OAI21xp33_ASAP7_75t_L g6678 ( 
.A1(n_5839),
.A2(n_5386),
.B(n_5687),
.Y(n_6678)
);

AOI22xp5_ASAP7_75t_L g6679 ( 
.A1(n_5839),
.A2(n_5607),
.B1(n_5555),
.B2(n_5597),
.Y(n_6679)
);

BUFx8_ASAP7_75t_SL g6680 ( 
.A(n_5905),
.Y(n_6680)
);

INVx3_ASAP7_75t_L g6681 ( 
.A(n_5800),
.Y(n_6681)
);

BUFx3_ASAP7_75t_L g6682 ( 
.A(n_5971),
.Y(n_6682)
);

CKINVDCx5p33_ASAP7_75t_R g6683 ( 
.A(n_6140),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6560),
.Y(n_6684)
);

AOI22xp33_ASAP7_75t_L g6685 ( 
.A1(n_6260),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6685)
);

AOI22xp33_ASAP7_75t_L g6686 ( 
.A1(n_6260),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6563),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6225),
.B(n_5524),
.Y(n_6688)
);

AOI22xp33_ASAP7_75t_L g6689 ( 
.A1(n_6398),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6689)
);

OAI22xp33_ASAP7_75t_L g6690 ( 
.A1(n_5998),
.A2(n_5555),
.B1(n_5597),
.B2(n_5575),
.Y(n_6690)
);

CKINVDCx5p33_ASAP7_75t_R g6691 ( 
.A(n_6140),
.Y(n_6691)
);

CKINVDCx20_ASAP7_75t_R g6692 ( 
.A(n_6142),
.Y(n_6692)
);

OAI21xp5_ASAP7_75t_L g6693 ( 
.A1(n_6476),
.A2(n_5518),
.B(n_5678),
.Y(n_6693)
);

INVx1_ASAP7_75t_SL g6694 ( 
.A(n_6432),
.Y(n_6694)
);

OAI22xp5_ASAP7_75t_L g6695 ( 
.A1(n_6476),
.A2(n_5555),
.B1(n_5538),
.B2(n_5605),
.Y(n_6695)
);

INVx2_ASAP7_75t_SL g6696 ( 
.A(n_5812),
.Y(n_6696)
);

INVx3_ASAP7_75t_L g6697 ( 
.A(n_5800),
.Y(n_6697)
);

OAI22xp33_ASAP7_75t_SL g6698 ( 
.A1(n_6118),
.A2(n_5657),
.B1(n_5667),
.B2(n_5547),
.Y(n_6698)
);

AOI22xp33_ASAP7_75t_SL g6699 ( 
.A1(n_5966),
.A2(n_6398),
.B1(n_5968),
.B2(n_6507),
.Y(n_6699)
);

BUFx6f_ASAP7_75t_L g6700 ( 
.A(n_6054),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_5790),
.Y(n_6701)
);

BUFx3_ASAP7_75t_L g6702 ( 
.A(n_5971),
.Y(n_6702)
);

OAI22xp5_ASAP7_75t_L g6703 ( 
.A1(n_6495),
.A2(n_5708),
.B1(n_5533),
.B2(n_5741),
.Y(n_6703)
);

BUFx2_ASAP7_75t_SL g6704 ( 
.A(n_5828),
.Y(n_6704)
);

INVx5_ASAP7_75t_L g6705 ( 
.A(n_6470),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6563),
.Y(n_6706)
);

BUFx8_ASAP7_75t_L g6707 ( 
.A(n_5809),
.Y(n_6707)
);

OAI22xp5_ASAP7_75t_SL g6708 ( 
.A1(n_5911),
.A2(n_5627),
.B1(n_5533),
.B2(n_5504),
.Y(n_6708)
);

BUFx12f_ASAP7_75t_L g6709 ( 
.A(n_5918),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_6573),
.Y(n_6710)
);

BUFx2_ASAP7_75t_SL g6711 ( 
.A(n_5828),
.Y(n_6711)
);

CKINVDCx16_ASAP7_75t_R g6712 ( 
.A(n_5915),
.Y(n_6712)
);

INVx4_ASAP7_75t_L g6713 ( 
.A(n_5971),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_5790),
.Y(n_6714)
);

AOI22xp33_ASAP7_75t_L g6715 ( 
.A1(n_5841),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_5790),
.Y(n_6716)
);

OAI22xp33_ASAP7_75t_L g6717 ( 
.A1(n_5998),
.A2(n_5575),
.B1(n_5662),
.B2(n_5711),
.Y(n_6717)
);

AOI22xp5_ASAP7_75t_SL g6718 ( 
.A1(n_6056),
.A2(n_5488),
.B1(n_5504),
.B2(n_5548),
.Y(n_6718)
);

CKINVDCx20_ASAP7_75t_R g6719 ( 
.A(n_6142),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_5790),
.Y(n_6720)
);

CKINVDCx11_ASAP7_75t_R g6721 ( 
.A(n_6145),
.Y(n_6721)
);

BUFx2_ASAP7_75t_L g6722 ( 
.A(n_6033),
.Y(n_6722)
);

INVx3_ASAP7_75t_L g6723 ( 
.A(n_5800),
.Y(n_6723)
);

BUFx3_ASAP7_75t_L g6724 ( 
.A(n_6111),
.Y(n_6724)
);

CKINVDCx20_ASAP7_75t_R g6725 ( 
.A(n_6145),
.Y(n_6725)
);

INVx6_ASAP7_75t_L g6726 ( 
.A(n_5846),
.Y(n_6726)
);

INVx6_ASAP7_75t_L g6727 ( 
.A(n_5846),
.Y(n_6727)
);

AOI22xp5_ASAP7_75t_L g6728 ( 
.A1(n_5841),
.A2(n_5525),
.B1(n_5696),
.B2(n_5575),
.Y(n_6728)
);

AOI22xp33_ASAP7_75t_L g6729 ( 
.A1(n_5968),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_5790),
.Y(n_6730)
);

OAI22xp5_ASAP7_75t_L g6731 ( 
.A1(n_6495),
.A2(n_5627),
.B1(n_5667),
.B2(n_5657),
.Y(n_6731)
);

BUFx6f_ASAP7_75t_L g6732 ( 
.A(n_6054),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6573),
.Y(n_6733)
);

OAI22xp5_ASAP7_75t_L g6734 ( 
.A1(n_6115),
.A2(n_5662),
.B1(n_5101),
.B2(n_5610),
.Y(n_6734)
);

INVx6_ASAP7_75t_L g6735 ( 
.A(n_5846),
.Y(n_6735)
);

BUFx10_ASAP7_75t_L g6736 ( 
.A(n_6344),
.Y(n_6736)
);

INVx3_ASAP7_75t_L g6737 ( 
.A(n_5800),
.Y(n_6737)
);

INVx4_ASAP7_75t_L g6738 ( 
.A(n_6111),
.Y(n_6738)
);

INVx4_ASAP7_75t_L g6739 ( 
.A(n_6111),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6579),
.Y(n_6740)
);

CKINVDCx11_ASAP7_75t_R g6741 ( 
.A(n_6134),
.Y(n_6741)
);

CKINVDCx8_ASAP7_75t_R g6742 ( 
.A(n_5915),
.Y(n_6742)
);

INVx4_ASAP7_75t_L g6743 ( 
.A(n_5844),
.Y(n_6743)
);

NAND2x1p5_ASAP7_75t_L g6744 ( 
.A(n_6321),
.B(n_5613),
.Y(n_6744)
);

AOI22xp33_ASAP7_75t_L g6745 ( 
.A1(n_6532),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6745)
);

INVx2_ASAP7_75t_SL g6746 ( 
.A(n_5812),
.Y(n_6746)
);

AOI22xp33_ASAP7_75t_L g6747 ( 
.A1(n_6532),
.A2(n_5347),
.B1(n_5318),
.B2(n_5317),
.Y(n_6747)
);

AND2x4_ASAP7_75t_L g6748 ( 
.A(n_6132),
.B(n_5221),
.Y(n_6748)
);

BUFx3_ASAP7_75t_L g6749 ( 
.A(n_6054),
.Y(n_6749)
);

CKINVDCx20_ASAP7_75t_R g6750 ( 
.A(n_6134),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6579),
.Y(n_6751)
);

OAI22xp5_ASAP7_75t_L g6752 ( 
.A1(n_6115),
.A2(n_5662),
.B1(n_5101),
.B2(n_5610),
.Y(n_6752)
);

AOI22xp33_ASAP7_75t_SL g6753 ( 
.A1(n_5966),
.A2(n_6507),
.B1(n_6670),
.B2(n_6522),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6585),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_5829),
.Y(n_6755)
);

OAI21xp33_ASAP7_75t_L g6756 ( 
.A1(n_6118),
.A2(n_5386),
.B(n_5480),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6225),
.B(n_5524),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6631),
.B(n_5195),
.Y(n_6758)
);

AOI22xp33_ASAP7_75t_SL g6759 ( 
.A1(n_6507),
.A2(n_5541),
.B1(n_5519),
.B2(n_5650),
.Y(n_6759)
);

INVx6_ASAP7_75t_L g6760 ( 
.A(n_5846),
.Y(n_6760)
);

OAI22xp5_ASAP7_75t_L g6761 ( 
.A1(n_6487),
.A2(n_5603),
.B1(n_5572),
.B2(n_5111),
.Y(n_6761)
);

BUFx12f_ASAP7_75t_L g6762 ( 
.A(n_6094),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6585),
.Y(n_6763)
);

OAI22xp5_ASAP7_75t_L g6764 ( 
.A1(n_6487),
.A2(n_5572),
.B1(n_5541),
.B2(n_5519),
.Y(n_6764)
);

BUFx6f_ASAP7_75t_L g6765 ( 
.A(n_6470),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6587),
.Y(n_6766)
);

CKINVDCx20_ASAP7_75t_R g6767 ( 
.A(n_6345),
.Y(n_6767)
);

BUFx12f_ASAP7_75t_L g6768 ( 
.A(n_6104),
.Y(n_6768)
);

OAI22xp33_ASAP7_75t_L g6769 ( 
.A1(n_6478),
.A2(n_5711),
.B1(n_5433),
.B2(n_5572),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6587),
.Y(n_6770)
);

BUFx8_ASAP7_75t_L g6771 ( 
.A(n_5809),
.Y(n_6771)
);

INVx6_ASAP7_75t_L g6772 ( 
.A(n_5953),
.Y(n_6772)
);

OAI22xp33_ASAP7_75t_L g6773 ( 
.A1(n_6478),
.A2(n_5711),
.B1(n_5433),
.B2(n_5519),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_L g6774 ( 
.A(n_6626),
.B(n_5524),
.Y(n_6774)
);

INVx4_ASAP7_75t_L g6775 ( 
.A(n_5844),
.Y(n_6775)
);

CKINVDCx6p67_ASAP7_75t_R g6776 ( 
.A(n_5809),
.Y(n_6776)
);

CKINVDCx5p33_ASAP7_75t_R g6777 ( 
.A(n_6106),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6674),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6674),
.Y(n_6779)
);

OAI22xp5_ASAP7_75t_L g6780 ( 
.A1(n_6405),
.A2(n_6254),
.B1(n_6489),
.B2(n_6483),
.Y(n_6780)
);

BUFx8_ASAP7_75t_L g6781 ( 
.A(n_5840),
.Y(n_6781)
);

AOI22xp33_ASAP7_75t_L g6782 ( 
.A1(n_6553),
.A2(n_5318),
.B1(n_5347),
.B2(n_5317),
.Y(n_6782)
);

CKINVDCx20_ASAP7_75t_R g6783 ( 
.A(n_6345),
.Y(n_6783)
);

OAI22xp33_ASAP7_75t_L g6784 ( 
.A1(n_6486),
.A2(n_5433),
.B1(n_5676),
.B2(n_5318),
.Y(n_6784)
);

BUFx4f_ASAP7_75t_L g6785 ( 
.A(n_5911),
.Y(n_6785)
);

BUFx6f_ASAP7_75t_L g6786 ( 
.A(n_6470),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_5797),
.Y(n_6787)
);

AOI22xp33_ASAP7_75t_SL g6788 ( 
.A1(n_6507),
.A2(n_5317),
.B1(n_5347),
.B2(n_5318),
.Y(n_6788)
);

CKINVDCx5p33_ASAP7_75t_R g6789 ( 
.A(n_6106),
.Y(n_6789)
);

OAI21xp5_ASAP7_75t_L g6790 ( 
.A1(n_6483),
.A2(n_5518),
.B(n_5613),
.Y(n_6790)
);

BUFx6f_ASAP7_75t_L g6791 ( 
.A(n_6470),
.Y(n_6791)
);

INVx1_ASAP7_75t_L g6792 ( 
.A(n_5797),
.Y(n_6792)
);

INVx6_ASAP7_75t_L g6793 ( 
.A(n_5953),
.Y(n_6793)
);

INVx1_ASAP7_75t_SL g6794 ( 
.A(n_6432),
.Y(n_6794)
);

INVx4_ASAP7_75t_L g6795 ( 
.A(n_5844),
.Y(n_6795)
);

AOI22xp33_ASAP7_75t_L g6796 ( 
.A1(n_6553),
.A2(n_5347),
.B1(n_5359),
.B2(n_5317),
.Y(n_6796)
);

INVx3_ASAP7_75t_L g6797 ( 
.A(n_5804),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_5802),
.Y(n_6798)
);

BUFx8_ASAP7_75t_SL g6799 ( 
.A(n_5786),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_5802),
.Y(n_6800)
);

AOI22xp33_ASAP7_75t_L g6801 ( 
.A1(n_6522),
.A2(n_6670),
.B1(n_6472),
.B2(n_6254),
.Y(n_6801)
);

AOI22xp33_ASAP7_75t_L g6802 ( 
.A1(n_6522),
.A2(n_5359),
.B1(n_5433),
.B2(n_5695),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_5807),
.Y(n_6803)
);

CKINVDCx5p33_ASAP7_75t_R g6804 ( 
.A(n_6234),
.Y(n_6804)
);

OAI22xp5_ASAP7_75t_L g6805 ( 
.A1(n_6405),
.A2(n_5690),
.B1(n_5729),
.B2(n_5724),
.Y(n_6805)
);

CKINVDCx5p33_ASAP7_75t_R g6806 ( 
.A(n_6234),
.Y(n_6806)
);

OAI22xp5_ASAP7_75t_L g6807 ( 
.A1(n_6489),
.A2(n_5724),
.B1(n_5743),
.B2(n_5729),
.Y(n_6807)
);

INVx3_ASAP7_75t_L g6808 ( 
.A(n_5804),
.Y(n_6808)
);

AND2x2_ASAP7_75t_L g6809 ( 
.A(n_6631),
.B(n_5195),
.Y(n_6809)
);

AOI22xp33_ASAP7_75t_L g6810 ( 
.A1(n_6522),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6810)
);

INVx2_ASAP7_75t_L g6811 ( 
.A(n_5829),
.Y(n_6811)
);

AOI22xp33_ASAP7_75t_L g6812 ( 
.A1(n_6670),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6812)
);

OR2x2_ASAP7_75t_L g6813 ( 
.A(n_5930),
.B(n_5328),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_5807),
.Y(n_6814)
);

INVx6_ASAP7_75t_L g6815 ( 
.A(n_5953),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_5811),
.Y(n_6816)
);

INVx2_ASAP7_75t_SL g6817 ( 
.A(n_5812),
.Y(n_6817)
);

INVx8_ASAP7_75t_L g6818 ( 
.A(n_6490),
.Y(n_6818)
);

INVx6_ASAP7_75t_L g6819 ( 
.A(n_5953),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_5811),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_5817),
.Y(n_6821)
);

BUFx12f_ASAP7_75t_L g6822 ( 
.A(n_6233),
.Y(n_6822)
);

CKINVDCx11_ASAP7_75t_R g6823 ( 
.A(n_6583),
.Y(n_6823)
);

OAI22xp5_ASAP7_75t_SL g6824 ( 
.A1(n_5911),
.A2(n_5725),
.B1(n_5548),
.B2(n_5530),
.Y(n_6824)
);

AND2x2_ASAP7_75t_L g6825 ( 
.A(n_6631),
.B(n_5195),
.Y(n_6825)
);

AOI22xp33_ASAP7_75t_L g6826 ( 
.A1(n_6670),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_5817),
.Y(n_6827)
);

AOI22xp33_ASAP7_75t_L g6828 ( 
.A1(n_6472),
.A2(n_6261),
.B1(n_6653),
.B2(n_6599),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_5818),
.Y(n_6829)
);

OAI22xp5_ASAP7_75t_L g6830 ( 
.A1(n_6492),
.A2(n_5724),
.B1(n_5743),
.B2(n_5729),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_5829),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_5818),
.Y(n_6832)
);

INVx1_ASAP7_75t_SL g6833 ( 
.A(n_6432),
.Y(n_6833)
);

INVx6_ASAP7_75t_L g6834 ( 
.A(n_5953),
.Y(n_6834)
);

CKINVDCx11_ASAP7_75t_R g6835 ( 
.A(n_6583),
.Y(n_6835)
);

INVx6_ASAP7_75t_L g6836 ( 
.A(n_6383),
.Y(n_6836)
);

AND2x4_ASAP7_75t_SL g6837 ( 
.A(n_5803),
.B(n_5434),
.Y(n_6837)
);

INVx6_ASAP7_75t_L g6838 ( 
.A(n_6383),
.Y(n_6838)
);

OAI22xp5_ASAP7_75t_L g6839 ( 
.A1(n_6492),
.A2(n_5743),
.B1(n_5755),
.B2(n_5753),
.Y(n_6839)
);

BUFx2_ASAP7_75t_SL g6840 ( 
.A(n_5828),
.Y(n_6840)
);

AOI22xp5_ASAP7_75t_L g6841 ( 
.A1(n_6261),
.A2(n_5725),
.B1(n_5289),
.B2(n_5302),
.Y(n_6841)
);

CKINVDCx20_ASAP7_75t_R g6842 ( 
.A(n_6079),
.Y(n_6842)
);

OAI22xp33_ASAP7_75t_L g6843 ( 
.A1(n_6486),
.A2(n_5359),
.B1(n_5289),
.B2(n_5302),
.Y(n_6843)
);

CKINVDCx5p33_ASAP7_75t_R g6844 ( 
.A(n_5819),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_5831),
.Y(n_6845)
);

AOI22xp33_ASAP7_75t_L g6846 ( 
.A1(n_6653),
.A2(n_6599),
.B1(n_6464),
.B2(n_6458),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_5831),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_5832),
.Y(n_6848)
);

AOI22xp33_ASAP7_75t_SL g6849 ( 
.A1(n_6494),
.A2(n_5359),
.B1(n_5620),
.B2(n_5434),
.Y(n_6849)
);

CKINVDCx20_ASAP7_75t_R g6850 ( 
.A(n_6079),
.Y(n_6850)
);

OR2x6_ASAP7_75t_L g6851 ( 
.A(n_6132),
.B(n_5242),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_5832),
.Y(n_6852)
);

AOI22xp33_ASAP7_75t_SL g6853 ( 
.A1(n_6494),
.A2(n_5789),
.B1(n_6617),
.B2(n_6618),
.Y(n_6853)
);

INVx6_ASAP7_75t_L g6854 ( 
.A(n_6383),
.Y(n_6854)
);

AOI22xp33_ASAP7_75t_L g6855 ( 
.A1(n_6464),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6855)
);

BUFx8_ASAP7_75t_L g6856 ( 
.A(n_5840),
.Y(n_6856)
);

INVx4_ASAP7_75t_L g6857 ( 
.A(n_5844),
.Y(n_6857)
);

AOI22xp33_ASAP7_75t_L g6858 ( 
.A1(n_6458),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6858)
);

AO22x1_ASAP7_75t_L g6859 ( 
.A1(n_5911),
.A2(n_5170),
.B1(n_5609),
.B2(n_5593),
.Y(n_6859)
);

CKINVDCx20_ASAP7_75t_R g6860 ( 
.A(n_6411),
.Y(n_6860)
);

BUFx8_ASAP7_75t_L g6861 ( 
.A(n_5840),
.Y(n_6861)
);

INVx1_ASAP7_75t_L g6862 ( 
.A(n_5834),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_5834),
.Y(n_6863)
);

CKINVDCx5p33_ASAP7_75t_R g6864 ( 
.A(n_6367),
.Y(n_6864)
);

INVx2_ASAP7_75t_SL g6865 ( 
.A(n_5812),
.Y(n_6865)
);

BUFx4f_ASAP7_75t_SL g6866 ( 
.A(n_6263),
.Y(n_6866)
);

INVx4_ASAP7_75t_L g6867 ( 
.A(n_5852),
.Y(n_6867)
);

INVx2_ASAP7_75t_SL g6868 ( 
.A(n_5812),
.Y(n_6868)
);

INVxp67_ASAP7_75t_L g6869 ( 
.A(n_5929),
.Y(n_6869)
);

AOI21xp5_ASAP7_75t_SL g6870 ( 
.A1(n_5912),
.A2(n_5500),
.B(n_5740),
.Y(n_6870)
);

AND2x4_ASAP7_75t_L g6871 ( 
.A(n_6132),
.B(n_5221),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_5838),
.Y(n_6872)
);

OAI22xp5_ASAP7_75t_L g6873 ( 
.A1(n_6384),
.A2(n_5753),
.B1(n_5778),
.B2(n_5755),
.Y(n_6873)
);

INVx2_ASAP7_75t_L g6874 ( 
.A(n_5829),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_5838),
.Y(n_6875)
);

AOI22xp33_ASAP7_75t_L g6876 ( 
.A1(n_6508),
.A2(n_5359),
.B1(n_5703),
.B2(n_5695),
.Y(n_6876)
);

INVx1_ASAP7_75t_L g6877 ( 
.A(n_5843),
.Y(n_6877)
);

BUFx2_ASAP7_75t_SL g6878 ( 
.A(n_5877),
.Y(n_6878)
);

AOI22xp33_ASAP7_75t_SL g6879 ( 
.A1(n_5789),
.A2(n_5434),
.B1(n_5620),
.B2(n_5693),
.Y(n_6879)
);

BUFx2_ASAP7_75t_L g6880 ( 
.A(n_6033),
.Y(n_6880)
);

INVx2_ASAP7_75t_L g6881 ( 
.A(n_5829),
.Y(n_6881)
);

BUFx6f_ASAP7_75t_L g6882 ( 
.A(n_6470),
.Y(n_6882)
);

AOI22xp5_ASAP7_75t_L g6883 ( 
.A1(n_6617),
.A2(n_5289),
.B1(n_5302),
.B2(n_5216),
.Y(n_6883)
);

BUFx2_ASAP7_75t_L g6884 ( 
.A(n_6033),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_5843),
.Y(n_6885)
);

OAI22xp5_ASAP7_75t_L g6886 ( 
.A1(n_6384),
.A2(n_5753),
.B1(n_5778),
.B2(n_5755),
.Y(n_6886)
);

AND2x2_ASAP7_75t_L g6887 ( 
.A(n_6632),
.B(n_5248),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_5849),
.Y(n_6888)
);

CKINVDCx5p33_ASAP7_75t_R g6889 ( 
.A(n_6368),
.Y(n_6889)
);

BUFx12f_ASAP7_75t_L g6890 ( 
.A(n_6262),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_5849),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_5863),
.Y(n_6892)
);

AOI22xp5_ASAP7_75t_L g6893 ( 
.A1(n_6508),
.A2(n_5289),
.B1(n_5302),
.B2(n_5216),
.Y(n_6893)
);

INVx1_ASAP7_75t_SL g6894 ( 
.A(n_6243),
.Y(n_6894)
);

AOI22xp33_ASAP7_75t_L g6895 ( 
.A1(n_5960),
.A2(n_6618),
.B1(n_6627),
.B2(n_6620),
.Y(n_6895)
);

NAND2x1p5_ASAP7_75t_L g6896 ( 
.A(n_6321),
.B(n_5618),
.Y(n_6896)
);

INVx1_ASAP7_75t_SL g6897 ( 
.A(n_6243),
.Y(n_6897)
);

AOI22xp33_ASAP7_75t_L g6898 ( 
.A1(n_5960),
.A2(n_5703),
.B1(n_5695),
.B2(n_5216),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_5863),
.Y(n_6899)
);

NAND2xp5_ASAP7_75t_L g6900 ( 
.A(n_6626),
.B(n_6506),
.Y(n_6900)
);

AOI22xp33_ASAP7_75t_SL g6901 ( 
.A1(n_6471),
.A2(n_5434),
.B1(n_5620),
.B2(n_5693),
.Y(n_6901)
);

OAI22xp33_ASAP7_75t_L g6902 ( 
.A1(n_6612),
.A2(n_5289),
.B1(n_5312),
.B2(n_5302),
.Y(n_6902)
);

INVx6_ASAP7_75t_L g6903 ( 
.A(n_6383),
.Y(n_6903)
);

INVx6_ASAP7_75t_L g6904 ( 
.A(n_6383),
.Y(n_6904)
);

OAI22xp33_ASAP7_75t_L g6905 ( 
.A1(n_6612),
.A2(n_5302),
.B1(n_5312),
.B2(n_5703),
.Y(n_6905)
);

OAI22xp33_ASAP7_75t_L g6906 ( 
.A1(n_6243),
.A2(n_5312),
.B1(n_5782),
.B2(n_5778),
.Y(n_6906)
);

OAI21xp33_ASAP7_75t_SL g6907 ( 
.A1(n_5923),
.A2(n_5435),
.B(n_5423),
.Y(n_6907)
);

AOI22xp33_ASAP7_75t_L g6908 ( 
.A1(n_6627),
.A2(n_5312),
.B1(n_5720),
.B2(n_5242),
.Y(n_6908)
);

OAI21xp5_ASAP7_75t_SL g6909 ( 
.A1(n_6586),
.A2(n_5530),
.B(n_5520),
.Y(n_6909)
);

HB1xp67_ASAP7_75t_L g6910 ( 
.A(n_5987),
.Y(n_6910)
);

CKINVDCx20_ASAP7_75t_R g6911 ( 
.A(n_6411),
.Y(n_6911)
);

INVx2_ASAP7_75t_L g6912 ( 
.A(n_5888),
.Y(n_6912)
);

AOI22xp33_ASAP7_75t_SL g6913 ( 
.A1(n_6471),
.A2(n_5434),
.B1(n_5620),
.B2(n_5693),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_5867),
.Y(n_6914)
);

BUFx2_ASAP7_75t_L g6915 ( 
.A(n_6033),
.Y(n_6915)
);

AOI22xp33_ASAP7_75t_L g6916 ( 
.A1(n_6620),
.A2(n_5312),
.B1(n_5720),
.B2(n_5242),
.Y(n_6916)
);

OAI22xp33_ASAP7_75t_L g6917 ( 
.A1(n_6243),
.A2(n_5312),
.B1(n_5782),
.B2(n_5435),
.Y(n_6917)
);

BUFx12f_ASAP7_75t_L g6918 ( 
.A(n_6263),
.Y(n_6918)
);

CKINVDCx20_ASAP7_75t_R g6919 ( 
.A(n_6420),
.Y(n_6919)
);

AOI22xp33_ASAP7_75t_SL g6920 ( 
.A1(n_6473),
.A2(n_5620),
.B1(n_5721),
.B2(n_5248),
.Y(n_6920)
);

AOI22xp33_ASAP7_75t_SL g6921 ( 
.A1(n_6473),
.A2(n_5620),
.B1(n_5721),
.B2(n_5248),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_5888),
.Y(n_6922)
);

BUFx4_ASAP7_75t_R g6923 ( 
.A(n_5852),
.Y(n_6923)
);

INVx2_ASAP7_75t_L g6924 ( 
.A(n_5888),
.Y(n_6924)
);

AND2x2_ASAP7_75t_L g6925 ( 
.A(n_6632),
.B(n_5556),
.Y(n_6925)
);

INVxp67_ASAP7_75t_SL g6926 ( 
.A(n_5987),
.Y(n_6926)
);

BUFx3_ASAP7_75t_L g6927 ( 
.A(n_5852),
.Y(n_6927)
);

OAI22xp5_ASAP7_75t_L g6928 ( 
.A1(n_6384),
.A2(n_5782),
.B1(n_5672),
.B2(n_5435),
.Y(n_6928)
);

OAI22xp5_ASAP7_75t_L g6929 ( 
.A1(n_6527),
.A2(n_5672),
.B1(n_5435),
.B2(n_5423),
.Y(n_6929)
);

NAND2xp5_ASAP7_75t_L g6930 ( 
.A(n_6506),
.B(n_5557),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_5888),
.Y(n_6931)
);

INVx8_ASAP7_75t_L g6932 ( 
.A(n_6490),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_5867),
.Y(n_6933)
);

BUFx8_ASAP7_75t_L g6934 ( 
.A(n_6263),
.Y(n_6934)
);

BUFx3_ASAP7_75t_L g6935 ( 
.A(n_5852),
.Y(n_6935)
);

INVx2_ASAP7_75t_L g6936 ( 
.A(n_5888),
.Y(n_6936)
);

AOI22xp33_ASAP7_75t_L g6937 ( 
.A1(n_6500),
.A2(n_5720),
.B1(n_5242),
.B2(n_5249),
.Y(n_6937)
);

CKINVDCx11_ASAP7_75t_R g6938 ( 
.A(n_6420),
.Y(n_6938)
);

INVx8_ASAP7_75t_L g6939 ( 
.A(n_6490),
.Y(n_6939)
);

AOI22xp33_ASAP7_75t_SL g6940 ( 
.A1(n_6520),
.A2(n_5721),
.B1(n_5187),
.B2(n_5189),
.Y(n_6940)
);

AOI22xp33_ASAP7_75t_L g6941 ( 
.A1(n_6500),
.A2(n_5720),
.B1(n_5249),
.B2(n_5165),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_5873),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_5873),
.Y(n_6943)
);

BUFx2_ASAP7_75t_L g6944 ( 
.A(n_6033),
.Y(n_6944)
);

AOI22xp33_ASAP7_75t_L g6945 ( 
.A1(n_5806),
.A2(n_5720),
.B1(n_5249),
.B2(n_5165),
.Y(n_6945)
);

AND2x2_ASAP7_75t_L g6946 ( 
.A(n_6632),
.B(n_5556),
.Y(n_6946)
);

AOI22xp33_ASAP7_75t_SL g6947 ( 
.A1(n_6520),
.A2(n_5187),
.B1(n_5189),
.B2(n_5423),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_5882),
.Y(n_6948)
);

NAND2x1p5_ASAP7_75t_L g6949 ( 
.A(n_6321),
.B(n_6324),
.Y(n_6949)
);

AOI22xp33_ASAP7_75t_L g6950 ( 
.A1(n_5806),
.A2(n_5720),
.B1(n_5249),
.B2(n_5165),
.Y(n_6950)
);

INVx3_ASAP7_75t_L g6951 ( 
.A(n_5804),
.Y(n_6951)
);

AOI22xp5_ASAP7_75t_L g6952 ( 
.A1(n_6056),
.A2(n_5714),
.B1(n_5341),
.B2(n_5520),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_5882),
.Y(n_6953)
);

BUFx2_ASAP7_75t_SL g6954 ( 
.A(n_5877),
.Y(n_6954)
);

INVx6_ASAP7_75t_L g6955 ( 
.A(n_5803),
.Y(n_6955)
);

OAI22xp5_ASAP7_75t_L g6956 ( 
.A1(n_6527),
.A2(n_5423),
.B1(n_5189),
.B2(n_5187),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_5894),
.Y(n_6957)
);

INVx1_ASAP7_75t_SL g6958 ( 
.A(n_5810),
.Y(n_6958)
);

AOI22xp33_ASAP7_75t_L g6959 ( 
.A1(n_6663),
.A2(n_5826),
.B1(n_5989),
.B2(n_6391),
.Y(n_6959)
);

INVx4_ASAP7_75t_L g6960 ( 
.A(n_6493),
.Y(n_6960)
);

BUFx12f_ASAP7_75t_L g6961 ( 
.A(n_6275),
.Y(n_6961)
);

AND2x4_ASAP7_75t_L g6962 ( 
.A(n_6132),
.B(n_5221),
.Y(n_6962)
);

INVx2_ASAP7_75t_L g6963 ( 
.A(n_5963),
.Y(n_6963)
);

CKINVDCx11_ASAP7_75t_R g6964 ( 
.A(n_6275),
.Y(n_6964)
);

BUFx12f_ASAP7_75t_L g6965 ( 
.A(n_6275),
.Y(n_6965)
);

BUFx6f_ASAP7_75t_L g6966 ( 
.A(n_6470),
.Y(n_6966)
);

AOI22xp33_ASAP7_75t_L g6967 ( 
.A1(n_6663),
.A2(n_5720),
.B1(n_5249),
.B2(n_5165),
.Y(n_6967)
);

NAND2x1p5_ASAP7_75t_L g6968 ( 
.A(n_6321),
.B(n_5618),
.Y(n_6968)
);

BUFx10_ASAP7_75t_L g6969 ( 
.A(n_6350),
.Y(n_6969)
);

OAI22xp5_ASAP7_75t_L g6970 ( 
.A1(n_6610),
.A2(n_5719),
.B1(n_5742),
.B2(n_5633),
.Y(n_6970)
);

INVx4_ASAP7_75t_L g6971 ( 
.A(n_6493),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_5894),
.Y(n_6972)
);

INVx1_ASAP7_75t_SL g6973 ( 
.A(n_5810),
.Y(n_6973)
);

INVx8_ASAP7_75t_L g6974 ( 
.A(n_6493),
.Y(n_6974)
);

AOI22xp33_ASAP7_75t_L g6975 ( 
.A1(n_5826),
.A2(n_5720),
.B1(n_5249),
.B2(n_5165),
.Y(n_6975)
);

INVx6_ASAP7_75t_L g6976 ( 
.A(n_5803),
.Y(n_6976)
);

NAND2xp5_ASAP7_75t_L g6977 ( 
.A(n_6514),
.B(n_5557),
.Y(n_6977)
);

OAI22xp5_ASAP7_75t_L g6978 ( 
.A1(n_6610),
.A2(n_5719),
.B1(n_5742),
.B2(n_5633),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_5901),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_5901),
.Y(n_6980)
);

INVx2_ASAP7_75t_L g6981 ( 
.A(n_5963),
.Y(n_6981)
);

AOI22xp33_ASAP7_75t_SL g6982 ( 
.A1(n_5893),
.A2(n_5092),
.B1(n_5669),
.B2(n_5634),
.Y(n_6982)
);

BUFx6f_ASAP7_75t_L g6983 ( 
.A(n_6470),
.Y(n_6983)
);

AOI22xp33_ASAP7_75t_L g6984 ( 
.A1(n_5989),
.A2(n_6402),
.B1(n_6408),
.B2(n_6391),
.Y(n_6984)
);

INVx4_ASAP7_75t_SL g6985 ( 
.A(n_6161),
.Y(n_6985)
);

INVx3_ASAP7_75t_SL g6986 ( 
.A(n_6356),
.Y(n_6986)
);

AOI22xp33_ASAP7_75t_SL g6987 ( 
.A1(n_5893),
.A2(n_5092),
.B1(n_5669),
.B2(n_5634),
.Y(n_6987)
);

AOI22xp33_ASAP7_75t_SL g6988 ( 
.A1(n_6116),
.A2(n_5092),
.B1(n_5669),
.B2(n_5166),
.Y(n_6988)
);

BUFx12f_ASAP7_75t_L g6989 ( 
.A(n_5939),
.Y(n_6989)
);

AND2x2_ASAP7_75t_L g6990 ( 
.A(n_6637),
.B(n_5556),
.Y(n_6990)
);

AOI22xp33_ASAP7_75t_L g6991 ( 
.A1(n_6391),
.A2(n_5165),
.B1(n_5279),
.B2(n_5177),
.Y(n_6991)
);

INVx6_ASAP7_75t_L g6992 ( 
.A(n_5803),
.Y(n_6992)
);

BUFx4_ASAP7_75t_R g6993 ( 
.A(n_5984),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_5903),
.Y(n_6994)
);

BUFx8_ASAP7_75t_L g6995 ( 
.A(n_5939),
.Y(n_6995)
);

HB1xp67_ASAP7_75t_L g6996 ( 
.A(n_6013),
.Y(n_6996)
);

CKINVDCx5p33_ASAP7_75t_R g6997 ( 
.A(n_5870),
.Y(n_6997)
);

OAI22xp5_ASAP7_75t_L g6998 ( 
.A1(n_6559),
.A2(n_5742),
.B1(n_5719),
.B2(n_5155),
.Y(n_6998)
);

INVxp67_ASAP7_75t_SL g6999 ( 
.A(n_6013),
.Y(n_6999)
);

OR2x2_ASAP7_75t_L g7000 ( 
.A(n_5930),
.B(n_5956),
.Y(n_7000)
);

AOI22xp33_ASAP7_75t_SL g7001 ( 
.A1(n_6116),
.A2(n_5166),
.B1(n_5331),
.B2(n_5326),
.Y(n_7001)
);

INVx5_ASAP7_75t_L g7002 ( 
.A(n_6470),
.Y(n_7002)
);

INVx2_ASAP7_75t_L g7003 ( 
.A(n_5963),
.Y(n_7003)
);

BUFx6f_ASAP7_75t_L g7004 ( 
.A(n_6480),
.Y(n_7004)
);

AOI22xp33_ASAP7_75t_L g7005 ( 
.A1(n_6402),
.A2(n_5148),
.B1(n_5400),
.B2(n_5177),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6637),
.B(n_5573),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_5903),
.Y(n_7007)
);

INVx2_ASAP7_75t_L g7008 ( 
.A(n_5963),
.Y(n_7008)
);

CKINVDCx20_ASAP7_75t_R g7009 ( 
.A(n_6351),
.Y(n_7009)
);

OAI22xp5_ASAP7_75t_L g7010 ( 
.A1(n_6559),
.A2(n_5742),
.B1(n_5719),
.B2(n_5155),
.Y(n_7010)
);

INVx1_ASAP7_75t_SL g7011 ( 
.A(n_5885),
.Y(n_7011)
);

INVx2_ASAP7_75t_L g7012 ( 
.A(n_5963),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6514),
.B(n_5557),
.Y(n_7013)
);

OAI22xp33_ASAP7_75t_L g7014 ( 
.A1(n_6636),
.A2(n_5090),
.B1(n_5104),
.B2(n_5148),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_5909),
.Y(n_7015)
);

AND2x4_ASAP7_75t_L g7016 ( 
.A(n_6132),
.B(n_6589),
.Y(n_7016)
);

CKINVDCx6p67_ASAP7_75t_R g7017 ( 
.A(n_5939),
.Y(n_7017)
);

BUFx4f_ASAP7_75t_SL g7018 ( 
.A(n_6101),
.Y(n_7018)
);

INVx1_ASAP7_75t_SL g7019 ( 
.A(n_5885),
.Y(n_7019)
);

BUFx6f_ASAP7_75t_L g7020 ( 
.A(n_6480),
.Y(n_7020)
);

AND2x2_ASAP7_75t_L g7021 ( 
.A(n_6637),
.B(n_6647),
.Y(n_7021)
);

OAI22xp33_ASAP7_75t_L g7022 ( 
.A1(n_6636),
.A2(n_5090),
.B1(n_5104),
.B2(n_5148),
.Y(n_7022)
);

OAI22xp33_ASAP7_75t_L g7023 ( 
.A1(n_6448),
.A2(n_5090),
.B1(n_5104),
.B2(n_5148),
.Y(n_7023)
);

INVx8_ASAP7_75t_L g7024 ( 
.A(n_6596),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_5909),
.Y(n_7025)
);

AOI22xp33_ASAP7_75t_SL g7026 ( 
.A1(n_5847),
.A2(n_5166),
.B1(n_5331),
.B2(n_5326),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_5910),
.Y(n_7027)
);

CKINVDCx20_ASAP7_75t_R g7028 ( 
.A(n_6351),
.Y(n_7028)
);

AND2x2_ASAP7_75t_L g7029 ( 
.A(n_6647),
.B(n_5573),
.Y(n_7029)
);

BUFx6f_ASAP7_75t_L g7030 ( 
.A(n_6480),
.Y(n_7030)
);

INVx2_ASAP7_75t_L g7031 ( 
.A(n_5974),
.Y(n_7031)
);

BUFx10_ASAP7_75t_L g7032 ( 
.A(n_5886),
.Y(n_7032)
);

CKINVDCx11_ASAP7_75t_R g7033 ( 
.A(n_6358),
.Y(n_7033)
);

AOI22xp33_ASAP7_75t_L g7034 ( 
.A1(n_6402),
.A2(n_5148),
.B1(n_5400),
.B2(n_5177),
.Y(n_7034)
);

BUFx4f_ASAP7_75t_SL g7035 ( 
.A(n_6101),
.Y(n_7035)
);

OAI22xp5_ASAP7_75t_L g7036 ( 
.A1(n_6448),
.A2(n_5155),
.B1(n_5124),
.B2(n_5126),
.Y(n_7036)
);

CKINVDCx20_ASAP7_75t_R g7037 ( 
.A(n_6358),
.Y(n_7037)
);

BUFx4_ASAP7_75t_SL g7038 ( 
.A(n_6373),
.Y(n_7038)
);

OAI22xp5_ASAP7_75t_L g7039 ( 
.A1(n_6511),
.A2(n_5155),
.B1(n_5124),
.B2(n_5126),
.Y(n_7039)
);

BUFx12f_ASAP7_75t_L g7040 ( 
.A(n_6101),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_SL g7041 ( 
.A1(n_5847),
.A2(n_5166),
.B1(n_5331),
.B2(n_5326),
.Y(n_7041)
);

INVx1_ASAP7_75t_SL g7042 ( 
.A(n_5938),
.Y(n_7042)
);

INVx5_ASAP7_75t_L g7043 ( 
.A(n_6480),
.Y(n_7043)
);

INVx3_ASAP7_75t_L g7044 ( 
.A(n_5804),
.Y(n_7044)
);

AOI22xp33_ASAP7_75t_L g7045 ( 
.A1(n_6408),
.A2(n_5148),
.B1(n_5400),
.B2(n_5177),
.Y(n_7045)
);

AOI22xp33_ASAP7_75t_L g7046 ( 
.A1(n_6408),
.A2(n_5400),
.B1(n_5415),
.B2(n_5177),
.Y(n_7046)
);

AOI22xp5_ASAP7_75t_L g7047 ( 
.A1(n_6590),
.A2(n_5714),
.B1(n_5341),
.B2(n_5424),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_5910),
.Y(n_7048)
);

BUFx3_ASAP7_75t_L g7049 ( 
.A(n_6401),
.Y(n_7049)
);

BUFx3_ASAP7_75t_L g7050 ( 
.A(n_6401),
.Y(n_7050)
);

INVx4_ASAP7_75t_L g7051 ( 
.A(n_6596),
.Y(n_7051)
);

AOI22xp33_ASAP7_75t_L g7052 ( 
.A1(n_5850),
.A2(n_5400),
.B1(n_5415),
.B2(n_5177),
.Y(n_7052)
);

CKINVDCx11_ASAP7_75t_R g7053 ( 
.A(n_6197),
.Y(n_7053)
);

NAND2xp5_ASAP7_75t_L g7054 ( 
.A(n_6416),
.B(n_5341),
.Y(n_7054)
);

AOI22xp33_ASAP7_75t_SL g7055 ( 
.A1(n_5868),
.A2(n_5166),
.B1(n_5349),
.B2(n_5331),
.Y(n_7055)
);

BUFx12f_ASAP7_75t_L g7056 ( 
.A(n_6197),
.Y(n_7056)
);

AOI22xp33_ASAP7_75t_SL g7057 ( 
.A1(n_5868),
.A2(n_5166),
.B1(n_5472),
.B2(n_5349),
.Y(n_7057)
);

INVx2_ASAP7_75t_L g7058 ( 
.A(n_5974),
.Y(n_7058)
);

INVx6_ASAP7_75t_L g7059 ( 
.A(n_5803),
.Y(n_7059)
);

OAI21xp5_ASAP7_75t_SL g7060 ( 
.A1(n_6586),
.A2(n_5716),
.B(n_5483),
.Y(n_7060)
);

INVx1_ASAP7_75t_SL g7061 ( 
.A(n_5938),
.Y(n_7061)
);

BUFx8_ASAP7_75t_L g7062 ( 
.A(n_6197),
.Y(n_7062)
);

NAND2x1p5_ASAP7_75t_L g7063 ( 
.A(n_6321),
.B(n_5618),
.Y(n_7063)
);

AOI22xp33_ASAP7_75t_SL g7064 ( 
.A1(n_5787),
.A2(n_5166),
.B1(n_5472),
.B2(n_5349),
.Y(n_7064)
);

OAI22xp5_ASAP7_75t_L g7065 ( 
.A1(n_6511),
.A2(n_5124),
.B1(n_5126),
.B2(n_5107),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_5920),
.Y(n_7066)
);

AOI22xp33_ASAP7_75t_L g7067 ( 
.A1(n_5850),
.A2(n_5415),
.B1(n_5462),
.B2(n_5400),
.Y(n_7067)
);

AOI22xp33_ASAP7_75t_L g7068 ( 
.A1(n_5850),
.A2(n_5462),
.B1(n_5471),
.B2(n_5415),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_5920),
.Y(n_7069)
);

INVx5_ASAP7_75t_L g7070 ( 
.A(n_6480),
.Y(n_7070)
);

BUFx12f_ASAP7_75t_L g7071 ( 
.A(n_6208),
.Y(n_7071)
);

CKINVDCx11_ASAP7_75t_R g7072 ( 
.A(n_6208),
.Y(n_7072)
);

INVx1_ASAP7_75t_SL g7073 ( 
.A(n_5940),
.Y(n_7073)
);

CKINVDCx20_ASAP7_75t_R g7074 ( 
.A(n_6457),
.Y(n_7074)
);

OAI22xp5_ASAP7_75t_L g7075 ( 
.A1(n_6209),
.A2(n_5107),
.B1(n_5143),
.B2(n_5133),
.Y(n_7075)
);

CKINVDCx11_ASAP7_75t_R g7076 ( 
.A(n_6208),
.Y(n_7076)
);

CKINVDCx11_ASAP7_75t_R g7077 ( 
.A(n_6401),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_5922),
.Y(n_7078)
);

NAND2x1p5_ASAP7_75t_L g7079 ( 
.A(n_6321),
.B(n_5655),
.Y(n_7079)
);

OAI22xp33_ASAP7_75t_L g7080 ( 
.A1(n_5954),
.A2(n_5462),
.B1(n_5471),
.B2(n_5415),
.Y(n_7080)
);

AOI22xp33_ASAP7_75t_L g7081 ( 
.A1(n_6159),
.A2(n_5462),
.B1(n_5471),
.B2(n_5415),
.Y(n_7081)
);

CKINVDCx20_ASAP7_75t_R g7082 ( 
.A(n_6552),
.Y(n_7082)
);

INVx5_ASAP7_75t_L g7083 ( 
.A(n_6480),
.Y(n_7083)
);

INVx2_ASAP7_75t_L g7084 ( 
.A(n_5974),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_5922),
.Y(n_7085)
);

INVx3_ASAP7_75t_L g7086 ( 
.A(n_5835),
.Y(n_7086)
);

INVx3_ASAP7_75t_L g7087 ( 
.A(n_5835),
.Y(n_7087)
);

BUFx3_ASAP7_75t_L g7088 ( 
.A(n_6421),
.Y(n_7088)
);

AOI22xp33_ASAP7_75t_SL g7089 ( 
.A1(n_5787),
.A2(n_5166),
.B1(n_5472),
.B2(n_5349),
.Y(n_7089)
);

INVx6_ASAP7_75t_L g7090 ( 
.A(n_5899),
.Y(n_7090)
);

AOI22xp33_ASAP7_75t_L g7091 ( 
.A1(n_6159),
.A2(n_5471),
.B1(n_5462),
.B2(n_5151),
.Y(n_7091)
);

INVx4_ASAP7_75t_SL g7092 ( 
.A(n_6161),
.Y(n_7092)
);

BUFx6f_ASAP7_75t_L g7093 ( 
.A(n_6480),
.Y(n_7093)
);

INVx2_ASAP7_75t_L g7094 ( 
.A(n_5974),
.Y(n_7094)
);

BUFx12f_ASAP7_75t_L g7095 ( 
.A(n_6421),
.Y(n_7095)
);

INVx1_ASAP7_75t_SL g7096 ( 
.A(n_5940),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_5934),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_5934),
.Y(n_7098)
);

OAI22xp5_ASAP7_75t_L g7099 ( 
.A1(n_6209),
.A2(n_5107),
.B1(n_5143),
.B2(n_5133),
.Y(n_7099)
);

BUFx3_ASAP7_75t_L g7100 ( 
.A(n_6421),
.Y(n_7100)
);

AOI22xp33_ASAP7_75t_L g7101 ( 
.A1(n_6162),
.A2(n_5471),
.B1(n_5462),
.B2(n_5151),
.Y(n_7101)
);

CKINVDCx11_ASAP7_75t_R g7102 ( 
.A(n_6430),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_5941),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_5941),
.Y(n_7104)
);

AOI22xp5_ASAP7_75t_L g7105 ( 
.A1(n_6590),
.A2(n_5341),
.B1(n_5424),
.B2(n_5471),
.Y(n_7105)
);

CKINVDCx11_ASAP7_75t_R g7106 ( 
.A(n_6430),
.Y(n_7106)
);

CKINVDCx11_ASAP7_75t_R g7107 ( 
.A(n_6430),
.Y(n_7107)
);

BUFx2_ASAP7_75t_L g7108 ( 
.A(n_5923),
.Y(n_7108)
);

BUFx8_ASAP7_75t_L g7109 ( 
.A(n_6453),
.Y(n_7109)
);

AOI22xp33_ASAP7_75t_L g7110 ( 
.A1(n_6162),
.A2(n_5151),
.B1(n_5206),
.B2(n_5152),
.Y(n_7110)
);

CKINVDCx20_ASAP7_75t_R g7111 ( 
.A(n_6578),
.Y(n_7111)
);

INVx2_ASAP7_75t_L g7112 ( 
.A(n_5974),
.Y(n_7112)
);

BUFx4f_ASAP7_75t_SL g7113 ( 
.A(n_6453),
.Y(n_7113)
);

AOI22xp33_ASAP7_75t_L g7114 ( 
.A1(n_6404),
.A2(n_5151),
.B1(n_5206),
.B2(n_5152),
.Y(n_7114)
);

BUFx6f_ASAP7_75t_L g7115 ( 
.A(n_6480),
.Y(n_7115)
);

AOI22xp33_ASAP7_75t_L g7116 ( 
.A1(n_6404),
.A2(n_5151),
.B1(n_5206),
.B2(n_5152),
.Y(n_7116)
);

CKINVDCx11_ASAP7_75t_R g7117 ( 
.A(n_6453),
.Y(n_7117)
);

AOI22xp33_ASAP7_75t_L g7118 ( 
.A1(n_5889),
.A2(n_5152),
.B1(n_5206),
.B2(n_5472),
.Y(n_7118)
);

CKINVDCx11_ASAP7_75t_R g7119 ( 
.A(n_6274),
.Y(n_7119)
);

INVx3_ASAP7_75t_L g7120 ( 
.A(n_5835),
.Y(n_7120)
);

OAI21xp5_ASAP7_75t_SL g7121 ( 
.A1(n_6576),
.A2(n_5716),
.B(n_5483),
.Y(n_7121)
);

BUFx3_ASAP7_75t_L g7122 ( 
.A(n_6596),
.Y(n_7122)
);

OAI22xp5_ASAP7_75t_L g7123 ( 
.A1(n_6604),
.A2(n_5143),
.B1(n_5158),
.B2(n_5133),
.Y(n_7123)
);

OAI22xp33_ASAP7_75t_SL g7124 ( 
.A1(n_5889),
.A2(n_5701),
.B1(n_5283),
.B2(n_5324),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_5946),
.Y(n_7125)
);

OAI22xp5_ASAP7_75t_L g7126 ( 
.A1(n_6604),
.A2(n_5158),
.B1(n_5480),
.B2(n_5776),
.Y(n_7126)
);

INVx6_ASAP7_75t_L g7127 ( 
.A(n_5899),
.Y(n_7127)
);

INVx2_ASAP7_75t_SL g7128 ( 
.A(n_5812),
.Y(n_7128)
);

CKINVDCx5p33_ASAP7_75t_R g7129 ( 
.A(n_6603),
.Y(n_7129)
);

INVx4_ASAP7_75t_L g7130 ( 
.A(n_6611),
.Y(n_7130)
);

CKINVDCx11_ASAP7_75t_R g7131 ( 
.A(n_6274),
.Y(n_7131)
);

INVx2_ASAP7_75t_L g7132 ( 
.A(n_6081),
.Y(n_7132)
);

INVx1_ASAP7_75t_SL g7133 ( 
.A(n_5947),
.Y(n_7133)
);

BUFx12f_ASAP7_75t_L g7134 ( 
.A(n_6659),
.Y(n_7134)
);

BUFx3_ASAP7_75t_L g7135 ( 
.A(n_6611),
.Y(n_7135)
);

OAI21xp33_ASAP7_75t_L g7136 ( 
.A1(n_5895),
.A2(n_5410),
.B(n_5701),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_6081),
.Y(n_7137)
);

AOI22xp33_ASAP7_75t_L g7138 ( 
.A1(n_6621),
.A2(n_5152),
.B1(n_5206),
.B2(n_5536),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_5946),
.Y(n_7139)
);

BUFx10_ASAP7_75t_L g7140 ( 
.A(n_6143),
.Y(n_7140)
);

INVx4_ASAP7_75t_SL g7141 ( 
.A(n_6161),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6081),
.Y(n_7142)
);

INVx4_ASAP7_75t_L g7143 ( 
.A(n_6611),
.Y(n_7143)
);

INVx2_ASAP7_75t_L g7144 ( 
.A(n_6081),
.Y(n_7144)
);

OAI22xp33_ASAP7_75t_L g7145 ( 
.A1(n_5954),
.A2(n_5437),
.B1(n_5410),
.B2(n_5701),
.Y(n_7145)
);

NAND2xp5_ASAP7_75t_L g7146 ( 
.A(n_6416),
.B(n_5310),
.Y(n_7146)
);

BUFx3_ASAP7_75t_L g7147 ( 
.A(n_5877),
.Y(n_7147)
);

BUFx6f_ASAP7_75t_L g7148 ( 
.A(n_6518),
.Y(n_7148)
);

INVx5_ASAP7_75t_L g7149 ( 
.A(n_6518),
.Y(n_7149)
);

CKINVDCx6p67_ASAP7_75t_R g7150 ( 
.A(n_6274),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_6647),
.B(n_5573),
.Y(n_7151)
);

NAND2x1p5_ASAP7_75t_L g7152 ( 
.A(n_6321),
.B(n_5655),
.Y(n_7152)
);

AOI22xp33_ASAP7_75t_L g7153 ( 
.A1(n_6621),
.A2(n_5152),
.B1(n_5206),
.B2(n_5536),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_5948),
.Y(n_7154)
);

AOI22xp33_ASAP7_75t_L g7155 ( 
.A1(n_6215),
.A2(n_5152),
.B1(n_5206),
.B2(n_5536),
.Y(n_7155)
);

BUFx4f_ASAP7_75t_SL g7156 ( 
.A(n_6274),
.Y(n_7156)
);

BUFx2_ASAP7_75t_L g7157 ( 
.A(n_5923),
.Y(n_7157)
);

AOI21xp33_ASAP7_75t_L g7158 ( 
.A1(n_6068),
.A2(n_5481),
.B(n_5410),
.Y(n_7158)
);

AOI21xp33_ASAP7_75t_L g7159 ( 
.A1(n_6068),
.A2(n_5481),
.B(n_5682),
.Y(n_7159)
);

AOI22xp5_ASAP7_75t_SL g7160 ( 
.A1(n_6519),
.A2(n_5593),
.B1(n_5609),
.B2(n_5170),
.Y(n_7160)
);

AOI22xp33_ASAP7_75t_L g7161 ( 
.A1(n_6215),
.A2(n_5152),
.B1(n_5206),
.B2(n_5536),
.Y(n_7161)
);

AOI22xp33_ASAP7_75t_L g7162 ( 
.A1(n_6216),
.A2(n_5152),
.B1(n_5206),
.B2(n_5183),
.Y(n_7162)
);

INVx1_ASAP7_75t_SL g7163 ( 
.A(n_5947),
.Y(n_7163)
);

AOI22xp33_ASAP7_75t_L g7164 ( 
.A1(n_6216),
.A2(n_5907),
.B1(n_5890),
.B2(n_6629),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_5948),
.Y(n_7165)
);

INVx2_ASAP7_75t_L g7166 ( 
.A(n_6081),
.Y(n_7166)
);

AOI22xp33_ASAP7_75t_L g7167 ( 
.A1(n_5907),
.A2(n_5152),
.B1(n_5206),
.B2(n_5183),
.Y(n_7167)
);

BUFx6f_ASAP7_75t_L g7168 ( 
.A(n_6518),
.Y(n_7168)
);

INVx2_ASAP7_75t_L g7169 ( 
.A(n_6181),
.Y(n_7169)
);

AOI22xp33_ASAP7_75t_L g7170 ( 
.A1(n_5890),
.A2(n_5105),
.B1(n_5096),
.B2(n_5102),
.Y(n_7170)
);

CKINVDCx20_ASAP7_75t_R g7171 ( 
.A(n_6341),
.Y(n_7171)
);

CKINVDCx20_ASAP7_75t_R g7172 ( 
.A(n_6341),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_5949),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_5949),
.Y(n_7174)
);

AOI22xp5_ASAP7_75t_L g7175 ( 
.A1(n_6349),
.A2(n_6446),
.B1(n_6477),
.B2(n_5859),
.Y(n_7175)
);

AOI22xp5_ASAP7_75t_L g7176 ( 
.A1(n_6349),
.A2(n_5422),
.B1(n_5416),
.B2(n_5170),
.Y(n_7176)
);

OAI22xp5_ASAP7_75t_L g7177 ( 
.A1(n_5895),
.A2(n_5898),
.B1(n_6474),
.B2(n_6452),
.Y(n_7177)
);

INVx2_ASAP7_75t_L g7178 ( 
.A(n_6181),
.Y(n_7178)
);

AOI22xp33_ASAP7_75t_L g7179 ( 
.A1(n_6629),
.A2(n_5105),
.B1(n_5096),
.B2(n_5102),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_5980),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_5980),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6181),
.Y(n_7182)
);

CKINVDCx6p67_ASAP7_75t_R g7183 ( 
.A(n_6335),
.Y(n_7183)
);

INVx3_ASAP7_75t_L g7184 ( 
.A(n_5835),
.Y(n_7184)
);

BUFx6f_ASAP7_75t_L g7185 ( 
.A(n_6518),
.Y(n_7185)
);

AOI22xp33_ASAP7_75t_SL g7186 ( 
.A1(n_6519),
.A2(n_5166),
.B1(n_5481),
.B2(n_5158),
.Y(n_7186)
);

CKINVDCx5p33_ASAP7_75t_R g7187 ( 
.A(n_6291),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_5982),
.Y(n_7188)
);

OAI22xp5_ASAP7_75t_L g7189 ( 
.A1(n_5898),
.A2(n_5776),
.B1(n_5766),
.B2(n_5683),
.Y(n_7189)
);

INVxp67_ASAP7_75t_SL g7190 ( 
.A(n_6036),
.Y(n_7190)
);

AOI22xp33_ASAP7_75t_L g7191 ( 
.A1(n_6089),
.A2(n_5169),
.B1(n_5105),
.B2(n_5096),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_5982),
.Y(n_7192)
);

AOI21xp5_ASAP7_75t_L g7193 ( 
.A1(n_5872),
.A2(n_5689),
.B(n_5283),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_5991),
.Y(n_7194)
);

AOI22xp33_ASAP7_75t_SL g7195 ( 
.A1(n_6556),
.A2(n_6160),
.B1(n_6276),
.B2(n_5975),
.Y(n_7195)
);

INVx1_ASAP7_75t_SL g7196 ( 
.A(n_5952),
.Y(n_7196)
);

BUFx12f_ASAP7_75t_L g7197 ( 
.A(n_6504),
.Y(n_7197)
);

INVx2_ASAP7_75t_L g7198 ( 
.A(n_6181),
.Y(n_7198)
);

CKINVDCx20_ASAP7_75t_R g7199 ( 
.A(n_6341),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_6526),
.B(n_5310),
.Y(n_7200)
);

OAI22xp5_ASAP7_75t_L g7201 ( 
.A1(n_6452),
.A2(n_5766),
.B1(n_5683),
.B2(n_5694),
.Y(n_7201)
);

AOI22xp33_ASAP7_75t_SL g7202 ( 
.A1(n_6556),
.A2(n_5481),
.B1(n_5245),
.B2(n_5559),
.Y(n_7202)
);

INVx6_ASAP7_75t_L g7203 ( 
.A(n_5899),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_5991),
.Y(n_7204)
);

AOI22xp33_ASAP7_75t_SL g7205 ( 
.A1(n_6160),
.A2(n_5481),
.B1(n_5245),
.B2(n_5689),
.Y(n_7205)
);

AOI22xp33_ASAP7_75t_L g7206 ( 
.A1(n_6089),
.A2(n_6240),
.B1(n_6252),
.B2(n_6016),
.Y(n_7206)
);

CKINVDCx16_ASAP7_75t_R g7207 ( 
.A(n_6346),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_5995),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_5995),
.Y(n_7209)
);

BUFx3_ASAP7_75t_L g7210 ( 
.A(n_6072),
.Y(n_7210)
);

OAI21xp5_ASAP7_75t_SL g7211 ( 
.A1(n_6576),
.A2(n_5259),
.B(n_5371),
.Y(n_7211)
);

INVx2_ASAP7_75t_L g7212 ( 
.A(n_6181),
.Y(n_7212)
);

BUFx2_ASAP7_75t_SL g7213 ( 
.A(n_6268),
.Y(n_7213)
);

AOI22xp33_ASAP7_75t_L g7214 ( 
.A1(n_6240),
.A2(n_5169),
.B1(n_5105),
.B2(n_5096),
.Y(n_7214)
);

CKINVDCx20_ASAP7_75t_R g7215 ( 
.A(n_6335),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_6206),
.Y(n_7216)
);

INVx3_ASAP7_75t_SL g7217 ( 
.A(n_6348),
.Y(n_7217)
);

INVx2_ASAP7_75t_L g7218 ( 
.A(n_6206),
.Y(n_7218)
);

CKINVDCx6p67_ASAP7_75t_R g7219 ( 
.A(n_6335),
.Y(n_7219)
);

OAI21xp5_ASAP7_75t_L g7220 ( 
.A1(n_5881),
.A2(n_5523),
.B(n_5281),
.Y(n_7220)
);

INVx6_ASAP7_75t_L g7221 ( 
.A(n_5899),
.Y(n_7221)
);

AOI22xp33_ASAP7_75t_SL g7222 ( 
.A1(n_6276),
.A2(n_5481),
.B1(n_5245),
.B2(n_5715),
.Y(n_7222)
);

AOI22xp33_ASAP7_75t_L g7223 ( 
.A1(n_6252),
.A2(n_5235),
.B1(n_5219),
.B2(n_5096),
.Y(n_7223)
);

INVx2_ASAP7_75t_L g7224 ( 
.A(n_6206),
.Y(n_7224)
);

BUFx6f_ASAP7_75t_L g7225 ( 
.A(n_6518),
.Y(n_7225)
);

AOI22xp33_ASAP7_75t_L g7226 ( 
.A1(n_6016),
.A2(n_6446),
.B1(n_6477),
.B2(n_6084),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_5999),
.Y(n_7227)
);

INVx2_ASAP7_75t_SL g7228 ( 
.A(n_5812),
.Y(n_7228)
);

BUFx2_ASAP7_75t_SL g7229 ( 
.A(n_6268),
.Y(n_7229)
);

INVx4_ASAP7_75t_L g7230 ( 
.A(n_6170),
.Y(n_7230)
);

CKINVDCx20_ASAP7_75t_R g7231 ( 
.A(n_6335),
.Y(n_7231)
);

INVx2_ASAP7_75t_L g7232 ( 
.A(n_6206),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_5999),
.Y(n_7233)
);

INVx8_ASAP7_75t_L g7234 ( 
.A(n_6161),
.Y(n_7234)
);

OAI22x1_ASAP7_75t_SL g7235 ( 
.A1(n_5805),
.A2(n_5675),
.B1(n_5651),
.B2(n_5508),
.Y(n_7235)
);

OAI22xp33_ASAP7_75t_L g7236 ( 
.A1(n_6153),
.A2(n_5437),
.B1(n_5332),
.B2(n_5430),
.Y(n_7236)
);

CKINVDCx11_ASAP7_75t_R g7237 ( 
.A(n_6601),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_L g7238 ( 
.A(n_6526),
.B(n_5323),
.Y(n_7238)
);

INVx1_ASAP7_75t_SL g7239 ( 
.A(n_5952),
.Y(n_7239)
);

INVx4_ASAP7_75t_L g7240 ( 
.A(n_6170),
.Y(n_7240)
);

INVx2_ASAP7_75t_L g7241 ( 
.A(n_6206),
.Y(n_7241)
);

CKINVDCx20_ASAP7_75t_R g7242 ( 
.A(n_6601),
.Y(n_7242)
);

AOI22xp33_ASAP7_75t_SL g7243 ( 
.A1(n_5975),
.A2(n_5715),
.B1(n_5752),
.B2(n_5727),
.Y(n_7243)
);

CKINVDCx6p67_ASAP7_75t_R g7244 ( 
.A(n_6601),
.Y(n_7244)
);

BUFx12f_ASAP7_75t_L g7245 ( 
.A(n_6504),
.Y(n_7245)
);

OAI21xp5_ASAP7_75t_SL g7246 ( 
.A1(n_6650),
.A2(n_5259),
.B(n_5371),
.Y(n_7246)
);

INVx2_ASAP7_75t_SL g7247 ( 
.A(n_5812),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_6001),
.Y(n_7248)
);

CKINVDCx16_ASAP7_75t_R g7249 ( 
.A(n_6346),
.Y(n_7249)
);

CKINVDCx11_ASAP7_75t_R g7250 ( 
.A(n_6601),
.Y(n_7250)
);

BUFx3_ASAP7_75t_L g7251 ( 
.A(n_6072),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6001),
.Y(n_7252)
);

INVx3_ASAP7_75t_L g7253 ( 
.A(n_6589),
.Y(n_7253)
);

INVx2_ASAP7_75t_SL g7254 ( 
.A(n_5887),
.Y(n_7254)
);

INVx2_ASAP7_75t_L g7255 ( 
.A(n_6222),
.Y(n_7255)
);

CKINVDCx5p33_ASAP7_75t_R g7256 ( 
.A(n_6291),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_6008),
.Y(n_7257)
);

AOI22xp33_ASAP7_75t_L g7258 ( 
.A1(n_6084),
.A2(n_5235),
.B1(n_5219),
.B2(n_5096),
.Y(n_7258)
);

AOI22xp33_ASAP7_75t_SL g7259 ( 
.A1(n_6669),
.A2(n_5715),
.B1(n_5752),
.B2(n_5727),
.Y(n_7259)
);

OAI22xp5_ASAP7_75t_L g7260 ( 
.A1(n_6452),
.A2(n_5674),
.B1(n_5698),
.B2(n_5694),
.Y(n_7260)
);

INVx2_ASAP7_75t_L g7261 ( 
.A(n_6222),
.Y(n_7261)
);

CKINVDCx11_ASAP7_75t_R g7262 ( 
.A(n_6516),
.Y(n_7262)
);

INVx2_ASAP7_75t_SL g7263 ( 
.A(n_5887),
.Y(n_7263)
);

OAI22xp5_ASAP7_75t_L g7264 ( 
.A1(n_6474),
.A2(n_6153),
.B1(n_5902),
.B2(n_6019),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_6008),
.Y(n_7265)
);

INVx1_ASAP7_75t_SL g7266 ( 
.A(n_6412),
.Y(n_7266)
);

AOI22xp33_ASAP7_75t_L g7267 ( 
.A1(n_6084),
.A2(n_5102),
.B1(n_5169),
.B2(n_5118),
.Y(n_7267)
);

OAI21xp5_ASAP7_75t_L g7268 ( 
.A1(n_5881),
.A2(n_5523),
.B(n_5281),
.Y(n_7268)
);

OAI22xp33_ASAP7_75t_L g7269 ( 
.A1(n_6019),
.A2(n_5437),
.B1(n_5430),
.B2(n_5332),
.Y(n_7269)
);

INVx6_ASAP7_75t_L g7270 ( 
.A(n_5899),
.Y(n_7270)
);

OAI21xp5_ASAP7_75t_SL g7271 ( 
.A1(n_6650),
.A2(n_5259),
.B(n_5371),
.Y(n_7271)
);

BUFx12f_ASAP7_75t_L g7272 ( 
.A(n_6516),
.Y(n_7272)
);

CKINVDCx11_ASAP7_75t_R g7273 ( 
.A(n_6538),
.Y(n_7273)
);

AOI22xp33_ASAP7_75t_SL g7274 ( 
.A1(n_6669),
.A2(n_5727),
.B1(n_5752),
.B2(n_5740),
.Y(n_7274)
);

BUFx2_ASAP7_75t_L g7275 ( 
.A(n_5923),
.Y(n_7275)
);

BUFx12f_ASAP7_75t_L g7276 ( 
.A(n_6538),
.Y(n_7276)
);

BUFx2_ASAP7_75t_SL g7277 ( 
.A(n_6646),
.Y(n_7277)
);

INVx4_ASAP7_75t_L g7278 ( 
.A(n_6170),
.Y(n_7278)
);

AOI22xp33_ASAP7_75t_L g7279 ( 
.A1(n_6084),
.A2(n_5102),
.B1(n_5169),
.B2(n_5118),
.Y(n_7279)
);

CKINVDCx20_ASAP7_75t_R g7280 ( 
.A(n_6297),
.Y(n_7280)
);

CKINVDCx5p33_ASAP7_75t_R g7281 ( 
.A(n_6297),
.Y(n_7281)
);

AOI22xp33_ASAP7_75t_SL g7282 ( 
.A1(n_6673),
.A2(n_5371),
.B1(n_5283),
.B2(n_5324),
.Y(n_7282)
);

OAI22xp33_ASAP7_75t_L g7283 ( 
.A1(n_5859),
.A2(n_5437),
.B1(n_5430),
.B2(n_5332),
.Y(n_7283)
);

INVx5_ASAP7_75t_L g7284 ( 
.A(n_6518),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6010),
.Y(n_7285)
);

NOR2xp33_ASAP7_75t_L g7286 ( 
.A(n_6557),
.B(n_5651),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_6517),
.B(n_5323),
.Y(n_7287)
);

OAI21xp5_ASAP7_75t_L g7288 ( 
.A1(n_5912),
.A2(n_5281),
.B(n_5280),
.Y(n_7288)
);

BUFx8_ASAP7_75t_L g7289 ( 
.A(n_6503),
.Y(n_7289)
);

OAI22xp33_ASAP7_75t_L g7290 ( 
.A1(n_6099),
.A2(n_5437),
.B1(n_5430),
.B2(n_5093),
.Y(n_7290)
);

OAI22xp33_ASAP7_75t_L g7291 ( 
.A1(n_6099),
.A2(n_5093),
.B1(n_5621),
.B2(n_5535),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_6222),
.Y(n_7292)
);

OAI22xp5_ASAP7_75t_L g7293 ( 
.A1(n_6474),
.A2(n_5674),
.B1(n_5706),
.B2(n_5698),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_6010),
.Y(n_7294)
);

INVx8_ASAP7_75t_L g7295 ( 
.A(n_6161),
.Y(n_7295)
);

AOI22xp33_ASAP7_75t_L g7296 ( 
.A1(n_6084),
.A2(n_5102),
.B1(n_5169),
.B2(n_5118),
.Y(n_7296)
);

NAND2x1p5_ASAP7_75t_L g7297 ( 
.A(n_6321),
.B(n_5655),
.Y(n_7297)
);

CKINVDCx11_ASAP7_75t_R g7298 ( 
.A(n_6668),
.Y(n_7298)
);

AOI22xp33_ASAP7_75t_L g7299 ( 
.A1(n_6084),
.A2(n_5102),
.B1(n_5169),
.B2(n_5118),
.Y(n_7299)
);

INVx6_ASAP7_75t_L g7300 ( 
.A(n_6454),
.Y(n_7300)
);

CKINVDCx16_ASAP7_75t_R g7301 ( 
.A(n_6156),
.Y(n_7301)
);

AND2x2_ASAP7_75t_L g7302 ( 
.A(n_6018),
.B(n_5537),
.Y(n_7302)
);

BUFx8_ASAP7_75t_L g7303 ( 
.A(n_6503),
.Y(n_7303)
);

BUFx2_ASAP7_75t_L g7304 ( 
.A(n_6595),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_6023),
.Y(n_7305)
);

OAI22xp33_ASAP7_75t_L g7306 ( 
.A1(n_6128),
.A2(n_5093),
.B1(n_5621),
.B2(n_5535),
.Y(n_7306)
);

OAI22xp33_ASAP7_75t_L g7307 ( 
.A1(n_6128),
.A2(n_5093),
.B1(n_5621),
.B2(n_5535),
.Y(n_7307)
);

INVx2_ASAP7_75t_L g7308 ( 
.A(n_6222),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_6023),
.Y(n_7309)
);

OAI22xp33_ASAP7_75t_L g7310 ( 
.A1(n_6113),
.A2(n_5535),
.B1(n_5621),
.B2(n_5283),
.Y(n_7310)
);

AOI22xp33_ASAP7_75t_L g7311 ( 
.A1(n_6084),
.A2(n_5183),
.B1(n_5219),
.B2(n_5118),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_6030),
.Y(n_7312)
);

BUFx8_ASAP7_75t_SL g7313 ( 
.A(n_6102),
.Y(n_7313)
);

AOI22xp33_ASAP7_75t_L g7314 ( 
.A1(n_6084),
.A2(n_5183),
.B1(n_5235),
.B2(n_5219),
.Y(n_7314)
);

AOI22xp33_ASAP7_75t_L g7315 ( 
.A1(n_6084),
.A2(n_5183),
.B1(n_5235),
.B2(n_5219),
.Y(n_7315)
);

OR2x2_ASAP7_75t_L g7316 ( 
.A(n_5930),
.B(n_5744),
.Y(n_7316)
);

AOI22xp33_ASAP7_75t_L g7317 ( 
.A1(n_6084),
.A2(n_5183),
.B1(n_5235),
.B2(n_5219),
.Y(n_7317)
);

INVx2_ASAP7_75t_L g7318 ( 
.A(n_6222),
.Y(n_7318)
);

INVx6_ASAP7_75t_L g7319 ( 
.A(n_6454),
.Y(n_7319)
);

AOI22xp33_ASAP7_75t_SL g7320 ( 
.A1(n_6673),
.A2(n_6113),
.B1(n_6584),
.B2(n_6571),
.Y(n_7320)
);

OAI22xp5_ASAP7_75t_L g7321 ( 
.A1(n_5902),
.A2(n_5722),
.B1(n_5759),
.B2(n_5706),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_6030),
.Y(n_7322)
);

AOI22xp33_ASAP7_75t_SL g7323 ( 
.A1(n_6571),
.A2(n_5283),
.B1(n_5324),
.B2(n_5170),
.Y(n_7323)
);

AND2x2_ASAP7_75t_L g7324 ( 
.A(n_6018),
.B(n_5537),
.Y(n_7324)
);

NAND2x1p5_ASAP7_75t_L g7325 ( 
.A(n_6324),
.B(n_5100),
.Y(n_7325)
);

OAI22xp5_ASAP7_75t_SL g7326 ( 
.A1(n_5929),
.A2(n_5675),
.B1(n_5759),
.B2(n_5722),
.Y(n_7326)
);

INVxp67_ASAP7_75t_SL g7327 ( 
.A(n_6036),
.Y(n_7327)
);

OAI22xp5_ASAP7_75t_L g7328 ( 
.A1(n_6009),
.A2(n_5112),
.B1(n_5305),
.B2(n_5284),
.Y(n_7328)
);

BUFx5_ASAP7_75t_L g7329 ( 
.A(n_6004),
.Y(n_7329)
);

CKINVDCx11_ASAP7_75t_R g7330 ( 
.A(n_6668),
.Y(n_7330)
);

CKINVDCx6p67_ASAP7_75t_R g7331 ( 
.A(n_6668),
.Y(n_7331)
);

AOI22xp33_ASAP7_75t_L g7332 ( 
.A1(n_6557),
.A2(n_5235),
.B1(n_5221),
.B2(n_5116),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6034),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_6034),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_6037),
.Y(n_7335)
);

AOI22xp33_ASAP7_75t_L g7336 ( 
.A1(n_6591),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7336)
);

OAI22xp33_ASAP7_75t_L g7337 ( 
.A1(n_6397),
.A2(n_5283),
.B1(n_5422),
.B2(n_5416),
.Y(n_7337)
);

BUFx10_ASAP7_75t_L g7338 ( 
.A(n_6518),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_6037),
.Y(n_7339)
);

CKINVDCx5p33_ASAP7_75t_R g7340 ( 
.A(n_6591),
.Y(n_7340)
);

INVx4_ASAP7_75t_L g7341 ( 
.A(n_6665),
.Y(n_7341)
);

AND2x2_ASAP7_75t_L g7342 ( 
.A(n_6018),
.B(n_5537),
.Y(n_7342)
);

BUFx10_ASAP7_75t_L g7343 ( 
.A(n_6518),
.Y(n_7343)
);

INVx2_ASAP7_75t_L g7344 ( 
.A(n_5794),
.Y(n_7344)
);

INVx4_ASAP7_75t_L g7345 ( 
.A(n_5805),
.Y(n_7345)
);

INVx2_ASAP7_75t_SL g7346 ( 
.A(n_5887),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_6042),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_6042),
.Y(n_7348)
);

OAI21xp5_ASAP7_75t_SL g7349 ( 
.A1(n_6645),
.A2(n_5259),
.B(n_5150),
.Y(n_7349)
);

AOI22xp33_ASAP7_75t_L g7350 ( 
.A1(n_6237),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_6043),
.Y(n_7351)
);

OAI22xp5_ASAP7_75t_L g7352 ( 
.A1(n_6009),
.A2(n_5112),
.B1(n_5305),
.B2(n_5284),
.Y(n_7352)
);

BUFx3_ASAP7_75t_L g7353 ( 
.A(n_6072),
.Y(n_7353)
);

AOI22xp33_ASAP7_75t_L g7354 ( 
.A1(n_6237),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7354)
);

AOI21xp33_ASAP7_75t_L g7355 ( 
.A1(n_6497),
.A2(n_5682),
.B(n_5283),
.Y(n_7355)
);

INVx1_ASAP7_75t_SL g7356 ( 
.A(n_6412),
.Y(n_7356)
);

AOI22xp33_ASAP7_75t_L g7357 ( 
.A1(n_6238),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7357)
);

CKINVDCx11_ASAP7_75t_R g7358 ( 
.A(n_6668),
.Y(n_7358)
);

INVx2_ASAP7_75t_L g7359 ( 
.A(n_5794),
.Y(n_7359)
);

AOI22xp33_ASAP7_75t_L g7360 ( 
.A1(n_6238),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7360)
);

OAI22xp5_ASAP7_75t_L g7361 ( 
.A1(n_6428),
.A2(n_5112),
.B1(n_5305),
.B2(n_5284),
.Y(n_7361)
);

BUFx6f_ASAP7_75t_L g7362 ( 
.A(n_6521),
.Y(n_7362)
);

AOI22xp33_ASAP7_75t_L g7363 ( 
.A1(n_6529),
.A2(n_5191),
.B1(n_5192),
.B2(n_5179),
.Y(n_7363)
);

INVx4_ASAP7_75t_L g7364 ( 
.A(n_6665),
.Y(n_7364)
);

INVx6_ASAP7_75t_L g7365 ( 
.A(n_6454),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_5794),
.Y(n_7366)
);

CKINVDCx11_ASAP7_75t_R g7367 ( 
.A(n_6102),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_6043),
.Y(n_7368)
);

CKINVDCx20_ASAP7_75t_R g7369 ( 
.A(n_6102),
.Y(n_7369)
);

BUFx6f_ASAP7_75t_L g7370 ( 
.A(n_6521),
.Y(n_7370)
);

AOI22xp33_ASAP7_75t_L g7371 ( 
.A1(n_6529),
.A2(n_5192),
.B1(n_5593),
.B2(n_5170),
.Y(n_7371)
);

INVx1_ASAP7_75t_SL g7372 ( 
.A(n_6412),
.Y(n_7372)
);

INVx6_ASAP7_75t_L g7373 ( 
.A(n_6454),
.Y(n_7373)
);

INVx6_ASAP7_75t_L g7374 ( 
.A(n_6454),
.Y(n_7374)
);

BUFx12f_ASAP7_75t_L g7375 ( 
.A(n_5805),
.Y(n_7375)
);

NAND2x1p5_ASAP7_75t_L g7376 ( 
.A(n_6324),
.B(n_5100),
.Y(n_7376)
);

AOI22xp33_ASAP7_75t_L g7377 ( 
.A1(n_6375),
.A2(n_5170),
.B1(n_5609),
.B2(n_5593),
.Y(n_7377)
);

CKINVDCx20_ASAP7_75t_R g7378 ( 
.A(n_6102),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_6069),
.Y(n_7379)
);

OAI22xp5_ASAP7_75t_L g7380 ( 
.A1(n_6428),
.A2(n_5112),
.B1(n_5305),
.B2(n_5284),
.Y(n_7380)
);

BUFx3_ASAP7_75t_L g7381 ( 
.A(n_6072),
.Y(n_7381)
);

AOI22xp33_ASAP7_75t_L g7382 ( 
.A1(n_6375),
.A2(n_5170),
.B1(n_5609),
.B2(n_5593),
.Y(n_7382)
);

BUFx12f_ASAP7_75t_L g7383 ( 
.A(n_5805),
.Y(n_7383)
);

AOI22xp33_ASAP7_75t_L g7384 ( 
.A1(n_6451),
.A2(n_5170),
.B1(n_5609),
.B2(n_5593),
.Y(n_7384)
);

BUFx3_ASAP7_75t_L g7385 ( 
.A(n_6072),
.Y(n_7385)
);

INVx2_ASAP7_75t_SL g7386 ( 
.A(n_5887),
.Y(n_7386)
);

INVx4_ASAP7_75t_L g7387 ( 
.A(n_6665),
.Y(n_7387)
);

OAI22xp33_ASAP7_75t_L g7388 ( 
.A1(n_6397),
.A2(n_5283),
.B1(n_5422),
.B2(n_5416),
.Y(n_7388)
);

OAI22xp33_ASAP7_75t_L g7389 ( 
.A1(n_6156),
.A2(n_5324),
.B1(n_5539),
.B2(n_5756),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_6069),
.Y(n_7390)
);

OAI21xp5_ASAP7_75t_L g7391 ( 
.A1(n_6497),
.A2(n_5280),
.B(n_5682),
.Y(n_7391)
);

OAI22xp5_ASAP7_75t_L g7392 ( 
.A1(n_6308),
.A2(n_5348),
.B1(n_5265),
.B2(n_5587),
.Y(n_7392)
);

BUFx2_ASAP7_75t_L g7393 ( 
.A(n_6595),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_6074),
.Y(n_7394)
);

CKINVDCx11_ASAP7_75t_R g7395 ( 
.A(n_6169),
.Y(n_7395)
);

AOI22xp33_ASAP7_75t_L g7396 ( 
.A1(n_6451),
.A2(n_5170),
.B1(n_5609),
.B2(n_5593),
.Y(n_7396)
);

INVx1_ASAP7_75t_L g7397 ( 
.A(n_6074),
.Y(n_7397)
);

INVx3_ASAP7_75t_L g7398 ( 
.A(n_6589),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_5794),
.Y(n_7399)
);

AOI22xp33_ASAP7_75t_L g7400 ( 
.A1(n_6278),
.A2(n_5609),
.B1(n_5679),
.B2(n_5593),
.Y(n_7400)
);

AOI21xp5_ASAP7_75t_L g7401 ( 
.A1(n_5872),
.A2(n_5324),
.B(n_5659),
.Y(n_7401)
);

BUFx2_ASAP7_75t_L g7402 ( 
.A(n_6595),
.Y(n_7402)
);

INVx2_ASAP7_75t_L g7403 ( 
.A(n_5796),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_6090),
.Y(n_7404)
);

BUFx3_ASAP7_75t_L g7405 ( 
.A(n_6072),
.Y(n_7405)
);

BUFx2_ASAP7_75t_SL g7406 ( 
.A(n_6646),
.Y(n_7406)
);

AOI22xp33_ASAP7_75t_SL g7407 ( 
.A1(n_6584),
.A2(n_5324),
.B1(n_5609),
.B2(n_5593),
.Y(n_7407)
);

AOI22xp33_ASAP7_75t_L g7408 ( 
.A1(n_6278),
.A2(n_5609),
.B1(n_5679),
.B2(n_5593),
.Y(n_7408)
);

AOI22xp33_ASAP7_75t_L g7409 ( 
.A1(n_6038),
.A2(n_5609),
.B1(n_5679),
.B2(n_5593),
.Y(n_7409)
);

CKINVDCx6p67_ASAP7_75t_R g7410 ( 
.A(n_6169),
.Y(n_7410)
);

BUFx4_ASAP7_75t_R g7411 ( 
.A(n_5984),
.Y(n_7411)
);

CKINVDCx11_ASAP7_75t_R g7412 ( 
.A(n_6169),
.Y(n_7412)
);

CKINVDCx5p33_ASAP7_75t_R g7413 ( 
.A(n_6662),
.Y(n_7413)
);

AOI22xp5_ASAP7_75t_L g7414 ( 
.A1(n_5801),
.A2(n_5609),
.B1(n_5679),
.B2(n_5593),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_6090),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_6095),
.Y(n_7416)
);

AOI22xp33_ASAP7_75t_L g7417 ( 
.A1(n_6038),
.A2(n_5609),
.B1(n_5679),
.B2(n_5593),
.Y(n_7417)
);

AND2x4_ASAP7_75t_L g7418 ( 
.A(n_6132),
.B(n_5292),
.Y(n_7418)
);

INVx2_ASAP7_75t_L g7419 ( 
.A(n_5796),
.Y(n_7419)
);

INVx2_ASAP7_75t_SL g7420 ( 
.A(n_5887),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_6095),
.Y(n_7421)
);

AND2x2_ASAP7_75t_L g7422 ( 
.A(n_6544),
.B(n_5537),
.Y(n_7422)
);

HB1xp67_ASAP7_75t_L g7423 ( 
.A(n_6137),
.Y(n_7423)
);

CKINVDCx11_ASAP7_75t_R g7424 ( 
.A(n_6169),
.Y(n_7424)
);

INVx2_ASAP7_75t_L g7425 ( 
.A(n_5796),
.Y(n_7425)
);

AOI22xp33_ASAP7_75t_SL g7426 ( 
.A1(n_5857),
.A2(n_5324),
.B1(n_5679),
.B2(n_5609),
.Y(n_7426)
);

CKINVDCx20_ASAP7_75t_R g7427 ( 
.A(n_6245),
.Y(n_7427)
);

AND2x2_ASAP7_75t_L g7428 ( 
.A(n_6544),
.B(n_5543),
.Y(n_7428)
);

OAI22xp33_ASAP7_75t_L g7429 ( 
.A1(n_6330),
.A2(n_5324),
.B1(n_5539),
.B2(n_5756),
.Y(n_7429)
);

AOI22xp33_ASAP7_75t_L g7430 ( 
.A1(n_5857),
.A2(n_5697),
.B1(n_5679),
.B2(n_5258),
.Y(n_7430)
);

INVx8_ASAP7_75t_L g7431 ( 
.A(n_6161),
.Y(n_7431)
);

INVx3_ASAP7_75t_L g7432 ( 
.A(n_6589),
.Y(n_7432)
);

BUFx4_ASAP7_75t_SL g7433 ( 
.A(n_6245),
.Y(n_7433)
);

INVx6_ASAP7_75t_L g7434 ( 
.A(n_6524),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_6112),
.Y(n_7435)
);

BUFx12f_ASAP7_75t_L g7436 ( 
.A(n_5805),
.Y(n_7436)
);

AOI22xp33_ASAP7_75t_L g7437 ( 
.A1(n_6048),
.A2(n_5697),
.B1(n_5679),
.B2(n_5258),
.Y(n_7437)
);

INVx5_ASAP7_75t_L g7438 ( 
.A(n_6521),
.Y(n_7438)
);

AOI22xp33_ASAP7_75t_L g7439 ( 
.A1(n_6048),
.A2(n_5697),
.B1(n_5679),
.B2(n_5258),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6112),
.Y(n_7440)
);

INVx2_ASAP7_75t_L g7441 ( 
.A(n_5796),
.Y(n_7441)
);

BUFx12f_ASAP7_75t_L g7442 ( 
.A(n_5848),
.Y(n_7442)
);

NAND2xp5_ASAP7_75t_L g7443 ( 
.A(n_6517),
.B(n_5323),
.Y(n_7443)
);

BUFx6f_ASAP7_75t_L g7444 ( 
.A(n_6521),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_6114),
.Y(n_7445)
);

AOI22xp33_ASAP7_75t_L g7446 ( 
.A1(n_6640),
.A2(n_6660),
.B1(n_6658),
.B2(n_5891),
.Y(n_7446)
);

HB1xp67_ASAP7_75t_L g7447 ( 
.A(n_6137),
.Y(n_7447)
);

INVx3_ASAP7_75t_L g7448 ( 
.A(n_6589),
.Y(n_7448)
);

BUFx2_ASAP7_75t_L g7449 ( 
.A(n_6595),
.Y(n_7449)
);

INVx1_ASAP7_75t_SL g7450 ( 
.A(n_5967),
.Y(n_7450)
);

AND2x2_ASAP7_75t_L g7451 ( 
.A(n_6544),
.B(n_5543),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_6114),
.Y(n_7452)
);

OAI22xp5_ASAP7_75t_L g7453 ( 
.A1(n_6308),
.A2(n_5348),
.B1(n_5265),
.B2(n_5587),
.Y(n_7453)
);

AOI22xp33_ASAP7_75t_SL g7454 ( 
.A1(n_6012),
.A2(n_5697),
.B1(n_5679),
.B2(n_5372),
.Y(n_7454)
);

BUFx2_ASAP7_75t_L g7455 ( 
.A(n_6595),
.Y(n_7455)
);

INVx6_ASAP7_75t_L g7456 ( 
.A(n_6524),
.Y(n_7456)
);

AOI22xp33_ASAP7_75t_L g7457 ( 
.A1(n_6640),
.A2(n_5697),
.B1(n_5679),
.B2(n_5258),
.Y(n_7457)
);

INVx1_ASAP7_75t_SL g7458 ( 
.A(n_5967),
.Y(n_7458)
);

BUFx4f_ASAP7_75t_SL g7459 ( 
.A(n_6245),
.Y(n_7459)
);

INVx2_ASAP7_75t_L g7460 ( 
.A(n_5808),
.Y(n_7460)
);

BUFx12f_ASAP7_75t_L g7461 ( 
.A(n_5848),
.Y(n_7461)
);

OAI22xp5_ASAP7_75t_L g7462 ( 
.A1(n_6310),
.A2(n_5348),
.B1(n_5265),
.B2(n_5587),
.Y(n_7462)
);

INVx3_ASAP7_75t_L g7463 ( 
.A(n_6598),
.Y(n_7463)
);

BUFx2_ASAP7_75t_SL g7464 ( 
.A(n_6521),
.Y(n_7464)
);

AND2x4_ASAP7_75t_L g7465 ( 
.A(n_6132),
.B(n_5292),
.Y(n_7465)
);

BUFx8_ASAP7_75t_L g7466 ( 
.A(n_6503),
.Y(n_7466)
);

BUFx2_ASAP7_75t_R g7467 ( 
.A(n_6245),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6138),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_6138),
.Y(n_7469)
);

INVx3_ASAP7_75t_L g7470 ( 
.A(n_6598),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_6141),
.Y(n_7471)
);

OAI22xp5_ASAP7_75t_L g7472 ( 
.A1(n_6310),
.A2(n_6207),
.B1(n_6135),
.B2(n_6040),
.Y(n_7472)
);

INVx1_ASAP7_75t_L g7473 ( 
.A(n_6141),
.Y(n_7473)
);

CKINVDCx6p67_ASAP7_75t_R g7474 ( 
.A(n_6247),
.Y(n_7474)
);

OAI22xp33_ASAP7_75t_L g7475 ( 
.A1(n_6330),
.A2(n_5539),
.B1(n_5381),
.B2(n_5384),
.Y(n_7475)
);

OAI22xp5_ASAP7_75t_SL g7476 ( 
.A1(n_6666),
.A2(n_5539),
.B1(n_5372),
.B2(n_5384),
.Y(n_7476)
);

INVx3_ASAP7_75t_L g7477 ( 
.A(n_6598),
.Y(n_7477)
);

OAI22xp5_ASAP7_75t_L g7478 ( 
.A1(n_6207),
.A2(n_6135),
.B1(n_6040),
.B2(n_6088),
.Y(n_7478)
);

AOI22xp33_ASAP7_75t_SL g7479 ( 
.A1(n_6012),
.A2(n_5697),
.B1(n_5679),
.B2(n_5372),
.Y(n_7479)
);

AOI22xp33_ASAP7_75t_L g7480 ( 
.A1(n_6660),
.A2(n_5697),
.B1(n_5679),
.B2(n_5258),
.Y(n_7480)
);

BUFx6f_ASAP7_75t_L g7481 ( 
.A(n_6521),
.Y(n_7481)
);

AOI22xp33_ASAP7_75t_SL g7482 ( 
.A1(n_5801),
.A2(n_5697),
.B1(n_5372),
.B2(n_5384),
.Y(n_7482)
);

OAI22xp5_ASAP7_75t_L g7483 ( 
.A1(n_6088),
.A2(n_5348),
.B1(n_5265),
.B2(n_5587),
.Y(n_7483)
);

INVx6_ASAP7_75t_L g7484 ( 
.A(n_6524),
.Y(n_7484)
);

INVx3_ASAP7_75t_L g7485 ( 
.A(n_6598),
.Y(n_7485)
);

BUFx3_ASAP7_75t_L g7486 ( 
.A(n_6360),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_6144),
.Y(n_7487)
);

BUFx8_ASAP7_75t_L g7488 ( 
.A(n_6503),
.Y(n_7488)
);

BUFx4f_ASAP7_75t_SL g7489 ( 
.A(n_6247),
.Y(n_7489)
);

OAI22xp33_ASAP7_75t_L g7490 ( 
.A1(n_6414),
.A2(n_5539),
.B1(n_5381),
.B2(n_5384),
.Y(n_7490)
);

INVx4_ASAP7_75t_L g7491 ( 
.A(n_6665),
.Y(n_7491)
);

AOI22xp33_ASAP7_75t_SL g7492 ( 
.A1(n_5833),
.A2(n_5697),
.B1(n_5372),
.B2(n_5384),
.Y(n_7492)
);

INVx1_ASAP7_75t_L g7493 ( 
.A(n_6144),
.Y(n_7493)
);

OAI22xp33_ASAP7_75t_L g7494 ( 
.A1(n_6414),
.A2(n_5381),
.B1(n_5384),
.B2(n_5372),
.Y(n_7494)
);

AOI21xp5_ASAP7_75t_L g7495 ( 
.A1(n_5879),
.A2(n_5734),
.B(n_5659),
.Y(n_7495)
);

INVx2_ASAP7_75t_L g7496 ( 
.A(n_5808),
.Y(n_7496)
);

BUFx2_ASAP7_75t_SL g7497 ( 
.A(n_6521),
.Y(n_7497)
);

OAI22xp5_ASAP7_75t_L g7498 ( 
.A1(n_5921),
.A2(n_5785),
.B1(n_5908),
.B2(n_5822),
.Y(n_7498)
);

OAI21xp33_ASAP7_75t_L g7499 ( 
.A1(n_6645),
.A2(n_5188),
.B(n_5185),
.Y(n_7499)
);

AOI22xp33_ASAP7_75t_L g7500 ( 
.A1(n_6658),
.A2(n_5697),
.B1(n_5258),
.B2(n_5665),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_6149),
.Y(n_7501)
);

OAI22xp33_ASAP7_75t_SL g7502 ( 
.A1(n_6174),
.A2(n_5185),
.B1(n_5194),
.B2(n_5188),
.Y(n_7502)
);

NAND2xp5_ASAP7_75t_L g7503 ( 
.A(n_6163),
.B(n_5125),
.Y(n_7503)
);

CKINVDCx5p33_ASAP7_75t_R g7504 ( 
.A(n_6662),
.Y(n_7504)
);

INVx1_ASAP7_75t_L g7505 ( 
.A(n_6149),
.Y(n_7505)
);

INVx2_ASAP7_75t_SL g7506 ( 
.A(n_5887),
.Y(n_7506)
);

INVx3_ASAP7_75t_L g7507 ( 
.A(n_6598),
.Y(n_7507)
);

AOI22xp33_ASAP7_75t_L g7508 ( 
.A1(n_5860),
.A2(n_5697),
.B1(n_5258),
.B2(n_5665),
.Y(n_7508)
);

NAND2x1p5_ASAP7_75t_L g7509 ( 
.A(n_6324),
.B(n_5100),
.Y(n_7509)
);

BUFx6f_ASAP7_75t_L g7510 ( 
.A(n_6521),
.Y(n_7510)
);

AOI22xp33_ASAP7_75t_L g7511 ( 
.A1(n_5860),
.A2(n_5697),
.B1(n_5730),
.B2(n_5665),
.Y(n_7511)
);

INVx6_ASAP7_75t_L g7512 ( 
.A(n_6524),
.Y(n_7512)
);

BUFx8_ASAP7_75t_SL g7513 ( 
.A(n_6247),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_6150),
.Y(n_7514)
);

AOI22xp33_ASAP7_75t_L g7515 ( 
.A1(n_5891),
.A2(n_5697),
.B1(n_5730),
.B2(n_5665),
.Y(n_7515)
);

OAI22xp5_ASAP7_75t_L g7516 ( 
.A1(n_5921),
.A2(n_5619),
.B1(n_5255),
.B2(n_5256),
.Y(n_7516)
);

OAI22xp5_ASAP7_75t_SL g7517 ( 
.A1(n_6666),
.A2(n_5372),
.B1(n_5384),
.B2(n_5381),
.Y(n_7517)
);

INVx3_ASAP7_75t_SL g7518 ( 
.A(n_6348),
.Y(n_7518)
);

CKINVDCx20_ASAP7_75t_R g7519 ( 
.A(n_6247),
.Y(n_7519)
);

AOI22xp33_ASAP7_75t_L g7520 ( 
.A1(n_6148),
.A2(n_5783),
.B1(n_5730),
.B2(n_5259),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_6150),
.Y(n_7521)
);

INVx2_ASAP7_75t_SL g7522 ( 
.A(n_5887),
.Y(n_7522)
);

BUFx3_ASAP7_75t_L g7523 ( 
.A(n_6360),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6152),
.Y(n_7524)
);

CKINVDCx11_ASAP7_75t_R g7525 ( 
.A(n_6288),
.Y(n_7525)
);

AOI22xp33_ASAP7_75t_L g7526 ( 
.A1(n_6148),
.A2(n_5783),
.B1(n_5730),
.B2(n_5313),
.Y(n_7526)
);

INVx6_ASAP7_75t_L g7527 ( 
.A(n_6524),
.Y(n_7527)
);

AOI22xp33_ASAP7_75t_L g7528 ( 
.A1(n_6255),
.A2(n_5783),
.B1(n_5313),
.B2(n_5333),
.Y(n_7528)
);

BUFx6f_ASAP7_75t_L g7529 ( 
.A(n_6548),
.Y(n_7529)
);

INVx1_ASAP7_75t_SL g7530 ( 
.A(n_5970),
.Y(n_7530)
);

BUFx3_ASAP7_75t_L g7531 ( 
.A(n_6360),
.Y(n_7531)
);

NAND2x1p5_ASAP7_75t_L g7532 ( 
.A(n_6324),
.B(n_5100),
.Y(n_7532)
);

NAND2x1p5_ASAP7_75t_L g7533 ( 
.A(n_6324),
.B(n_5100),
.Y(n_7533)
);

BUFx6f_ASAP7_75t_L g7534 ( 
.A(n_6548),
.Y(n_7534)
);

AOI22xp33_ASAP7_75t_L g7535 ( 
.A1(n_6255),
.A2(n_5783),
.B1(n_5313),
.B2(n_5333),
.Y(n_7535)
);

BUFx3_ASAP7_75t_L g7536 ( 
.A(n_6360),
.Y(n_7536)
);

AOI22xp33_ASAP7_75t_L g7537 ( 
.A1(n_5833),
.A2(n_5313),
.B1(n_5333),
.B2(n_5309),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_6152),
.Y(n_7538)
);

BUFx2_ASAP7_75t_L g7539 ( 
.A(n_6161),
.Y(n_7539)
);

AOI22xp33_ASAP7_75t_L g7540 ( 
.A1(n_5862),
.A2(n_5924),
.B1(n_5945),
.B2(n_5883),
.Y(n_7540)
);

BUFx3_ASAP7_75t_L g7541 ( 
.A(n_6360),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_6157),
.Y(n_7542)
);

CKINVDCx20_ASAP7_75t_R g7543 ( 
.A(n_6288),
.Y(n_7543)
);

NAND2xp5_ASAP7_75t_L g7544 ( 
.A(n_6163),
.B(n_5125),
.Y(n_7544)
);

INVx2_ASAP7_75t_L g7545 ( 
.A(n_5808),
.Y(n_7545)
);

AOI22xp33_ASAP7_75t_L g7546 ( 
.A1(n_5862),
.A2(n_5924),
.B1(n_5945),
.B2(n_5883),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_5808),
.Y(n_7547)
);

AOI22xp33_ASAP7_75t_L g7548 ( 
.A1(n_5862),
.A2(n_5313),
.B1(n_5333),
.B2(n_5309),
.Y(n_7548)
);

OAI22xp5_ASAP7_75t_L g7549 ( 
.A1(n_5785),
.A2(n_5619),
.B1(n_5255),
.B2(n_5256),
.Y(n_7549)
);

AOI22xp5_ASAP7_75t_L g7550 ( 
.A1(n_5788),
.A2(n_5736),
.B1(n_5748),
.B2(n_5585),
.Y(n_7550)
);

AOI22xp33_ASAP7_75t_L g7551 ( 
.A1(n_5862),
.A2(n_5924),
.B1(n_5945),
.B2(n_5883),
.Y(n_7551)
);

AOI22xp5_ASAP7_75t_L g7552 ( 
.A1(n_5788),
.A2(n_5736),
.B1(n_5748),
.B2(n_5585),
.Y(n_7552)
);

CKINVDCx6p67_ASAP7_75t_R g7553 ( 
.A(n_6288),
.Y(n_7553)
);

INVx1_ASAP7_75t_L g7554 ( 
.A(n_6157),
.Y(n_7554)
);

CKINVDCx11_ASAP7_75t_R g7555 ( 
.A(n_6288),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_6165),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_6165),
.Y(n_7557)
);

INVx4_ASAP7_75t_L g7558 ( 
.A(n_5848),
.Y(n_7558)
);

INVx4_ASAP7_75t_L g7559 ( 
.A(n_5848),
.Y(n_7559)
);

INVx4_ASAP7_75t_L g7560 ( 
.A(n_5848),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_6180),
.Y(n_7561)
);

INVx2_ASAP7_75t_L g7562 ( 
.A(n_5814),
.Y(n_7562)
);

AOI22xp5_ASAP7_75t_L g7563 ( 
.A1(n_6105),
.A2(n_5585),
.B1(n_5381),
.B2(n_5384),
.Y(n_7563)
);

INVx4_ASAP7_75t_L g7564 ( 
.A(n_5865),
.Y(n_7564)
);

BUFx3_ASAP7_75t_L g7565 ( 
.A(n_6360),
.Y(n_7565)
);

OAI22xp5_ASAP7_75t_L g7566 ( 
.A1(n_5785),
.A2(n_5619),
.B1(n_5255),
.B2(n_5256),
.Y(n_7566)
);

CKINVDCx6p67_ASAP7_75t_R g7567 ( 
.A(n_6289),
.Y(n_7567)
);

OAI21xp5_ASAP7_75t_SL g7568 ( 
.A1(n_6178),
.A2(n_5150),
.B(n_5585),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_6180),
.Y(n_7569)
);

BUFx10_ASAP7_75t_L g7570 ( 
.A(n_6548),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_6182),
.Y(n_7571)
);

INVx4_ASAP7_75t_L g7572 ( 
.A(n_6665),
.Y(n_7572)
);

AOI22xp5_ASAP7_75t_L g7573 ( 
.A1(n_6105),
.A2(n_5381),
.B1(n_5384),
.B2(n_5372),
.Y(n_7573)
);

BUFx2_ASAP7_75t_SL g7574 ( 
.A(n_6548),
.Y(n_7574)
);

BUFx12f_ASAP7_75t_L g7575 ( 
.A(n_5865),
.Y(n_7575)
);

BUFx6f_ASAP7_75t_L g7576 ( 
.A(n_6548),
.Y(n_7576)
);

BUFx4f_ASAP7_75t_SL g7577 ( 
.A(n_6289),
.Y(n_7577)
);

AOI22xp33_ASAP7_75t_L g7578 ( 
.A1(n_5883),
.A2(n_5313),
.B1(n_5333),
.B2(n_5309),
.Y(n_7578)
);

AOI22xp33_ASAP7_75t_L g7579 ( 
.A1(n_5924),
.A2(n_5313),
.B1(n_5333),
.B2(n_5309),
.Y(n_7579)
);

INVx3_ASAP7_75t_L g7580 ( 
.A(n_6602),
.Y(n_7580)
);

INVx1_ASAP7_75t_SL g7581 ( 
.A(n_5970),
.Y(n_7581)
);

INVx1_ASAP7_75t_L g7582 ( 
.A(n_6182),
.Y(n_7582)
);

NAND2xp5_ASAP7_75t_L g7583 ( 
.A(n_6217),
.B(n_5130),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_6185),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_6185),
.Y(n_7585)
);

HB1xp67_ASAP7_75t_L g7586 ( 
.A(n_6193),
.Y(n_7586)
);

INVx6_ASAP7_75t_L g7587 ( 
.A(n_6548),
.Y(n_7587)
);

AOI22xp33_ASAP7_75t_L g7588 ( 
.A1(n_5945),
.A2(n_5333),
.B1(n_5342),
.B2(n_5309),
.Y(n_7588)
);

BUFx4f_ASAP7_75t_L g7589 ( 
.A(n_6597),
.Y(n_7589)
);

BUFx12f_ASAP7_75t_L g7590 ( 
.A(n_5865),
.Y(n_7590)
);

OAI22xp5_ASAP7_75t_L g7591 ( 
.A1(n_5822),
.A2(n_5619),
.B1(n_5255),
.B2(n_5256),
.Y(n_7591)
);

INVx2_ASAP7_75t_L g7592 ( 
.A(n_5814),
.Y(n_7592)
);

NAND2xp5_ASAP7_75t_L g7593 ( 
.A(n_6217),
.B(n_6609),
.Y(n_7593)
);

INVx6_ASAP7_75t_L g7594 ( 
.A(n_6548),
.Y(n_7594)
);

INVx2_ASAP7_75t_L g7595 ( 
.A(n_5814),
.Y(n_7595)
);

AOI22xp5_ASAP7_75t_L g7596 ( 
.A1(n_6046),
.A2(n_5774),
.B1(n_5775),
.B2(n_5767),
.Y(n_7596)
);

AOI22xp33_ASAP7_75t_SL g7597 ( 
.A1(n_5822),
.A2(n_5381),
.B1(n_5384),
.B2(n_5372),
.Y(n_7597)
);

AOI22xp5_ASAP7_75t_L g7598 ( 
.A1(n_6046),
.A2(n_5774),
.B1(n_5775),
.B2(n_5767),
.Y(n_7598)
);

OAI21xp33_ASAP7_75t_L g7599 ( 
.A1(n_6309),
.A2(n_5188),
.B(n_5185),
.Y(n_7599)
);

AOI22xp33_ASAP7_75t_L g7600 ( 
.A1(n_5962),
.A2(n_5342),
.B1(n_5309),
.B2(n_5343),
.Y(n_7600)
);

OAI22x1_ASAP7_75t_L g7601 ( 
.A1(n_6187),
.A2(n_5194),
.B1(n_5224),
.B2(n_5215),
.Y(n_7601)
);

AOI22xp33_ASAP7_75t_L g7602 ( 
.A1(n_5962),
.A2(n_5342),
.B1(n_5309),
.B2(n_5343),
.Y(n_7602)
);

INVx2_ASAP7_75t_L g7603 ( 
.A(n_5814),
.Y(n_7603)
);

INVx2_ASAP7_75t_L g7604 ( 
.A(n_5858),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_6190),
.Y(n_7605)
);

NAND2xp5_ASAP7_75t_L g7606 ( 
.A(n_6609),
.B(n_5130),
.Y(n_7606)
);

OAI22xp5_ASAP7_75t_L g7607 ( 
.A1(n_5908),
.A2(n_5241),
.B1(n_5198),
.B2(n_5193),
.Y(n_7607)
);

BUFx3_ASAP7_75t_L g7608 ( 
.A(n_6628),
.Y(n_7608)
);

BUFx2_ASAP7_75t_L g7609 ( 
.A(n_6161),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_6190),
.Y(n_7610)
);

CKINVDCx20_ASAP7_75t_R g7611 ( 
.A(n_6289),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_6192),
.Y(n_7612)
);

AND2x2_ASAP7_75t_L g7613 ( 
.A(n_6545),
.B(n_5543),
.Y(n_7613)
);

AOI22xp33_ASAP7_75t_L g7614 ( 
.A1(n_5962),
.A2(n_5997),
.B1(n_6015),
.B2(n_5972),
.Y(n_7614)
);

BUFx2_ASAP7_75t_SL g7615 ( 
.A(n_6548),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_6192),
.Y(n_7616)
);

INVx6_ASAP7_75t_L g7617 ( 
.A(n_6592),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_5858),
.Y(n_7618)
);

CKINVDCx6p67_ASAP7_75t_R g7619 ( 
.A(n_6289),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_6199),
.Y(n_7620)
);

INVx1_ASAP7_75t_SL g7621 ( 
.A(n_6006),
.Y(n_7621)
);

BUFx8_ASAP7_75t_L g7622 ( 
.A(n_6503),
.Y(n_7622)
);

AOI22xp33_ASAP7_75t_SL g7623 ( 
.A1(n_5908),
.A2(n_5381),
.B1(n_5402),
.B2(n_5372),
.Y(n_7623)
);

INVx6_ASAP7_75t_L g7624 ( 
.A(n_6592),
.Y(n_7624)
);

BUFx4_ASAP7_75t_R g7625 ( 
.A(n_6292),
.Y(n_7625)
);

INVx2_ASAP7_75t_L g7626 ( 
.A(n_5858),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_6199),
.Y(n_7627)
);

BUFx8_ASAP7_75t_SL g7628 ( 
.A(n_6292),
.Y(n_7628)
);

AOI22xp33_ASAP7_75t_SL g7629 ( 
.A1(n_6000),
.A2(n_5402),
.B1(n_5404),
.B2(n_5381),
.Y(n_7629)
);

OAI22xp5_ASAP7_75t_L g7630 ( 
.A1(n_6000),
.A2(n_6120),
.B1(n_6127),
.B2(n_6087),
.Y(n_7630)
);

INVx2_ASAP7_75t_L g7631 ( 
.A(n_5858),
.Y(n_7631)
);

AOI21xp5_ASAP7_75t_L g7632 ( 
.A1(n_5879),
.A2(n_5734),
.B(n_5659),
.Y(n_7632)
);

NAND2x1_ASAP7_75t_L g7633 ( 
.A(n_6161),
.B(n_5272),
.Y(n_7633)
);

CKINVDCx20_ASAP7_75t_R g7634 ( 
.A(n_6292),
.Y(n_7634)
);

OAI22xp5_ASAP7_75t_L g7635 ( 
.A1(n_6000),
.A2(n_5241),
.B1(n_5198),
.B2(n_5193),
.Y(n_7635)
);

NAND2xp5_ASAP7_75t_SL g7636 ( 
.A(n_6547),
.B(n_5268),
.Y(n_7636)
);

BUFx3_ASAP7_75t_L g7637 ( 
.A(n_6628),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_5874),
.Y(n_7638)
);

BUFx3_ASAP7_75t_L g7639 ( 
.A(n_6628),
.Y(n_7639)
);

CKINVDCx20_ASAP7_75t_R g7640 ( 
.A(n_6292),
.Y(n_7640)
);

INVx6_ASAP7_75t_L g7641 ( 
.A(n_6592),
.Y(n_7641)
);

AOI22xp33_ASAP7_75t_L g7642 ( 
.A1(n_5962),
.A2(n_5342),
.B1(n_5344),
.B2(n_5343),
.Y(n_7642)
);

INVx3_ASAP7_75t_L g7643 ( 
.A(n_6602),
.Y(n_7643)
);

INVx6_ASAP7_75t_L g7644 ( 
.A(n_6592),
.Y(n_7644)
);

INVx4_ASAP7_75t_L g7645 ( 
.A(n_5865),
.Y(n_7645)
);

INVx1_ASAP7_75t_SL g7646 ( 
.A(n_6006),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_6214),
.Y(n_7647)
);

OAI22xp33_ASAP7_75t_L g7648 ( 
.A1(n_6414),
.A2(n_5402),
.B1(n_5411),
.B2(n_5404),
.Y(n_7648)
);

OAI22xp33_ASAP7_75t_L g7649 ( 
.A1(n_6641),
.A2(n_6256),
.B1(n_6191),
.B2(n_6305),
.Y(n_7649)
);

INVx2_ASAP7_75t_SL g7650 ( 
.A(n_5887),
.Y(n_7650)
);

INVx3_ASAP7_75t_L g7651 ( 
.A(n_6602),
.Y(n_7651)
);

INVx2_ASAP7_75t_L g7652 ( 
.A(n_5874),
.Y(n_7652)
);

CKINVDCx11_ASAP7_75t_R g7653 ( 
.A(n_6320),
.Y(n_7653)
);

OAI21xp33_ASAP7_75t_L g7654 ( 
.A1(n_6309),
.A2(n_5215),
.B(n_5194),
.Y(n_7654)
);

BUFx6f_ASAP7_75t_L g7655 ( 
.A(n_6592),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_5874),
.Y(n_7656)
);

AOI22xp33_ASAP7_75t_L g7657 ( 
.A1(n_5972),
.A2(n_5342),
.B1(n_5344),
.B2(n_5343),
.Y(n_7657)
);

BUFx2_ASAP7_75t_L g7658 ( 
.A(n_6161),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_6214),
.Y(n_7659)
);

OAI22xp5_ASAP7_75t_L g7660 ( 
.A1(n_6059),
.A2(n_5241),
.B1(n_5198),
.B2(n_5193),
.Y(n_7660)
);

BUFx6f_ASAP7_75t_L g7661 ( 
.A(n_6592),
.Y(n_7661)
);

BUFx3_ASAP7_75t_L g7662 ( 
.A(n_6628),
.Y(n_7662)
);

BUFx10_ASAP7_75t_L g7663 ( 
.A(n_6592),
.Y(n_7663)
);

INVx6_ASAP7_75t_L g7664 ( 
.A(n_6592),
.Y(n_7664)
);

AOI22xp33_ASAP7_75t_L g7665 ( 
.A1(n_5972),
.A2(n_5342),
.B1(n_5344),
.B2(n_5343),
.Y(n_7665)
);

INVx3_ASAP7_75t_L g7666 ( 
.A(n_6602),
.Y(n_7666)
);

BUFx12f_ASAP7_75t_L g7667 ( 
.A(n_5865),
.Y(n_7667)
);

AOI22xp33_ASAP7_75t_L g7668 ( 
.A1(n_5972),
.A2(n_5342),
.B1(n_5344),
.B2(n_5343),
.Y(n_7668)
);

CKINVDCx5p33_ASAP7_75t_R g7669 ( 
.A(n_6662),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_6232),
.Y(n_7670)
);

INVx1_ASAP7_75t_SL g7671 ( 
.A(n_6049),
.Y(n_7671)
);

AOI22xp33_ASAP7_75t_L g7672 ( 
.A1(n_5997),
.A2(n_5344),
.B1(n_5343),
.B2(n_5292),
.Y(n_7672)
);

INVx2_ASAP7_75t_L g7673 ( 
.A(n_5874),
.Y(n_7673)
);

INVx6_ASAP7_75t_L g7674 ( 
.A(n_6597),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_5875),
.Y(n_7675)
);

HB1xp67_ASAP7_75t_L g7676 ( 
.A(n_6193),
.Y(n_7676)
);

AOI22xp33_ASAP7_75t_L g7677 ( 
.A1(n_5997),
.A2(n_5344),
.B1(n_5292),
.B2(n_5304),
.Y(n_7677)
);

BUFx2_ASAP7_75t_L g7678 ( 
.A(n_5997),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_6232),
.Y(n_7679)
);

AOI22xp33_ASAP7_75t_SL g7680 ( 
.A1(n_6087),
.A2(n_5402),
.B1(n_5404),
.B2(n_5381),
.Y(n_7680)
);

CKINVDCx6p67_ASAP7_75t_R g7681 ( 
.A(n_6320),
.Y(n_7681)
);

CKINVDCx20_ASAP7_75t_R g7682 ( 
.A(n_6320),
.Y(n_7682)
);

INVx6_ASAP7_75t_L g7683 ( 
.A(n_6597),
.Y(n_7683)
);

INVx8_ASAP7_75t_L g7684 ( 
.A(n_5798),
.Y(n_7684)
);

INVx2_ASAP7_75t_L g7685 ( 
.A(n_5875),
.Y(n_7685)
);

BUFx3_ASAP7_75t_L g7686 ( 
.A(n_6628),
.Y(n_7686)
);

INVx1_ASAP7_75t_L g7687 ( 
.A(n_6244),
.Y(n_7687)
);

INVx4_ASAP7_75t_L g7688 ( 
.A(n_5919),
.Y(n_7688)
);

INVx4_ASAP7_75t_L g7689 ( 
.A(n_5919),
.Y(n_7689)
);

OAI22xp5_ASAP7_75t_SL g7690 ( 
.A1(n_6619),
.A2(n_5404),
.B1(n_5406),
.B2(n_5402),
.Y(n_7690)
);

BUFx6f_ASAP7_75t_L g7691 ( 
.A(n_6597),
.Y(n_7691)
);

AOI22xp33_ASAP7_75t_L g7692 ( 
.A1(n_6015),
.A2(n_5344),
.B1(n_5304),
.B2(n_5272),
.Y(n_7692)
);

AOI22xp5_ASAP7_75t_L g7693 ( 
.A1(n_6431),
.A2(n_5402),
.B1(n_5406),
.B2(n_5404),
.Y(n_7693)
);

INVx1_ASAP7_75t_L g7694 ( 
.A(n_6244),
.Y(n_7694)
);

AND2x2_ASAP7_75t_L g7695 ( 
.A(n_6545),
.B(n_5543),
.Y(n_7695)
);

INVx2_ASAP7_75t_L g7696 ( 
.A(n_5875),
.Y(n_7696)
);

AOI22xp33_ASAP7_75t_SL g7697 ( 
.A1(n_6087),
.A2(n_5404),
.B1(n_5406),
.B2(n_5402),
.Y(n_7697)
);

CKINVDCx14_ASAP7_75t_R g7698 ( 
.A(n_6628),
.Y(n_7698)
);

BUFx12f_ASAP7_75t_L g7699 ( 
.A(n_5919),
.Y(n_7699)
);

NOR3xp33_ASAP7_75t_L g7700 ( 
.A(n_6641),
.B(n_6121),
.C(n_6080),
.Y(n_7700)
);

NAND2xp5_ASAP7_75t_L g7701 ( 
.A(n_6619),
.B(n_5200),
.Y(n_7701)
);

AOI22xp33_ASAP7_75t_L g7702 ( 
.A1(n_6015),
.A2(n_5304),
.B1(n_5354),
.B2(n_5272),
.Y(n_7702)
);

BUFx12f_ASAP7_75t_L g7703 ( 
.A(n_5919),
.Y(n_7703)
);

INVx4_ASAP7_75t_SL g7704 ( 
.A(n_6004),
.Y(n_7704)
);

OAI22xp5_ASAP7_75t_L g7705 ( 
.A1(n_6120),
.A2(n_5241),
.B1(n_5198),
.B2(n_5193),
.Y(n_7705)
);

NAND2xp5_ASAP7_75t_L g7706 ( 
.A(n_6643),
.B(n_5723),
.Y(n_7706)
);

OAI22xp33_ASAP7_75t_L g7707 ( 
.A1(n_6256),
.A2(n_5404),
.B1(n_5406),
.B2(n_5402),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_6249),
.Y(n_7708)
);

NAND2xp5_ASAP7_75t_L g7709 ( 
.A(n_6643),
.B(n_5723),
.Y(n_7709)
);

CKINVDCx11_ASAP7_75t_R g7710 ( 
.A(n_6320),
.Y(n_7710)
);

BUFx6f_ASAP7_75t_L g7711 ( 
.A(n_6597),
.Y(n_7711)
);

OAI22x1_ASAP7_75t_SL g7712 ( 
.A1(n_5919),
.A2(n_5595),
.B1(n_5677),
.B2(n_5608),
.Y(n_7712)
);

CKINVDCx16_ASAP7_75t_R g7713 ( 
.A(n_6323),
.Y(n_7713)
);

BUFx6f_ASAP7_75t_L g7714 ( 
.A(n_6597),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_6249),
.Y(n_7715)
);

BUFx2_ASAP7_75t_L g7716 ( 
.A(n_6015),
.Y(n_7716)
);

OAI22xp33_ASAP7_75t_L g7717 ( 
.A1(n_6191),
.A2(n_5404),
.B1(n_5406),
.B2(n_5402),
.Y(n_7717)
);

AOI22xp33_ASAP7_75t_L g7718 ( 
.A1(n_6052),
.A2(n_5304),
.B1(n_5354),
.B2(n_5272),
.Y(n_7718)
);

INVx3_ASAP7_75t_L g7719 ( 
.A(n_6602),
.Y(n_7719)
);

CKINVDCx11_ASAP7_75t_R g7720 ( 
.A(n_6323),
.Y(n_7720)
);

AOI22xp33_ASAP7_75t_SL g7721 ( 
.A1(n_6059),
.A2(n_5404),
.B1(n_5406),
.B2(n_5402),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_6266),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_6266),
.Y(n_7723)
);

AOI22xp33_ASAP7_75t_L g7724 ( 
.A1(n_6052),
.A2(n_5354),
.B1(n_5379),
.B2(n_5361),
.Y(n_7724)
);

INVx6_ASAP7_75t_L g7725 ( 
.A(n_6597),
.Y(n_7725)
);

CKINVDCx11_ASAP7_75t_R g7726 ( 
.A(n_6323),
.Y(n_7726)
);

INVx1_ASAP7_75t_SL g7727 ( 
.A(n_6049),
.Y(n_7727)
);

BUFx10_ASAP7_75t_L g7728 ( 
.A(n_6597),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_6270),
.Y(n_7729)
);

AOI22xp33_ASAP7_75t_L g7730 ( 
.A1(n_6052),
.A2(n_5354),
.B1(n_5379),
.B2(n_5361),
.Y(n_7730)
);

INVx1_ASAP7_75t_L g7731 ( 
.A(n_6270),
.Y(n_7731)
);

INVx6_ASAP7_75t_L g7732 ( 
.A(n_6638),
.Y(n_7732)
);

AOI22xp33_ASAP7_75t_L g7733 ( 
.A1(n_6052),
.A2(n_5379),
.B1(n_5361),
.B2(n_5600),
.Y(n_7733)
);

AOI22xp5_ASAP7_75t_L g7734 ( 
.A1(n_6431),
.A2(n_5406),
.B1(n_5411),
.B2(n_5404),
.Y(n_7734)
);

BUFx8_ASAP7_75t_L g7735 ( 
.A(n_6503),
.Y(n_7735)
);

BUFx12f_ASAP7_75t_L g7736 ( 
.A(n_5985),
.Y(n_7736)
);

INVx1_ASAP7_75t_L g7737 ( 
.A(n_6281),
.Y(n_7737)
);

AOI22xp33_ASAP7_75t_SL g7738 ( 
.A1(n_6059),
.A2(n_5411),
.B1(n_5417),
.B2(n_5406),
.Y(n_7738)
);

NAND2xp5_ASAP7_75t_L g7739 ( 
.A(n_6644),
.B(n_5601),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6281),
.Y(n_7740)
);

INVx1_ASAP7_75t_SL g7741 ( 
.A(n_6086),
.Y(n_7741)
);

CKINVDCx11_ASAP7_75t_R g7742 ( 
.A(n_6323),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_6644),
.B(n_5601),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_6285),
.Y(n_7744)
);

OAI21xp5_ASAP7_75t_SL g7745 ( 
.A1(n_6178),
.A2(n_6061),
.B(n_6242),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_6285),
.Y(n_7746)
);

NAND2xp5_ASAP7_75t_L g7747 ( 
.A(n_6655),
.B(n_5602),
.Y(n_7747)
);

AOI22xp33_ASAP7_75t_L g7748 ( 
.A1(n_6064),
.A2(n_5379),
.B1(n_5361),
.B2(n_5600),
.Y(n_7748)
);

INVx2_ASAP7_75t_L g7749 ( 
.A(n_5875),
.Y(n_7749)
);

INVx6_ASAP7_75t_L g7750 ( 
.A(n_6638),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_6655),
.B(n_5602),
.Y(n_7751)
);

CKINVDCx20_ASAP7_75t_R g7752 ( 
.A(n_6371),
.Y(n_7752)
);

INVx1_ASAP7_75t_L g7753 ( 
.A(n_6294),
.Y(n_7753)
);

BUFx12f_ASAP7_75t_L g7754 ( 
.A(n_5985),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_6294),
.Y(n_7755)
);

AOI22xp33_ASAP7_75t_L g7756 ( 
.A1(n_6064),
.A2(n_6098),
.B1(n_6067),
.B2(n_6396),
.Y(n_7756)
);

INVx6_ASAP7_75t_L g7757 ( 
.A(n_6638),
.Y(n_7757)
);

BUFx8_ASAP7_75t_SL g7758 ( 
.A(n_6371),
.Y(n_7758)
);

BUFx4f_ASAP7_75t_L g7759 ( 
.A(n_6638),
.Y(n_7759)
);

OAI22xp33_ASAP7_75t_L g7760 ( 
.A1(n_6305),
.A2(n_5411),
.B1(n_5417),
.B2(n_5406),
.Y(n_7760)
);

BUFx2_ASAP7_75t_L g7761 ( 
.A(n_6064),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_5904),
.Y(n_7762)
);

INVx1_ASAP7_75t_L g7763 ( 
.A(n_6300),
.Y(n_7763)
);

AOI22xp33_ASAP7_75t_SL g7764 ( 
.A1(n_6071),
.A2(n_5411),
.B1(n_5417),
.B2(n_5406),
.Y(n_7764)
);

OAI22x1_ASAP7_75t_L g7765 ( 
.A1(n_6071),
.A2(n_5215),
.B1(n_5229),
.B2(n_5224),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_6300),
.Y(n_7766)
);

INVx2_ASAP7_75t_SL g7767 ( 
.A(n_5931),
.Y(n_7767)
);

INVx2_ASAP7_75t_L g7768 ( 
.A(n_5904),
.Y(n_7768)
);

BUFx10_ASAP7_75t_L g7769 ( 
.A(n_6638),
.Y(n_7769)
);

AOI22xp33_ASAP7_75t_L g7770 ( 
.A1(n_6064),
.A2(n_5635),
.B1(n_5656),
.B2(n_5600),
.Y(n_7770)
);

INVx2_ASAP7_75t_L g7771 ( 
.A(n_5904),
.Y(n_7771)
);

AOI22xp33_ASAP7_75t_L g7772 ( 
.A1(n_6067),
.A2(n_5635),
.B1(n_5656),
.B2(n_5600),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_6301),
.Y(n_7773)
);

AOI22xp33_ASAP7_75t_L g7774 ( 
.A1(n_6067),
.A2(n_5635),
.B1(n_5656),
.B2(n_5600),
.Y(n_7774)
);

BUFx3_ASAP7_75t_L g7775 ( 
.A(n_6642),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_6301),
.Y(n_7776)
);

INVx6_ASAP7_75t_L g7777 ( 
.A(n_6638),
.Y(n_7777)
);

AOI22xp33_ASAP7_75t_SL g7778 ( 
.A1(n_6071),
.A2(n_5417),
.B1(n_5420),
.B2(n_5411),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_6322),
.Y(n_7779)
);

BUFx4_ASAP7_75t_SL g7780 ( 
.A(n_6371),
.Y(n_7780)
);

CKINVDCx6p67_ASAP7_75t_R g7781 ( 
.A(n_6371),
.Y(n_7781)
);

INVx8_ASAP7_75t_L g7782 ( 
.A(n_5798),
.Y(n_7782)
);

INVx6_ASAP7_75t_L g7783 ( 
.A(n_6638),
.Y(n_7783)
);

INVx6_ASAP7_75t_L g7784 ( 
.A(n_6638),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_6322),
.Y(n_7785)
);

AOI22xp33_ASAP7_75t_SL g7786 ( 
.A1(n_6120),
.A2(n_5417),
.B1(n_5420),
.B2(n_5411),
.Y(n_7786)
);

CKINVDCx5p33_ASAP7_75t_R g7787 ( 
.A(n_6662),
.Y(n_7787)
);

INVx1_ASAP7_75t_SL g7788 ( 
.A(n_6086),
.Y(n_7788)
);

AOI22xp33_ASAP7_75t_L g7789 ( 
.A1(n_6067),
.A2(n_5635),
.B1(n_5656),
.B2(n_5600),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_6326),
.Y(n_7790)
);

BUFx12f_ASAP7_75t_L g7791 ( 
.A(n_5985),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_6326),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_6778),
.Y(n_7793)
);

INVx2_ASAP7_75t_L g7794 ( 
.A(n_7344),
.Y(n_7794)
);

OAI21x1_ASAP7_75t_L g7795 ( 
.A1(n_6949),
.A2(n_6543),
.B(n_6575),
.Y(n_7795)
);

OR2x6_ASAP7_75t_L g7796 ( 
.A(n_6870),
.B(n_6635),
.Y(n_7796)
);

INVx1_ASAP7_75t_L g7797 ( 
.A(n_6778),
.Y(n_7797)
);

BUFx8_ASAP7_75t_L g7798 ( 
.A(n_6918),
.Y(n_7798)
);

NAND2xp5_ASAP7_75t_L g7799 ( 
.A(n_6900),
.B(n_6657),
.Y(n_7799)
);

INVx1_ASAP7_75t_L g7800 ( 
.A(n_6779),
.Y(n_7800)
);

BUFx4f_ASAP7_75t_L g7801 ( 
.A(n_6776),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_6779),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_7344),
.Y(n_7803)
);

CKINVDCx5p33_ASAP7_75t_R g7804 ( 
.A(n_6721),
.Y(n_7804)
);

OAI21x1_ASAP7_75t_L g7805 ( 
.A1(n_6949),
.A2(n_6543),
.B(n_6575),
.Y(n_7805)
);

INVx1_ASAP7_75t_L g7806 ( 
.A(n_6675),
.Y(n_7806)
);

BUFx2_ASAP7_75t_L g7807 ( 
.A(n_6907),
.Y(n_7807)
);

INVx2_ASAP7_75t_L g7808 ( 
.A(n_7344),
.Y(n_7808)
);

CKINVDCx5p33_ASAP7_75t_R g7809 ( 
.A(n_6741),
.Y(n_7809)
);

CKINVDCx5p33_ASAP7_75t_R g7810 ( 
.A(n_6938),
.Y(n_7810)
);

AOI22xp33_ASAP7_75t_L g7811 ( 
.A1(n_6780),
.A2(n_6109),
.B1(n_6041),
.B2(n_6080),
.Y(n_7811)
);

HB1xp67_ASAP7_75t_L g7812 ( 
.A(n_6910),
.Y(n_7812)
);

INVx2_ASAP7_75t_L g7813 ( 
.A(n_7359),
.Y(n_7813)
);

AO21x2_ASAP7_75t_L g7814 ( 
.A1(n_7158),
.A2(n_5784),
.B(n_5935),
.Y(n_7814)
);

INVx2_ASAP7_75t_L g7815 ( 
.A(n_7359),
.Y(n_7815)
);

INVx4_ASAP7_75t_L g7816 ( 
.A(n_6713),
.Y(n_7816)
);

INVx3_ASAP7_75t_SL g7817 ( 
.A(n_6776),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_6675),
.Y(n_7818)
);

INVx2_ASAP7_75t_L g7819 ( 
.A(n_7359),
.Y(n_7819)
);

INVx3_ASAP7_75t_L g7820 ( 
.A(n_7633),
.Y(n_7820)
);

INVx2_ASAP7_75t_SL g7821 ( 
.A(n_6705),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_6684),
.Y(n_7822)
);

HB1xp67_ASAP7_75t_L g7823 ( 
.A(n_6910),
.Y(n_7823)
);

NAND2xp5_ASAP7_75t_L g7824 ( 
.A(n_6900),
.B(n_6657),
.Y(n_7824)
);

AOI221xp5_ASAP7_75t_L g7825 ( 
.A1(n_6780),
.A2(n_6109),
.B1(n_6219),
.B2(n_6224),
.C(n_6218),
.Y(n_7825)
);

BUFx6f_ASAP7_75t_L g7826 ( 
.A(n_6700),
.Y(n_7826)
);

AOI22xp33_ASAP7_75t_L g7827 ( 
.A1(n_6853),
.A2(n_6041),
.B1(n_5825),
.B2(n_6083),
.Y(n_7827)
);

AO21x1_ASAP7_75t_SL g7828 ( 
.A1(n_6790),
.A2(n_6295),
.B(n_6172),
.Y(n_7828)
);

INVx3_ASAP7_75t_L g7829 ( 
.A(n_7633),
.Y(n_7829)
);

AOI22xp5_ASAP7_75t_L g7830 ( 
.A1(n_6846),
.A2(n_6061),
.B1(n_6229),
.B2(n_6213),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_6684),
.Y(n_7831)
);

INVx2_ASAP7_75t_SL g7832 ( 
.A(n_6705),
.Y(n_7832)
);

BUFx3_ASAP7_75t_L g7833 ( 
.A(n_7197),
.Y(n_7833)
);

AND2x2_ASAP7_75t_L g7834 ( 
.A(n_7021),
.B(n_6127),
.Y(n_7834)
);

OAI21x1_ASAP7_75t_L g7835 ( 
.A1(n_6949),
.A2(n_6543),
.B(n_6575),
.Y(n_7835)
);

INVx1_ASAP7_75t_L g7836 ( 
.A(n_6687),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_6687),
.Y(n_7837)
);

AO21x2_ASAP7_75t_L g7838 ( 
.A1(n_7158),
.A2(n_5784),
.B(n_5935),
.Y(n_7838)
);

AO21x2_ASAP7_75t_L g7839 ( 
.A1(n_7494),
.A2(n_7648),
.B(n_7159),
.Y(n_7839)
);

BUFx6f_ASAP7_75t_L g7840 ( 
.A(n_6700),
.Y(n_7840)
);

OAI21xp5_ASAP7_75t_L g7841 ( 
.A1(n_6699),
.A2(n_6242),
.B(n_6029),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_6706),
.Y(n_7842)
);

INVx2_ASAP7_75t_L g7843 ( 
.A(n_7366),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_6853),
.A2(n_6041),
.B1(n_5825),
.B2(n_6083),
.Y(n_7844)
);

BUFx2_ASAP7_75t_L g7845 ( 
.A(n_6907),
.Y(n_7845)
);

INVx1_ASAP7_75t_L g7846 ( 
.A(n_6706),
.Y(n_7846)
);

AND2x2_ASAP7_75t_L g7847 ( 
.A(n_7021),
.B(n_7302),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_6710),
.Y(n_7848)
);

INVx2_ASAP7_75t_L g7849 ( 
.A(n_7366),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_6710),
.Y(n_7850)
);

BUFx3_ASAP7_75t_L g7851 ( 
.A(n_7197),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_L g7852 ( 
.A(n_7593),
.B(n_6396),
.Y(n_7852)
);

INVx2_ASAP7_75t_L g7853 ( 
.A(n_7366),
.Y(n_7853)
);

INVx2_ASAP7_75t_L g7854 ( 
.A(n_7399),
.Y(n_7854)
);

INVx1_ASAP7_75t_L g7855 ( 
.A(n_6733),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_6733),
.Y(n_7856)
);

AOI22xp33_ASAP7_75t_SL g7857 ( 
.A1(n_7289),
.A2(n_6187),
.B1(n_6127),
.B2(n_6136),
.Y(n_7857)
);

BUFx2_ASAP7_75t_SL g7858 ( 
.A(n_6742),
.Y(n_7858)
);

INVx2_ASAP7_75t_L g7859 ( 
.A(n_7399),
.Y(n_7859)
);

INVx1_ASAP7_75t_L g7860 ( 
.A(n_6740),
.Y(n_7860)
);

OR2x2_ASAP7_75t_L g7861 ( 
.A(n_7630),
.B(n_6187),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_6740),
.Y(n_7862)
);

AND2x4_ASAP7_75t_L g7863 ( 
.A(n_7704),
.B(n_6985),
.Y(n_7863)
);

INVx1_ASAP7_75t_L g7864 ( 
.A(n_6751),
.Y(n_7864)
);

OAI22xp5_ASAP7_75t_L g7865 ( 
.A1(n_6699),
.A2(n_6352),
.B1(n_6050),
.B2(n_6382),
.Y(n_7865)
);

INVx2_ASAP7_75t_L g7866 ( 
.A(n_7399),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_6751),
.Y(n_7867)
);

AND2x2_ASAP7_75t_L g7868 ( 
.A(n_7021),
.B(n_6272),
.Y(n_7868)
);

INVx2_ASAP7_75t_L g7869 ( 
.A(n_7403),
.Y(n_7869)
);

INVx2_ASAP7_75t_L g7870 ( 
.A(n_7403),
.Y(n_7870)
);

AOI22xp5_ASAP7_75t_L g7871 ( 
.A1(n_6828),
.A2(n_6229),
.B1(n_6213),
.B2(n_6174),
.Y(n_7871)
);

INVx2_ASAP7_75t_L g7872 ( 
.A(n_7403),
.Y(n_7872)
);

NAND2x1p5_ASAP7_75t_L g7873 ( 
.A(n_6705),
.B(n_6324),
.Y(n_7873)
);

BUFx2_ASAP7_75t_SL g7874 ( 
.A(n_6742),
.Y(n_7874)
);

AOI22xp33_ASAP7_75t_L g7875 ( 
.A1(n_6678),
.A2(n_5825),
.B1(n_6223),
.B2(n_6136),
.Y(n_7875)
);

BUFx3_ASAP7_75t_L g7876 ( 
.A(n_7197),
.Y(n_7876)
);

NAND2xp5_ASAP7_75t_L g7877 ( 
.A(n_7593),
.B(n_6218),
.Y(n_7877)
);

INVx2_ASAP7_75t_L g7878 ( 
.A(n_7419),
.Y(n_7878)
);

NAND2xp5_ASAP7_75t_L g7879 ( 
.A(n_7054),
.B(n_6219),
.Y(n_7879)
);

OAI21xp5_ASAP7_75t_L g7880 ( 
.A1(n_7164),
.A2(n_6029),
.B(n_6224),
.Y(n_7880)
);

HB1xp67_ASAP7_75t_L g7881 ( 
.A(n_6996),
.Y(n_7881)
);

HB1xp67_ASAP7_75t_L g7882 ( 
.A(n_6996),
.Y(n_7882)
);

OR2x2_ASAP7_75t_L g7883 ( 
.A(n_7630),
.B(n_6537),
.Y(n_7883)
);

CKINVDCx9p33_ASAP7_75t_R g7884 ( 
.A(n_6923),
.Y(n_7884)
);

AOI22xp33_ASAP7_75t_L g7885 ( 
.A1(n_6678),
.A2(n_5825),
.B1(n_6223),
.B2(n_6664),
.Y(n_7885)
);

INVx4_ASAP7_75t_L g7886 ( 
.A(n_6713),
.Y(n_7886)
);

OR2x2_ASAP7_75t_L g7887 ( 
.A(n_7607),
.B(n_6537),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_6754),
.Y(n_7888)
);

INVx2_ASAP7_75t_L g7889 ( 
.A(n_7419),
.Y(n_7889)
);

AOI22xp33_ASAP7_75t_L g7890 ( 
.A1(n_6695),
.A2(n_5825),
.B1(n_6671),
.B2(n_6664),
.Y(n_7890)
);

INVx2_ASAP7_75t_L g7891 ( 
.A(n_7419),
.Y(n_7891)
);

AOI21x1_ASAP7_75t_L g7892 ( 
.A1(n_7498),
.A2(n_6859),
.B(n_6205),
.Y(n_7892)
);

BUFx2_ASAP7_75t_L g7893 ( 
.A(n_7289),
.Y(n_7893)
);

AND2x2_ASAP7_75t_L g7894 ( 
.A(n_7302),
.B(n_6272),
.Y(n_7894)
);

INVx3_ASAP7_75t_L g7895 ( 
.A(n_6949),
.Y(n_7895)
);

OAI21x1_ASAP7_75t_L g7896 ( 
.A1(n_7401),
.A2(n_6017),
.B(n_6531),
.Y(n_7896)
);

HB1xp67_ASAP7_75t_L g7897 ( 
.A(n_7423),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_6754),
.Y(n_7898)
);

AO21x2_ASAP7_75t_L g7899 ( 
.A1(n_7494),
.A2(n_5978),
.B(n_5927),
.Y(n_7899)
);

BUFx2_ASAP7_75t_L g7900 ( 
.A(n_7289),
.Y(n_7900)
);

INVx3_ASAP7_75t_L g7901 ( 
.A(n_7234),
.Y(n_7901)
);

HB1xp67_ASAP7_75t_L g7902 ( 
.A(n_7423),
.Y(n_7902)
);

AO21x2_ASAP7_75t_L g7903 ( 
.A1(n_7648),
.A2(n_7159),
.B(n_7490),
.Y(n_7903)
);

INVx3_ASAP7_75t_L g7904 ( 
.A(n_7234),
.Y(n_7904)
);

INVx2_ASAP7_75t_L g7905 ( 
.A(n_7425),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_6763),
.Y(n_7906)
);

INVx1_ASAP7_75t_L g7907 ( 
.A(n_6763),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_6766),
.Y(n_7908)
);

CKINVDCx6p67_ASAP7_75t_R g7909 ( 
.A(n_7245),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_6766),
.Y(n_7910)
);

AOI22xp33_ASAP7_75t_L g7911 ( 
.A1(n_6695),
.A2(n_5825),
.B1(n_6671),
.B2(n_5951),
.Y(n_7911)
);

INVx1_ASAP7_75t_L g7912 ( 
.A(n_6770),
.Y(n_7912)
);

INVx3_ASAP7_75t_L g7913 ( 
.A(n_7234),
.Y(n_7913)
);

INVx2_ASAP7_75t_L g7914 ( 
.A(n_7425),
.Y(n_7914)
);

OAI21x1_ASAP7_75t_L g7915 ( 
.A1(n_7401),
.A2(n_6017),
.B(n_6531),
.Y(n_7915)
);

AO21x2_ASAP7_75t_L g7916 ( 
.A1(n_7490),
.A2(n_5978),
.B(n_5927),
.Y(n_7916)
);

OR2x6_ASAP7_75t_L g7917 ( 
.A(n_6870),
.B(n_6635),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_6770),
.Y(n_7918)
);

INVx3_ASAP7_75t_L g7919 ( 
.A(n_7234),
.Y(n_7919)
);

AOI22xp5_ASAP7_75t_SL g7920 ( 
.A1(n_6805),
.A2(n_6378),
.B1(n_6427),
.B2(n_6319),
.Y(n_7920)
);

INVx3_ASAP7_75t_L g7921 ( 
.A(n_7234),
.Y(n_7921)
);

INVx2_ASAP7_75t_L g7922 ( 
.A(n_7425),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_6787),
.Y(n_7923)
);

INVx2_ASAP7_75t_L g7924 ( 
.A(n_7441),
.Y(n_7924)
);

BUFx3_ASAP7_75t_L g7925 ( 
.A(n_7276),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_6787),
.Y(n_7926)
);

BUFx6f_ASAP7_75t_SL g7927 ( 
.A(n_6713),
.Y(n_7927)
);

OA21x2_ASAP7_75t_L g7928 ( 
.A1(n_7193),
.A2(n_6017),
.B(n_6513),
.Y(n_7928)
);

OAI22xp5_ASAP7_75t_L g7929 ( 
.A1(n_6984),
.A2(n_6352),
.B1(n_6050),
.B2(n_6382),
.Y(n_7929)
);

AOI21x1_ASAP7_75t_L g7930 ( 
.A1(n_7498),
.A2(n_6205),
.B(n_6122),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_6792),
.Y(n_7931)
);

INVx2_ASAP7_75t_SL g7932 ( 
.A(n_6705),
.Y(n_7932)
);

HB1xp67_ASAP7_75t_L g7933 ( 
.A(n_7447),
.Y(n_7933)
);

INVx2_ASAP7_75t_L g7934 ( 
.A(n_7441),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_6792),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_6798),
.Y(n_7936)
);

INVx1_ASAP7_75t_L g7937 ( 
.A(n_6798),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_6800),
.Y(n_7938)
);

INVxp67_ASAP7_75t_L g7939 ( 
.A(n_6774),
.Y(n_7939)
);

INVx2_ASAP7_75t_L g7940 ( 
.A(n_7441),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_6800),
.Y(n_7941)
);

INVx2_ASAP7_75t_L g7942 ( 
.A(n_7460),
.Y(n_7942)
);

AND2x2_ASAP7_75t_L g7943 ( 
.A(n_7302),
.B(n_6272),
.Y(n_7943)
);

INVx1_ASAP7_75t_L g7944 ( 
.A(n_6803),
.Y(n_7944)
);

NAND2xp5_ASAP7_75t_L g7945 ( 
.A(n_7054),
.B(n_7446),
.Y(n_7945)
);

INVx4_ASAP7_75t_SL g7946 ( 
.A(n_6676),
.Y(n_7946)
);

INVx2_ASAP7_75t_L g7947 ( 
.A(n_7460),
.Y(n_7947)
);

INVx3_ASAP7_75t_L g7948 ( 
.A(n_7234),
.Y(n_7948)
);

HB1xp67_ASAP7_75t_L g7949 ( 
.A(n_7447),
.Y(n_7949)
);

INVx1_ASAP7_75t_L g7950 ( 
.A(n_6803),
.Y(n_7950)
);

OA21x2_ASAP7_75t_L g7951 ( 
.A1(n_7193),
.A2(n_6528),
.B(n_6513),
.Y(n_7951)
);

CKINVDCx20_ASAP7_75t_R g7952 ( 
.A(n_7033),
.Y(n_7952)
);

NAND2x1p5_ASAP7_75t_L g7953 ( 
.A(n_6705),
.B(n_6324),
.Y(n_7953)
);

NAND2xp5_ASAP7_75t_L g7954 ( 
.A(n_6869),
.B(n_6235),
.Y(n_7954)
);

INVx2_ASAP7_75t_SL g7955 ( 
.A(n_6705),
.Y(n_7955)
);

INVx2_ASAP7_75t_L g7956 ( 
.A(n_7460),
.Y(n_7956)
);

INVx2_ASAP7_75t_L g7957 ( 
.A(n_7496),
.Y(n_7957)
);

AND2x4_ASAP7_75t_L g7958 ( 
.A(n_7704),
.B(n_6456),
.Y(n_7958)
);

INVx1_ASAP7_75t_L g7959 ( 
.A(n_6814),
.Y(n_7959)
);

INVx1_ASAP7_75t_L g7960 ( 
.A(n_6814),
.Y(n_7960)
);

INVx1_ASAP7_75t_L g7961 ( 
.A(n_6816),
.Y(n_7961)
);

AND2x2_ASAP7_75t_L g7962 ( 
.A(n_7324),
.B(n_7342),
.Y(n_7962)
);

INVx1_ASAP7_75t_L g7963 ( 
.A(n_6816),
.Y(n_7963)
);

AOI21x1_ASAP7_75t_L g7964 ( 
.A1(n_6859),
.A2(n_6205),
.B(n_6122),
.Y(n_7964)
);

AND2x2_ASAP7_75t_L g7965 ( 
.A(n_7324),
.B(n_6651),
.Y(n_7965)
);

INVx1_ASAP7_75t_L g7966 ( 
.A(n_6820),
.Y(n_7966)
);

BUFx3_ASAP7_75t_L g7967 ( 
.A(n_7245),
.Y(n_7967)
);

AOI22xp33_ASAP7_75t_SL g7968 ( 
.A1(n_7289),
.A2(n_6246),
.B1(n_6235),
.B2(n_6250),
.Y(n_7968)
);

INVx3_ASAP7_75t_L g7969 ( 
.A(n_7295),
.Y(n_7969)
);

AOI22xp33_ASAP7_75t_L g7970 ( 
.A1(n_6895),
.A2(n_5951),
.B1(n_6151),
.B2(n_6147),
.Y(n_7970)
);

AO21x1_ASAP7_75t_SL g7971 ( 
.A1(n_6790),
.A2(n_6295),
.B(n_6172),
.Y(n_7971)
);

OAI21xp5_ASAP7_75t_L g7972 ( 
.A1(n_6959),
.A2(n_6246),
.B(n_6202),
.Y(n_7972)
);

INVx11_ASAP7_75t_L g7973 ( 
.A(n_6707),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_6820),
.Y(n_7974)
);

INVx1_ASAP7_75t_L g7975 ( 
.A(n_6821),
.Y(n_7975)
);

AND2x4_ASAP7_75t_L g7976 ( 
.A(n_7704),
.B(n_6456),
.Y(n_7976)
);

INVx6_ASAP7_75t_L g7977 ( 
.A(n_6707),
.Y(n_7977)
);

NAND2xp5_ASAP7_75t_L g7978 ( 
.A(n_6869),
.B(n_5792),
.Y(n_7978)
);

AOI22xp5_ASAP7_75t_L g7979 ( 
.A1(n_6679),
.A2(n_6435),
.B1(n_6418),
.B2(n_6313),
.Y(n_7979)
);

BUFx3_ASAP7_75t_L g7980 ( 
.A(n_7245),
.Y(n_7980)
);

INVx2_ASAP7_75t_L g7981 ( 
.A(n_7496),
.Y(n_7981)
);

OAI222xp33_ASAP7_75t_L g7982 ( 
.A1(n_7320),
.A2(n_6679),
.B1(n_7175),
.B2(n_6805),
.C1(n_7478),
.C2(n_6728),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_7496),
.Y(n_7983)
);

INVx1_ASAP7_75t_L g7984 ( 
.A(n_6821),
.Y(n_7984)
);

INVx1_ASAP7_75t_L g7985 ( 
.A(n_6827),
.Y(n_7985)
);

HB1xp67_ASAP7_75t_L g7986 ( 
.A(n_7586),
.Y(n_7986)
);

INVx2_ASAP7_75t_SL g7987 ( 
.A(n_6705),
.Y(n_7987)
);

INVx3_ASAP7_75t_L g7988 ( 
.A(n_7295),
.Y(n_7988)
);

INVx1_ASAP7_75t_L g7989 ( 
.A(n_6827),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_6829),
.Y(n_7990)
);

OAI21x1_ASAP7_75t_L g7991 ( 
.A1(n_7325),
.A2(n_6558),
.B(n_6550),
.Y(n_7991)
);

BUFx2_ASAP7_75t_L g7992 ( 
.A(n_7303),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_6829),
.Y(n_7993)
);

INVx1_ASAP7_75t_L g7994 ( 
.A(n_6832),
.Y(n_7994)
);

AND2x2_ASAP7_75t_L g7995 ( 
.A(n_7324),
.B(n_6651),
.Y(n_7995)
);

AOI22xp33_ASAP7_75t_L g7996 ( 
.A1(n_7478),
.A2(n_5951),
.B1(n_6151),
.B2(n_6147),
.Y(n_7996)
);

HB1xp67_ASAP7_75t_L g7997 ( 
.A(n_7586),
.Y(n_7997)
);

INVx1_ASAP7_75t_L g7998 ( 
.A(n_6832),
.Y(n_7998)
);

INVx2_ASAP7_75t_L g7999 ( 
.A(n_7545),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_6845),
.Y(n_8000)
);

AOI22xp33_ASAP7_75t_L g8001 ( 
.A1(n_6690),
.A2(n_5951),
.B1(n_6167),
.B2(n_6435),
.Y(n_8001)
);

INVx2_ASAP7_75t_L g8002 ( 
.A(n_7545),
.Y(n_8002)
);

INVx1_ASAP7_75t_L g8003 ( 
.A(n_6845),
.Y(n_8003)
);

INVx3_ASAP7_75t_L g8004 ( 
.A(n_7295),
.Y(n_8004)
);

HB1xp67_ASAP7_75t_L g8005 ( 
.A(n_7676),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_6847),
.Y(n_8006)
);

NAND2x1_ASAP7_75t_L g8007 ( 
.A(n_7587),
.B(n_6672),
.Y(n_8007)
);

INVx2_ASAP7_75t_L g8008 ( 
.A(n_7545),
.Y(n_8008)
);

INVx1_ASAP7_75t_L g8009 ( 
.A(n_6847),
.Y(n_8009)
);

INVx1_ASAP7_75t_L g8010 ( 
.A(n_6848),
.Y(n_8010)
);

INVx2_ASAP7_75t_L g8011 ( 
.A(n_7547),
.Y(n_8011)
);

BUFx4f_ASAP7_75t_L g8012 ( 
.A(n_6776),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_6848),
.Y(n_8013)
);

INVx1_ASAP7_75t_L g8014 ( 
.A(n_6852),
.Y(n_8014)
);

AOI22xp33_ASAP7_75t_L g8015 ( 
.A1(n_6690),
.A2(n_5951),
.B1(n_6167),
.B2(n_5824),
.Y(n_8015)
);

BUFx3_ASAP7_75t_L g8016 ( 
.A(n_7272),
.Y(n_8016)
);

INVx2_ASAP7_75t_SL g8017 ( 
.A(n_7002),
.Y(n_8017)
);

INVx2_ASAP7_75t_L g8018 ( 
.A(n_7547),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_6852),
.Y(n_8019)
);

AO21x2_ASAP7_75t_L g8020 ( 
.A1(n_7700),
.A2(n_5917),
.B(n_5854),
.Y(n_8020)
);

INVx3_ASAP7_75t_L g8021 ( 
.A(n_7295),
.Y(n_8021)
);

NAND2x1_ASAP7_75t_L g8022 ( 
.A(n_7587),
.B(n_6672),
.Y(n_8022)
);

INVx2_ASAP7_75t_L g8023 ( 
.A(n_7547),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_6862),
.Y(n_8024)
);

BUFx2_ASAP7_75t_L g8025 ( 
.A(n_7303),
.Y(n_8025)
);

INVx2_ASAP7_75t_L g8026 ( 
.A(n_7562),
.Y(n_8026)
);

BUFx2_ASAP7_75t_L g8027 ( 
.A(n_7303),
.Y(n_8027)
);

NAND2xp5_ASAP7_75t_L g8028 ( 
.A(n_7606),
.B(n_5792),
.Y(n_8028)
);

INVx2_ASAP7_75t_L g8029 ( 
.A(n_7562),
.Y(n_8029)
);

BUFx2_ASAP7_75t_L g8030 ( 
.A(n_7303),
.Y(n_8030)
);

HB1xp67_ASAP7_75t_L g8031 ( 
.A(n_7676),
.Y(n_8031)
);

INVx1_ASAP7_75t_L g8032 ( 
.A(n_6862),
.Y(n_8032)
);

AO21x1_ASAP7_75t_SL g8033 ( 
.A1(n_6693),
.A2(n_5892),
.B(n_6283),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_6863),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_6863),
.Y(n_8035)
);

OAI21x1_ASAP7_75t_L g8036 ( 
.A1(n_7325),
.A2(n_6558),
.B(n_6550),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_6872),
.Y(n_8037)
);

BUFx6f_ASAP7_75t_L g8038 ( 
.A(n_6700),
.Y(n_8038)
);

AO21x2_ASAP7_75t_L g8039 ( 
.A1(n_7700),
.A2(n_5917),
.B(n_5854),
.Y(n_8039)
);

BUFx12f_ASAP7_75t_L g8040 ( 
.A(n_6964),
.Y(n_8040)
);

NOR2x1_ASAP7_75t_R g8041 ( 
.A(n_7077),
.B(n_5985),
.Y(n_8041)
);

BUFx2_ASAP7_75t_L g8042 ( 
.A(n_7466),
.Y(n_8042)
);

AOI22xp33_ASAP7_75t_SL g8043 ( 
.A1(n_7735),
.A2(n_6250),
.B1(n_6183),
.B2(n_6188),
.Y(n_8043)
);

AND2x2_ASAP7_75t_L g8044 ( 
.A(n_7342),
.B(n_6651),
.Y(n_8044)
);

INVx3_ASAP7_75t_L g8045 ( 
.A(n_7295),
.Y(n_8045)
);

OAI21x1_ASAP7_75t_L g8046 ( 
.A1(n_7325),
.A2(n_6566),
.B(n_6565),
.Y(n_8046)
);

INVx1_ASAP7_75t_L g8047 ( 
.A(n_6872),
.Y(n_8047)
);

BUFx3_ASAP7_75t_L g8048 ( 
.A(n_7272),
.Y(n_8048)
);

NAND2xp5_ASAP7_75t_L g8049 ( 
.A(n_7606),
.B(n_6307),
.Y(n_8049)
);

BUFx2_ASAP7_75t_L g8050 ( 
.A(n_7466),
.Y(n_8050)
);

AND2x4_ASAP7_75t_L g8051 ( 
.A(n_7704),
.B(n_6456),
.Y(n_8051)
);

INVx1_ASAP7_75t_L g8052 ( 
.A(n_6875),
.Y(n_8052)
);

INVx2_ASAP7_75t_L g8053 ( 
.A(n_7562),
.Y(n_8053)
);

INVx1_ASAP7_75t_L g8054 ( 
.A(n_6875),
.Y(n_8054)
);

AOI221xp5_ASAP7_75t_L g8055 ( 
.A1(n_6830),
.A2(n_6304),
.B1(n_6299),
.B2(n_6551),
.C(n_6546),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_6877),
.Y(n_8056)
);

INVx3_ASAP7_75t_L g8057 ( 
.A(n_7295),
.Y(n_8057)
);

INVx6_ASAP7_75t_L g8058 ( 
.A(n_6707),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_7592),
.Y(n_8059)
);

BUFx6f_ASAP7_75t_L g8060 ( 
.A(n_6700),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_6877),
.Y(n_8061)
);

INVx1_ASAP7_75t_L g8062 ( 
.A(n_6885),
.Y(n_8062)
);

INVx2_ASAP7_75t_SL g8063 ( 
.A(n_7002),
.Y(n_8063)
);

INVx1_ASAP7_75t_L g8064 ( 
.A(n_6885),
.Y(n_8064)
);

INVx1_ASAP7_75t_L g8065 ( 
.A(n_6888),
.Y(n_8065)
);

NAND2x1_ASAP7_75t_L g8066 ( 
.A(n_7587),
.B(n_6672),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_6888),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_6891),
.Y(n_8068)
);

INVx2_ASAP7_75t_L g8069 ( 
.A(n_7592),
.Y(n_8069)
);

INVx2_ASAP7_75t_L g8070 ( 
.A(n_7592),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_6891),
.Y(n_8071)
);

HB1xp67_ASAP7_75t_L g8072 ( 
.A(n_6892),
.Y(n_8072)
);

INVx1_ASAP7_75t_L g8073 ( 
.A(n_6892),
.Y(n_8073)
);

INVx2_ASAP7_75t_L g8074 ( 
.A(n_7595),
.Y(n_8074)
);

HB1xp67_ASAP7_75t_L g8075 ( 
.A(n_6899),
.Y(n_8075)
);

INVx4_ASAP7_75t_L g8076 ( 
.A(n_6713),
.Y(n_8076)
);

INVx4_ASAP7_75t_L g8077 ( 
.A(n_6738),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_6899),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_6914),
.Y(n_8079)
);

INVx2_ASAP7_75t_L g8080 ( 
.A(n_7595),
.Y(n_8080)
);

OAI21x1_ASAP7_75t_L g8081 ( 
.A1(n_7325),
.A2(n_6566),
.B(n_6565),
.Y(n_8081)
);

INVx1_ASAP7_75t_L g8082 ( 
.A(n_6914),
.Y(n_8082)
);

HB1xp67_ASAP7_75t_L g8083 ( 
.A(n_6933),
.Y(n_8083)
);

INVx2_ASAP7_75t_L g8084 ( 
.A(n_7595),
.Y(n_8084)
);

AOI22xp33_ASAP7_75t_L g8085 ( 
.A1(n_6717),
.A2(n_5951),
.B1(n_5824),
.B2(n_5906),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_6933),
.Y(n_8086)
);

BUFx8_ASAP7_75t_SL g8087 ( 
.A(n_6680),
.Y(n_8087)
);

INVx2_ASAP7_75t_L g8088 ( 
.A(n_7603),
.Y(n_8088)
);

INVx2_ASAP7_75t_L g8089 ( 
.A(n_7603),
.Y(n_8089)
);

OAI21x1_ASAP7_75t_L g8090 ( 
.A1(n_7376),
.A2(n_6582),
.B(n_6574),
.Y(n_8090)
);

OAI21x1_ASAP7_75t_L g8091 ( 
.A1(n_7376),
.A2(n_6582),
.B(n_6574),
.Y(n_8091)
);

INVx1_ASAP7_75t_L g8092 ( 
.A(n_6942),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_6942),
.Y(n_8093)
);

AOI22xp33_ASAP7_75t_SL g8094 ( 
.A1(n_7466),
.A2(n_6175),
.B1(n_6188),
.B2(n_6183),
.Y(n_8094)
);

INVx2_ASAP7_75t_SL g8095 ( 
.A(n_7002),
.Y(n_8095)
);

HB1xp67_ASAP7_75t_L g8096 ( 
.A(n_6943),
.Y(n_8096)
);

INVx2_ASAP7_75t_L g8097 ( 
.A(n_7603),
.Y(n_8097)
);

INVx1_ASAP7_75t_L g8098 ( 
.A(n_6943),
.Y(n_8098)
);

NAND2x1_ASAP7_75t_L g8099 ( 
.A(n_7587),
.B(n_6672),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_6948),
.Y(n_8100)
);

INVx2_ASAP7_75t_SL g8101 ( 
.A(n_7002),
.Y(n_8101)
);

INVx1_ASAP7_75t_L g8102 ( 
.A(n_6948),
.Y(n_8102)
);

AO21x2_ASAP7_75t_L g8103 ( 
.A1(n_7355),
.A2(n_5845),
.B(n_6528),
.Y(n_8103)
);

BUFx2_ASAP7_75t_L g8104 ( 
.A(n_7466),
.Y(n_8104)
);

INVx2_ASAP7_75t_SL g8105 ( 
.A(n_7002),
.Y(n_8105)
);

NOR2xp33_ASAP7_75t_L g8106 ( 
.A(n_6712),
.B(n_6002),
.Y(n_8106)
);

INVx3_ASAP7_75t_L g8107 ( 
.A(n_7431),
.Y(n_8107)
);

AOI22xp33_ASAP7_75t_L g8108 ( 
.A1(n_6717),
.A2(n_5906),
.B1(n_6418),
.B2(n_6540),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7604),
.Y(n_8109)
);

BUFx3_ASAP7_75t_L g8110 ( 
.A(n_7272),
.Y(n_8110)
);

BUFx2_ASAP7_75t_L g8111 ( 
.A(n_7488),
.Y(n_8111)
);

AOI21x1_ASAP7_75t_L g8112 ( 
.A1(n_7636),
.A2(n_6212),
.B(n_5955),
.Y(n_8112)
);

INVx3_ASAP7_75t_L g8113 ( 
.A(n_7431),
.Y(n_8113)
);

INVx1_ASAP7_75t_L g8114 ( 
.A(n_6953),
.Y(n_8114)
);

INVx1_ASAP7_75t_L g8115 ( 
.A(n_6953),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7604),
.Y(n_8116)
);

INVx3_ASAP7_75t_L g8117 ( 
.A(n_7431),
.Y(n_8117)
);

AND2x2_ASAP7_75t_L g8118 ( 
.A(n_7342),
.B(n_6545),
.Y(n_8118)
);

BUFx6f_ASAP7_75t_L g8119 ( 
.A(n_6700),
.Y(n_8119)
);

INVx2_ASAP7_75t_L g8120 ( 
.A(n_7604),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_6957),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_6957),
.Y(n_8122)
);

INVx2_ASAP7_75t_L g8123 ( 
.A(n_7618),
.Y(n_8123)
);

AND2x2_ASAP7_75t_L g8124 ( 
.A(n_6925),
.B(n_6600),
.Y(n_8124)
);

INVx1_ASAP7_75t_L g8125 ( 
.A(n_6972),
.Y(n_8125)
);

INVx2_ASAP7_75t_SL g8126 ( 
.A(n_7002),
.Y(n_8126)
);

OR2x6_ASAP7_75t_L g8127 ( 
.A(n_7431),
.B(n_7177),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_6972),
.Y(n_8128)
);

AND2x2_ASAP7_75t_L g8129 ( 
.A(n_6925),
.B(n_6600),
.Y(n_8129)
);

INVx2_ASAP7_75t_L g8130 ( 
.A(n_7618),
.Y(n_8130)
);

OAI21x1_ASAP7_75t_SL g8131 ( 
.A1(n_7745),
.A2(n_6580),
.B(n_6287),
.Y(n_8131)
);

INVx2_ASAP7_75t_L g8132 ( 
.A(n_7618),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_6979),
.Y(n_8133)
);

INVx1_ASAP7_75t_L g8134 ( 
.A(n_6979),
.Y(n_8134)
);

CKINVDCx8_ASAP7_75t_R g8135 ( 
.A(n_7207),
.Y(n_8135)
);

AO21x1_ASAP7_75t_SL g8136 ( 
.A1(n_6693),
.A2(n_5892),
.B(n_6283),
.Y(n_8136)
);

INVxp67_ASAP7_75t_L g8137 ( 
.A(n_6774),
.Y(n_8137)
);

NOR2xp33_ASAP7_75t_L g8138 ( 
.A(n_6712),
.B(n_6002),
.Y(n_8138)
);

INVxp33_ASAP7_75t_L g8139 ( 
.A(n_6718),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_6980),
.Y(n_8140)
);

AND2x2_ASAP7_75t_L g8141 ( 
.A(n_6925),
.B(n_6600),
.Y(n_8141)
);

AOI22xp33_ASAP7_75t_L g8142 ( 
.A1(n_7320),
.A2(n_5906),
.B1(n_6540),
.B2(n_5892),
.Y(n_8142)
);

INVx2_ASAP7_75t_L g8143 ( 
.A(n_7626),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_6980),
.Y(n_8144)
);

BUFx2_ASAP7_75t_SL g8145 ( 
.A(n_6742),
.Y(n_8145)
);

HB1xp67_ASAP7_75t_L g8146 ( 
.A(n_6994),
.Y(n_8146)
);

BUFx3_ASAP7_75t_L g8147 ( 
.A(n_7276),
.Y(n_8147)
);

OAI21x1_ASAP7_75t_L g8148 ( 
.A1(n_7376),
.A2(n_6607),
.B(n_6593),
.Y(n_8148)
);

NOR2xp33_ASAP7_75t_L g8149 ( 
.A(n_6743),
.B(n_6525),
.Y(n_8149)
);

INVx2_ASAP7_75t_SL g8150 ( 
.A(n_7002),
.Y(n_8150)
);

BUFx3_ASAP7_75t_L g8151 ( 
.A(n_7276),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_6994),
.Y(n_8152)
);

AND2x2_ASAP7_75t_L g8153 ( 
.A(n_6946),
.B(n_6630),
.Y(n_8153)
);

INVx2_ASAP7_75t_L g8154 ( 
.A(n_7626),
.Y(n_8154)
);

INVx2_ASAP7_75t_L g8155 ( 
.A(n_7626),
.Y(n_8155)
);

INVx2_ASAP7_75t_L g8156 ( 
.A(n_7631),
.Y(n_8156)
);

HB1xp67_ASAP7_75t_SL g8157 ( 
.A(n_6707),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_7007),
.Y(n_8158)
);

OAI22xp5_ASAP7_75t_L g8159 ( 
.A1(n_6728),
.A2(n_6753),
.B1(n_6801),
.B2(n_7175),
.Y(n_8159)
);

INVx2_ASAP7_75t_L g8160 ( 
.A(n_7631),
.Y(n_8160)
);

INVx2_ASAP7_75t_L g8161 ( 
.A(n_7631),
.Y(n_8161)
);

INVx3_ASAP7_75t_L g8162 ( 
.A(n_7431),
.Y(n_8162)
);

CKINVDCx20_ASAP7_75t_R g8163 ( 
.A(n_6823),
.Y(n_8163)
);

INVx2_ASAP7_75t_L g8164 ( 
.A(n_7638),
.Y(n_8164)
);

AND2x2_ASAP7_75t_L g8165 ( 
.A(n_6946),
.B(n_6630),
.Y(n_8165)
);

INVx1_ASAP7_75t_SL g8166 ( 
.A(n_7467),
.Y(n_8166)
);

OAI21x1_ASAP7_75t_L g8167 ( 
.A1(n_7376),
.A2(n_6607),
.B(n_6593),
.Y(n_8167)
);

INVx2_ASAP7_75t_L g8168 ( 
.A(n_7638),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7007),
.Y(n_8169)
);

AOI21xp33_ASAP7_75t_L g8170 ( 
.A1(n_7177),
.A2(n_5913),
.B(n_6108),
.Y(n_8170)
);

CKINVDCx12_ASAP7_75t_R g8171 ( 
.A(n_6718),
.Y(n_8171)
);

INVx2_ASAP7_75t_L g8172 ( 
.A(n_7638),
.Y(n_8172)
);

INVx3_ASAP7_75t_L g8173 ( 
.A(n_7431),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_7015),
.Y(n_8174)
);

BUFx2_ASAP7_75t_SL g8175 ( 
.A(n_6682),
.Y(n_8175)
);

INVx2_ASAP7_75t_L g8176 ( 
.A(n_7652),
.Y(n_8176)
);

INVx3_ASAP7_75t_L g8177 ( 
.A(n_6765),
.Y(n_8177)
);

BUFx3_ASAP7_75t_L g8178 ( 
.A(n_6771),
.Y(n_8178)
);

AND2x2_ASAP7_75t_L g8179 ( 
.A(n_6946),
.B(n_6630),
.Y(n_8179)
);

INVx2_ASAP7_75t_SL g8180 ( 
.A(n_7043),
.Y(n_8180)
);

OAI21xp5_ASAP7_75t_L g8181 ( 
.A1(n_6830),
.A2(n_6202),
.B(n_6121),
.Y(n_8181)
);

INVx2_ASAP7_75t_L g8182 ( 
.A(n_7652),
.Y(n_8182)
);

INVx2_ASAP7_75t_L g8183 ( 
.A(n_7652),
.Y(n_8183)
);

AND2x2_ASAP7_75t_L g8184 ( 
.A(n_6990),
.B(n_7006),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7015),
.Y(n_8185)
);

AO21x1_ASAP7_75t_L g8186 ( 
.A1(n_7472),
.A2(n_6839),
.B(n_7745),
.Y(n_8186)
);

HB1xp67_ASAP7_75t_L g8187 ( 
.A(n_7025),
.Y(n_8187)
);

INVx2_ASAP7_75t_L g8188 ( 
.A(n_7656),
.Y(n_8188)
);

INVx2_ASAP7_75t_L g8189 ( 
.A(n_7656),
.Y(n_8189)
);

AOI22xp33_ASAP7_75t_SL g8190 ( 
.A1(n_7488),
.A2(n_6175),
.B1(n_6025),
.B2(n_6540),
.Y(n_8190)
);

OR2x6_ASAP7_75t_L g8191 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8191)
);

INVx2_ASAP7_75t_L g8192 ( 
.A(n_7656),
.Y(n_8192)
);

INVx1_ASAP7_75t_SL g8193 ( 
.A(n_7467),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7025),
.Y(n_8194)
);

INVx2_ASAP7_75t_L g8195 ( 
.A(n_7673),
.Y(n_8195)
);

OAI22xp33_ASAP7_75t_L g8196 ( 
.A1(n_6839),
.A2(n_6313),
.B1(n_6284),
.B2(n_6343),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_7027),
.Y(n_8197)
);

AND2x2_ASAP7_75t_L g8198 ( 
.A(n_6990),
.B(n_6031),
.Y(n_8198)
);

AND2x2_ASAP7_75t_L g8199 ( 
.A(n_6990),
.B(n_6031),
.Y(n_8199)
);

AND2x2_ASAP7_75t_L g8200 ( 
.A(n_7006),
.B(n_6031),
.Y(n_8200)
);

INVx2_ASAP7_75t_L g8201 ( 
.A(n_7673),
.Y(n_8201)
);

BUFx3_ASAP7_75t_L g8202 ( 
.A(n_6771),
.Y(n_8202)
);

INVx3_ASAP7_75t_L g8203 ( 
.A(n_6765),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7027),
.Y(n_8204)
);

INVx1_ASAP7_75t_L g8205 ( 
.A(n_7048),
.Y(n_8205)
);

OAI21x1_ASAP7_75t_L g8206 ( 
.A1(n_7509),
.A2(n_6616),
.B(n_6613),
.Y(n_8206)
);

OR2x6_ASAP7_75t_L g8207 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_7673),
.Y(n_8208)
);

OA21x2_ASAP7_75t_L g8209 ( 
.A1(n_7599),
.A2(n_6661),
.B(n_6447),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_7048),
.Y(n_8210)
);

AND2x2_ASAP7_75t_L g8211 ( 
.A(n_7006),
.B(n_6031),
.Y(n_8211)
);

BUFx2_ASAP7_75t_R g8212 ( 
.A(n_6799),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_7066),
.Y(n_8213)
);

OAI21x1_ASAP7_75t_L g8214 ( 
.A1(n_7509),
.A2(n_6616),
.B(n_6613),
.Y(n_8214)
);

INVx2_ASAP7_75t_L g8215 ( 
.A(n_7675),
.Y(n_8215)
);

OA21x2_ASAP7_75t_L g8216 ( 
.A1(n_7599),
.A2(n_6661),
.B(n_6447),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_7066),
.Y(n_8217)
);

AND2x2_ASAP7_75t_L g8218 ( 
.A(n_7029),
.B(n_6031),
.Y(n_8218)
);

INVx3_ASAP7_75t_L g8219 ( 
.A(n_6765),
.Y(n_8219)
);

INVx2_ASAP7_75t_L g8220 ( 
.A(n_7675),
.Y(n_8220)
);

AND2x4_ASAP7_75t_SL g8221 ( 
.A(n_7150),
.B(n_5985),
.Y(n_8221)
);

INVx3_ASAP7_75t_L g8222 ( 
.A(n_6765),
.Y(n_8222)
);

OAI21x1_ASAP7_75t_L g8223 ( 
.A1(n_7509),
.A2(n_6572),
.B(n_5957),
.Y(n_8223)
);

OAI22xp33_ASAP7_75t_L g8224 ( 
.A1(n_7060),
.A2(n_6284),
.B1(n_6343),
.B2(n_5986),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7069),
.Y(n_8225)
);

OAI22xp33_ASAP7_75t_L g8226 ( 
.A1(n_7060),
.A2(n_5986),
.B1(n_6298),
.B2(n_6319),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7069),
.Y(n_8227)
);

INVx3_ASAP7_75t_L g8228 ( 
.A(n_6765),
.Y(n_8228)
);

AOI22xp33_ASAP7_75t_SL g8229 ( 
.A1(n_7488),
.A2(n_6025),
.B1(n_6540),
.B2(n_6503),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7078),
.Y(n_8230)
);

BUFx2_ASAP7_75t_L g8231 ( 
.A(n_7488),
.Y(n_8231)
);

INVx2_ASAP7_75t_L g8232 ( 
.A(n_7675),
.Y(n_8232)
);

INVx3_ASAP7_75t_L g8233 ( 
.A(n_6765),
.Y(n_8233)
);

INVx2_ASAP7_75t_L g8234 ( 
.A(n_7685),
.Y(n_8234)
);

NAND2x1p5_ASAP7_75t_L g8235 ( 
.A(n_7043),
.B(n_5931),
.Y(n_8235)
);

INVx3_ASAP7_75t_L g8236 ( 
.A(n_6765),
.Y(n_8236)
);

INVx1_ASAP7_75t_L g8237 ( 
.A(n_7078),
.Y(n_8237)
);

AOI22xp33_ASAP7_75t_SL g8238 ( 
.A1(n_7622),
.A2(n_6540),
.B1(n_6503),
.B2(n_6378),
.Y(n_8238)
);

INVx3_ASAP7_75t_L g8239 ( 
.A(n_6786),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_7085),
.Y(n_8240)
);

OR2x6_ASAP7_75t_L g8241 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8241)
);

INVx1_ASAP7_75t_SL g8242 ( 
.A(n_6894),
.Y(n_8242)
);

INVx1_ASAP7_75t_L g8243 ( 
.A(n_7085),
.Y(n_8243)
);

INVx2_ASAP7_75t_L g8244 ( 
.A(n_7685),
.Y(n_8244)
);

BUFx12f_ASAP7_75t_L g8245 ( 
.A(n_7102),
.Y(n_8245)
);

CKINVDCx16_ASAP7_75t_R g8246 ( 
.A(n_7207),
.Y(n_8246)
);

INVx1_ASAP7_75t_L g8247 ( 
.A(n_7097),
.Y(n_8247)
);

BUFx2_ASAP7_75t_L g8248 ( 
.A(n_7622),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_7097),
.Y(n_8249)
);

INVx1_ASAP7_75t_L g8250 ( 
.A(n_7098),
.Y(n_8250)
);

INVx2_ASAP7_75t_L g8251 ( 
.A(n_7685),
.Y(n_8251)
);

INVx6_ASAP7_75t_L g8252 ( 
.A(n_6771),
.Y(n_8252)
);

NAND2xp5_ASAP7_75t_L g8253 ( 
.A(n_7701),
.B(n_6307),
.Y(n_8253)
);

INVx2_ASAP7_75t_L g8254 ( 
.A(n_7696),
.Y(n_8254)
);

OR2x2_ASAP7_75t_L g8255 ( 
.A(n_7607),
.B(n_6546),
.Y(n_8255)
);

INVx3_ASAP7_75t_L g8256 ( 
.A(n_6786),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7098),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7103),
.Y(n_8258)
);

INVx2_ASAP7_75t_L g8259 ( 
.A(n_7696),
.Y(n_8259)
);

NAND2xp5_ASAP7_75t_L g8260 ( 
.A(n_7701),
.B(n_6314),
.Y(n_8260)
);

OA21x2_ASAP7_75t_L g8261 ( 
.A1(n_7654),
.A2(n_6445),
.B(n_6510),
.Y(n_8261)
);

HB1xp67_ASAP7_75t_L g8262 ( 
.A(n_7103),
.Y(n_8262)
);

INVx3_ASAP7_75t_L g8263 ( 
.A(n_6786),
.Y(n_8263)
);

INVx2_ASAP7_75t_L g8264 ( 
.A(n_7696),
.Y(n_8264)
);

AND2x2_ASAP7_75t_L g8265 ( 
.A(n_7029),
.B(n_7151),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_7104),
.Y(n_8266)
);

INVx1_ASAP7_75t_L g8267 ( 
.A(n_7104),
.Y(n_8267)
);

INVx1_ASAP7_75t_L g8268 ( 
.A(n_7125),
.Y(n_8268)
);

HB1xp67_ASAP7_75t_L g8269 ( 
.A(n_7125),
.Y(n_8269)
);

INVx2_ASAP7_75t_L g8270 ( 
.A(n_7749),
.Y(n_8270)
);

AND2x2_ASAP7_75t_L g8271 ( 
.A(n_7029),
.B(n_6031),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_7739),
.B(n_6314),
.Y(n_8272)
);

AOI22xp33_ASAP7_75t_SL g8273 ( 
.A1(n_7622),
.A2(n_6540),
.B1(n_6427),
.B2(n_6248),
.Y(n_8273)
);

INVx4_ASAP7_75t_L g8274 ( 
.A(n_6738),
.Y(n_8274)
);

OR2x2_ASAP7_75t_L g8275 ( 
.A(n_7635),
.B(n_6551),
.Y(n_8275)
);

HB1xp67_ASAP7_75t_L g8276 ( 
.A(n_7139),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_7139),
.Y(n_8277)
);

BUFx3_ASAP7_75t_L g8278 ( 
.A(n_6771),
.Y(n_8278)
);

HB1xp67_ASAP7_75t_L g8279 ( 
.A(n_7154),
.Y(n_8279)
);

BUFx6f_ASAP7_75t_L g8280 ( 
.A(n_6700),
.Y(n_8280)
);

AO21x2_ASAP7_75t_L g8281 ( 
.A1(n_7355),
.A2(n_5845),
.B(n_6510),
.Y(n_8281)
);

INVx2_ASAP7_75t_SL g8282 ( 
.A(n_7043),
.Y(n_8282)
);

INVx2_ASAP7_75t_L g8283 ( 
.A(n_7749),
.Y(n_8283)
);

AND2x2_ASAP7_75t_L g8284 ( 
.A(n_7151),
.B(n_6031),
.Y(n_8284)
);

CKINVDCx5p33_ASAP7_75t_R g8285 ( 
.A(n_6835),
.Y(n_8285)
);

INVx2_ASAP7_75t_L g8286 ( 
.A(n_7749),
.Y(n_8286)
);

INVx2_ASAP7_75t_L g8287 ( 
.A(n_7762),
.Y(n_8287)
);

AOI222xp33_ASAP7_75t_L g8288 ( 
.A1(n_6807),
.A2(n_6279),
.B1(n_6248),
.B2(n_6108),
.C1(n_5913),
.C2(n_6374),
.Y(n_8288)
);

NAND2xp5_ASAP7_75t_L g8289 ( 
.A(n_7739),
.B(n_6353),
.Y(n_8289)
);

OAI21xp5_ASAP7_75t_L g8290 ( 
.A1(n_7472),
.A2(n_6093),
.B(n_6077),
.Y(n_8290)
);

INVx2_ASAP7_75t_L g8291 ( 
.A(n_7762),
.Y(n_8291)
);

BUFx12f_ASAP7_75t_L g8292 ( 
.A(n_7106),
.Y(n_8292)
);

AOI22xp33_ASAP7_75t_L g8293 ( 
.A1(n_7264),
.A2(n_5906),
.B1(n_6649),
.B2(n_6164),
.Y(n_8293)
);

BUFx3_ASAP7_75t_L g8294 ( 
.A(n_6781),
.Y(n_8294)
);

AOI22xp33_ASAP7_75t_L g8295 ( 
.A1(n_7264),
.A2(n_5906),
.B1(n_6649),
.B2(n_6164),
.Y(n_8295)
);

INVx2_ASAP7_75t_L g8296 ( 
.A(n_7762),
.Y(n_8296)
);

HB1xp67_ASAP7_75t_L g8297 ( 
.A(n_7154),
.Y(n_8297)
);

AOI22xp33_ASAP7_75t_SL g8298 ( 
.A1(n_7622),
.A2(n_6502),
.B1(n_6654),
.B2(n_6394),
.Y(n_8298)
);

INVx2_ASAP7_75t_L g8299 ( 
.A(n_7768),
.Y(n_8299)
);

NAND2xp5_ASAP7_75t_L g8300 ( 
.A(n_7743),
.B(n_6353),
.Y(n_8300)
);

OAI21xp5_ASAP7_75t_L g8301 ( 
.A1(n_7195),
.A2(n_6093),
.B(n_6077),
.Y(n_8301)
);

INVx2_ASAP7_75t_L g8302 ( 
.A(n_7768),
.Y(n_8302)
);

BUFx3_ASAP7_75t_L g8303 ( 
.A(n_6781),
.Y(n_8303)
);

INVx3_ASAP7_75t_L g8304 ( 
.A(n_6786),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_7165),
.Y(n_8305)
);

INVx3_ASAP7_75t_L g8306 ( 
.A(n_6786),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_7165),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_7173),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_7173),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7174),
.Y(n_8310)
);

INVx2_ASAP7_75t_L g8311 ( 
.A(n_7768),
.Y(n_8311)
);

OA21x2_ASAP7_75t_L g8312 ( 
.A1(n_7654),
.A2(n_6445),
.B(n_6251),
.Y(n_8312)
);

OAI21x1_ASAP7_75t_L g8313 ( 
.A1(n_7509),
.A2(n_6572),
.B(n_5957),
.Y(n_8313)
);

INVx1_ASAP7_75t_L g8314 ( 
.A(n_7174),
.Y(n_8314)
);

NAND2xp5_ASAP7_75t_L g8315 ( 
.A(n_7743),
.B(n_6562),
.Y(n_8315)
);

INVx2_ASAP7_75t_L g8316 ( 
.A(n_7771),
.Y(n_8316)
);

BUFx2_ASAP7_75t_L g8317 ( 
.A(n_7735),
.Y(n_8317)
);

INVx2_ASAP7_75t_L g8318 ( 
.A(n_7771),
.Y(n_8318)
);

INVx1_ASAP7_75t_L g8319 ( 
.A(n_7180),
.Y(n_8319)
);

INVx1_ASAP7_75t_L g8320 ( 
.A(n_7180),
.Y(n_8320)
);

AOI22xp33_ASAP7_75t_L g8321 ( 
.A1(n_6734),
.A2(n_5906),
.B1(n_6279),
.B2(n_6194),
.Y(n_8321)
);

INVx2_ASAP7_75t_L g8322 ( 
.A(n_7771),
.Y(n_8322)
);

INVx3_ASAP7_75t_L g8323 ( 
.A(n_6786),
.Y(n_8323)
);

BUFx10_ASAP7_75t_L g8324 ( 
.A(n_6676),
.Y(n_8324)
);

INVx2_ASAP7_75t_L g8325 ( 
.A(n_6701),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7181),
.Y(n_8326)
);

AOI22xp33_ASAP7_75t_L g8327 ( 
.A1(n_6734),
.A2(n_6194),
.B1(n_6133),
.B2(n_6020),
.Y(n_8327)
);

INVx2_ASAP7_75t_L g8328 ( 
.A(n_6701),
.Y(n_8328)
);

INVx1_ASAP7_75t_L g8329 ( 
.A(n_7181),
.Y(n_8329)
);

OAI22xp33_ASAP7_75t_L g8330 ( 
.A1(n_7249),
.A2(n_6298),
.B1(n_6547),
.B2(n_6580),
.Y(n_8330)
);

INVx2_ASAP7_75t_L g8331 ( 
.A(n_6701),
.Y(n_8331)
);

INVx1_ASAP7_75t_L g8332 ( 
.A(n_7188),
.Y(n_8332)
);

INVx2_ASAP7_75t_L g8333 ( 
.A(n_6714),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_7188),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7192),
.Y(n_8335)
);

HB1xp67_ASAP7_75t_L g8336 ( 
.A(n_7192),
.Y(n_8336)
);

INVx1_ASAP7_75t_L g8337 ( 
.A(n_7194),
.Y(n_8337)
);

INVx2_ASAP7_75t_L g8338 ( 
.A(n_6714),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_7194),
.Y(n_8339)
);

INVx2_ASAP7_75t_L g8340 ( 
.A(n_6714),
.Y(n_8340)
);

HB1xp67_ASAP7_75t_L g8341 ( 
.A(n_7204),
.Y(n_8341)
);

BUFx3_ASAP7_75t_L g8342 ( 
.A(n_6781),
.Y(n_8342)
);

OAI22xp33_ASAP7_75t_L g8343 ( 
.A1(n_7249),
.A2(n_6304),
.B1(n_6299),
.B2(n_6316),
.Y(n_8343)
);

OR2x2_ASAP7_75t_L g8344 ( 
.A(n_7635),
.B(n_6562),
.Y(n_8344)
);

INVx2_ASAP7_75t_L g8345 ( 
.A(n_6716),
.Y(n_8345)
);

AND2x4_ASAP7_75t_L g8346 ( 
.A(n_7704),
.B(n_6456),
.Y(n_8346)
);

AND2x2_ASAP7_75t_L g8347 ( 
.A(n_7151),
.B(n_6031),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_7204),
.Y(n_8348)
);

AOI22xp33_ASAP7_75t_SL g8349 ( 
.A1(n_7735),
.A2(n_6807),
.B1(n_6886),
.B2(n_6873),
.Y(n_8349)
);

INVx2_ASAP7_75t_L g8350 ( 
.A(n_6716),
.Y(n_8350)
);

INVx2_ASAP7_75t_L g8351 ( 
.A(n_6716),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_7208),
.Y(n_8352)
);

NAND2x1p5_ASAP7_75t_L g8353 ( 
.A(n_7043),
.B(n_5931),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_7208),
.Y(n_8354)
);

AND2x2_ASAP7_75t_L g8355 ( 
.A(n_6758),
.B(n_6469),
.Y(n_8355)
);

OA21x2_ASAP7_75t_L g8356 ( 
.A1(n_7349),
.A2(n_6251),
.B(n_6269),
.Y(n_8356)
);

OR2x2_ASAP7_75t_L g8357 ( 
.A(n_7660),
.B(n_6594),
.Y(n_8357)
);

INVx1_ASAP7_75t_L g8358 ( 
.A(n_7209),
.Y(n_8358)
);

AND2x2_ASAP7_75t_L g8359 ( 
.A(n_6758),
.B(n_6469),
.Y(n_8359)
);

INVx2_ASAP7_75t_L g8360 ( 
.A(n_6720),
.Y(n_8360)
);

INVx1_ASAP7_75t_SL g8361 ( 
.A(n_6894),
.Y(n_8361)
);

INVx2_ASAP7_75t_L g8362 ( 
.A(n_6720),
.Y(n_8362)
);

AND2x2_ASAP7_75t_L g8363 ( 
.A(n_6758),
.B(n_6469),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7209),
.Y(n_8364)
);

INVx1_ASAP7_75t_L g8365 ( 
.A(n_7227),
.Y(n_8365)
);

HB1xp67_ASAP7_75t_L g8366 ( 
.A(n_7227),
.Y(n_8366)
);

INVx2_ASAP7_75t_L g8367 ( 
.A(n_6720),
.Y(n_8367)
);

OA21x2_ASAP7_75t_L g8368 ( 
.A1(n_7349),
.A2(n_6269),
.B(n_6123),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_7233),
.Y(n_8369)
);

OAI21x1_ASAP7_75t_L g8370 ( 
.A1(n_7532),
.A2(n_6572),
.B(n_6126),
.Y(n_8370)
);

AOI22xp33_ASAP7_75t_SL g8371 ( 
.A1(n_7735),
.A2(n_6394),
.B1(n_6654),
.B2(n_6502),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_7233),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7248),
.Y(n_8373)
);

BUFx3_ASAP7_75t_L g8374 ( 
.A(n_6781),
.Y(n_8374)
);

INVx3_ASAP7_75t_L g8375 ( 
.A(n_6786),
.Y(n_8375)
);

AOI22xp33_ASAP7_75t_SL g8376 ( 
.A1(n_6873),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8376)
);

INVx3_ASAP7_75t_SL g8377 ( 
.A(n_7017),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_7248),
.Y(n_8378)
);

INVx1_ASAP7_75t_L g8379 ( 
.A(n_7252),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7252),
.Y(n_8380)
);

HB1xp67_ASAP7_75t_L g8381 ( 
.A(n_7257),
.Y(n_8381)
);

CKINVDCx14_ASAP7_75t_R g8382 ( 
.A(n_7262),
.Y(n_8382)
);

AND2x2_ASAP7_75t_L g8383 ( 
.A(n_6809),
.B(n_6496),
.Y(n_8383)
);

INVx3_ASAP7_75t_L g8384 ( 
.A(n_6966),
.Y(n_8384)
);

INVx1_ASAP7_75t_L g8385 ( 
.A(n_7257),
.Y(n_8385)
);

INVx1_ASAP7_75t_L g8386 ( 
.A(n_7265),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7265),
.Y(n_8387)
);

BUFx3_ASAP7_75t_L g8388 ( 
.A(n_6856),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7285),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7285),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_7294),
.Y(n_8391)
);

INVx3_ASAP7_75t_L g8392 ( 
.A(n_6966),
.Y(n_8392)
);

OA21x2_ASAP7_75t_L g8393 ( 
.A1(n_7246),
.A2(n_6123),
.B(n_6372),
.Y(n_8393)
);

OAI22xp5_ASAP7_75t_L g8394 ( 
.A1(n_6753),
.A2(n_6027),
.B1(n_6020),
.B2(n_6133),
.Y(n_8394)
);

HB1xp67_ASAP7_75t_L g8395 ( 
.A(n_7294),
.Y(n_8395)
);

INVx2_ASAP7_75t_L g8396 ( 
.A(n_6730),
.Y(n_8396)
);

INVx2_ASAP7_75t_L g8397 ( 
.A(n_6730),
.Y(n_8397)
);

HB1xp67_ASAP7_75t_L g8398 ( 
.A(n_7305),
.Y(n_8398)
);

AND2x2_ASAP7_75t_L g8399 ( 
.A(n_6809),
.B(n_6496),
.Y(n_8399)
);

AND2x2_ASAP7_75t_L g8400 ( 
.A(n_6809),
.B(n_6496),
.Y(n_8400)
);

OAI21xp5_ASAP7_75t_L g8401 ( 
.A1(n_7195),
.A2(n_6093),
.B(n_6070),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_6730),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_7305),
.Y(n_8403)
);

NAND2xp5_ASAP7_75t_L g8404 ( 
.A(n_7747),
.B(n_6594),
.Y(n_8404)
);

AOI22xp33_ASAP7_75t_L g8405 ( 
.A1(n_6752),
.A2(n_6131),
.B1(n_6539),
.B2(n_5932),
.Y(n_8405)
);

CKINVDCx20_ASAP7_75t_R g8406 ( 
.A(n_7009),
.Y(n_8406)
);

AND2x4_ASAP7_75t_L g8407 ( 
.A(n_6985),
.B(n_6456),
.Y(n_8407)
);

OAI21xp33_ASAP7_75t_SL g8408 ( 
.A1(n_7206),
.A2(n_7034),
.B(n_7005),
.Y(n_8408)
);

INVx8_ASAP7_75t_L g8409 ( 
.A(n_6818),
.Y(n_8409)
);

BUFx6f_ASAP7_75t_L g8410 ( 
.A(n_6700),
.Y(n_8410)
);

AND2x2_ASAP7_75t_L g8411 ( 
.A(n_6825),
.B(n_6515),
.Y(n_8411)
);

HB1xp67_ASAP7_75t_L g8412 ( 
.A(n_7309),
.Y(n_8412)
);

AO21x2_ASAP7_75t_L g8413 ( 
.A1(n_7391),
.A2(n_5996),
.B(n_6103),
.Y(n_8413)
);

INVx3_ASAP7_75t_L g8414 ( 
.A(n_6966),
.Y(n_8414)
);

BUFx12f_ASAP7_75t_L g8415 ( 
.A(n_7107),
.Y(n_8415)
);

INVx1_ASAP7_75t_L g8416 ( 
.A(n_7309),
.Y(n_8416)
);

INVx2_ASAP7_75t_L g8417 ( 
.A(n_6755),
.Y(n_8417)
);

BUFx6f_ASAP7_75t_L g8418 ( 
.A(n_6732),
.Y(n_8418)
);

NAND2x1p5_ASAP7_75t_L g8419 ( 
.A(n_7043),
.B(n_5931),
.Y(n_8419)
);

NAND2x1p5_ASAP7_75t_L g8420 ( 
.A(n_7043),
.B(n_5931),
.Y(n_8420)
);

BUFx10_ASAP7_75t_L g8421 ( 
.A(n_6676),
.Y(n_8421)
);

INVx3_ASAP7_75t_L g8422 ( 
.A(n_6966),
.Y(n_8422)
);

BUFx3_ASAP7_75t_L g8423 ( 
.A(n_6856),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_7312),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_6755),
.Y(n_8425)
);

AND2x2_ASAP7_75t_L g8426 ( 
.A(n_6825),
.B(n_6515),
.Y(n_8426)
);

BUFx4f_ASAP7_75t_SL g8427 ( 
.A(n_6709),
.Y(n_8427)
);

AND2x2_ASAP7_75t_L g8428 ( 
.A(n_6825),
.B(n_6515),
.Y(n_8428)
);

INVx2_ASAP7_75t_L g8429 ( 
.A(n_6755),
.Y(n_8429)
);

OAI22xp5_ASAP7_75t_L g8430 ( 
.A1(n_7001),
.A2(n_6027),
.B1(n_6210),
.B2(n_6131),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_7312),
.Y(n_8431)
);

NAND2xp5_ASAP7_75t_L g8432 ( 
.A(n_7747),
.B(n_7751),
.Y(n_8432)
);

INVx2_ASAP7_75t_SL g8433 ( 
.A(n_7043),
.Y(n_8433)
);

AOI22xp33_ASAP7_75t_SL g8434 ( 
.A1(n_6886),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8434)
);

INVx2_ASAP7_75t_L g8435 ( 
.A(n_6811),
.Y(n_8435)
);

OAI22xp33_ASAP7_75t_L g8436 ( 
.A1(n_7301),
.A2(n_6327),
.B1(n_6316),
.B2(n_6253),
.Y(n_8436)
);

AND2x2_ASAP7_75t_L g8437 ( 
.A(n_6887),
.B(n_6536),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7322),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_7322),
.Y(n_8439)
);

INVx2_ASAP7_75t_L g8440 ( 
.A(n_6811),
.Y(n_8440)
);

HB1xp67_ASAP7_75t_L g8441 ( 
.A(n_7333),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_7333),
.Y(n_8442)
);

INVx1_ASAP7_75t_L g8443 ( 
.A(n_7334),
.Y(n_8443)
);

INVx1_ASAP7_75t_L g8444 ( 
.A(n_7334),
.Y(n_8444)
);

BUFx3_ASAP7_75t_L g8445 ( 
.A(n_6856),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_7335),
.Y(n_8446)
);

INVx4_ASAP7_75t_L g8447 ( 
.A(n_6738),
.Y(n_8447)
);

AO21x1_ASAP7_75t_SL g8448 ( 
.A1(n_6883),
.A2(n_5969),
.B(n_6338),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_7335),
.Y(n_8449)
);

INVx2_ASAP7_75t_SL g8450 ( 
.A(n_7070),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_7339),
.Y(n_8451)
);

INVx2_ASAP7_75t_L g8452 ( 
.A(n_6811),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_7339),
.Y(n_8453)
);

OR2x6_ASAP7_75t_L g8454 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8454)
);

AOI22xp33_ASAP7_75t_L g8455 ( 
.A1(n_6752),
.A2(n_6539),
.B1(n_5932),
.B2(n_5897),
.Y(n_8455)
);

BUFx5_ASAP7_75t_L g8456 ( 
.A(n_7140),
.Y(n_8456)
);

AOI322xp5_ASAP7_75t_L g8457 ( 
.A1(n_7649),
.A2(n_5224),
.A3(n_5231),
.B1(n_5229),
.B2(n_6342),
.C1(n_6338),
.C2(n_6419),
.Y(n_8457)
);

BUFx8_ASAP7_75t_SL g8458 ( 
.A(n_6709),
.Y(n_8458)
);

INVx1_ASAP7_75t_L g8459 ( 
.A(n_7347),
.Y(n_8459)
);

INVx1_ASAP7_75t_L g8460 ( 
.A(n_7347),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_7348),
.Y(n_8461)
);

AOI222xp33_ASAP7_75t_L g8462 ( 
.A1(n_6708),
.A2(n_6374),
.B1(n_6306),
.B2(n_6332),
.C1(n_6354),
.C2(n_6342),
.Y(n_8462)
);

INVx1_ASAP7_75t_L g8463 ( 
.A(n_7348),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_7351),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_L g8465 ( 
.A(n_7751),
.B(n_6327),
.Y(n_8465)
);

AOI22xp33_ASAP7_75t_L g8466 ( 
.A1(n_6756),
.A2(n_5897),
.B1(n_6354),
.B2(n_6117),
.Y(n_8466)
);

INVx2_ASAP7_75t_L g8467 ( 
.A(n_6831),
.Y(n_8467)
);

OAI22xp33_ASAP7_75t_L g8468 ( 
.A1(n_7301),
.A2(n_6253),
.B1(n_6450),
.B2(n_6377),
.Y(n_8468)
);

BUFx3_ASAP7_75t_L g8469 ( 
.A(n_6856),
.Y(n_8469)
);

INVx2_ASAP7_75t_L g8470 ( 
.A(n_6831),
.Y(n_8470)
);

AOI22xp33_ASAP7_75t_L g8471 ( 
.A1(n_6756),
.A2(n_7649),
.B1(n_6731),
.B2(n_6703),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_6831),
.Y(n_8472)
);

HB1xp67_ASAP7_75t_L g8473 ( 
.A(n_7351),
.Y(n_8473)
);

INVx1_ASAP7_75t_L g8474 ( 
.A(n_7368),
.Y(n_8474)
);

INVx2_ASAP7_75t_L g8475 ( 
.A(n_6874),
.Y(n_8475)
);

HB1xp67_ASAP7_75t_L g8476 ( 
.A(n_7368),
.Y(n_8476)
);

OAI21x1_ASAP7_75t_L g8477 ( 
.A1(n_7532),
.A2(n_6126),
.B(n_5996),
.Y(n_8477)
);

INVx1_ASAP7_75t_L g8478 ( 
.A(n_7379),
.Y(n_8478)
);

HB1xp67_ASAP7_75t_L g8479 ( 
.A(n_7379),
.Y(n_8479)
);

AOI21xp33_ASAP7_75t_L g8480 ( 
.A1(n_6731),
.A2(n_6296),
.B(n_6287),
.Y(n_8480)
);

INVx2_ASAP7_75t_L g8481 ( 
.A(n_6874),
.Y(n_8481)
);

BUFx8_ASAP7_75t_L g8482 ( 
.A(n_6918),
.Y(n_8482)
);

HB1xp67_ASAP7_75t_L g8483 ( 
.A(n_7390),
.Y(n_8483)
);

INVx2_ASAP7_75t_L g8484 ( 
.A(n_6874),
.Y(n_8484)
);

OAI21x1_ASAP7_75t_L g8485 ( 
.A1(n_7532),
.A2(n_6124),
.B(n_6107),
.Y(n_8485)
);

OA21x2_ASAP7_75t_L g8486 ( 
.A1(n_7246),
.A2(n_6461),
.B(n_6372),
.Y(n_8486)
);

AOI22xp33_ASAP7_75t_SL g8487 ( 
.A1(n_6703),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8487)
);

OAI22xp5_ASAP7_75t_L g8488 ( 
.A1(n_7001),
.A2(n_6210),
.B1(n_5969),
.B2(n_6117),
.Y(n_8488)
);

INVx1_ASAP7_75t_L g8489 ( 
.A(n_7390),
.Y(n_8489)
);

INVx2_ASAP7_75t_L g8490 ( 
.A(n_6881),
.Y(n_8490)
);

INVx2_ASAP7_75t_L g8491 ( 
.A(n_6881),
.Y(n_8491)
);

AOI21x1_ASAP7_75t_L g8492 ( 
.A1(n_7495),
.A2(n_6273),
.B(n_6459),
.Y(n_8492)
);

NAND2xp5_ASAP7_75t_L g8493 ( 
.A(n_7706),
.B(n_6475),
.Y(n_8493)
);

INVx1_ASAP7_75t_L g8494 ( 
.A(n_7394),
.Y(n_8494)
);

INVx2_ASAP7_75t_L g8495 ( 
.A(n_6881),
.Y(n_8495)
);

INVx8_ASAP7_75t_L g8496 ( 
.A(n_6818),
.Y(n_8496)
);

OAI22xp33_ASAP7_75t_L g8497 ( 
.A1(n_7105),
.A2(n_6377),
.B1(n_6569),
.B2(n_6450),
.Y(n_8497)
);

AOI21x1_ASAP7_75t_L g8498 ( 
.A1(n_7495),
.A2(n_6273),
.B(n_6459),
.Y(n_8498)
);

AO21x2_ASAP7_75t_L g8499 ( 
.A1(n_7391),
.A2(n_6107),
.B(n_6103),
.Y(n_8499)
);

OAI21x1_ASAP7_75t_L g8500 ( 
.A1(n_7532),
.A2(n_6124),
.B(n_6005),
.Y(n_8500)
);

INVx2_ASAP7_75t_L g8501 ( 
.A(n_6912),
.Y(n_8501)
);

AND2x2_ASAP7_75t_L g8502 ( 
.A(n_6887),
.B(n_6536),
.Y(n_8502)
);

OAI21x1_ASAP7_75t_L g8503 ( 
.A1(n_7533),
.A2(n_6005),
.B(n_5936),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_7394),
.Y(n_8504)
);

INVx1_ASAP7_75t_L g8505 ( 
.A(n_7397),
.Y(n_8505)
);

OAI21x1_ASAP7_75t_L g8506 ( 
.A1(n_7533),
.A2(n_5936),
.B(n_6091),
.Y(n_8506)
);

AO21x1_ASAP7_75t_L g8507 ( 
.A1(n_6698),
.A2(n_6542),
.B(n_6541),
.Y(n_8507)
);

HB1xp67_ASAP7_75t_L g8508 ( 
.A(n_7397),
.Y(n_8508)
);

BUFx2_ASAP7_75t_L g8509 ( 
.A(n_7712),
.Y(n_8509)
);

AND2x2_ASAP7_75t_L g8510 ( 
.A(n_6887),
.B(n_6536),
.Y(n_8510)
);

AOI22xp5_ASAP7_75t_L g8511 ( 
.A1(n_6708),
.A2(n_5793),
.B1(n_6648),
.B2(n_6014),
.Y(n_8511)
);

AO21x2_ASAP7_75t_L g8512 ( 
.A1(n_7717),
.A2(n_6461),
.B(n_6463),
.Y(n_8512)
);

HB1xp67_ASAP7_75t_L g8513 ( 
.A(n_7404),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_7404),
.Y(n_8514)
);

INVx1_ASAP7_75t_L g8515 ( 
.A(n_7415),
.Y(n_8515)
);

INVx2_ASAP7_75t_SL g8516 ( 
.A(n_7070),
.Y(n_8516)
);

OAI21x1_ASAP7_75t_L g8517 ( 
.A1(n_7533),
.A2(n_6091),
.B(n_6110),
.Y(n_8517)
);

INVx1_ASAP7_75t_L g8518 ( 
.A(n_7415),
.Y(n_8518)
);

AOI22xp5_ASAP7_75t_SL g8519 ( 
.A1(n_7280),
.A2(n_6098),
.B1(n_6442),
.B2(n_6425),
.Y(n_8519)
);

OAI21x1_ASAP7_75t_L g8520 ( 
.A1(n_7533),
.A2(n_6110),
.B(n_6039),
.Y(n_8520)
);

INVx2_ASAP7_75t_L g8521 ( 
.A(n_6912),
.Y(n_8521)
);

AND2x2_ASAP7_75t_L g8522 ( 
.A(n_7422),
.B(n_6534),
.Y(n_8522)
);

OAI21x1_ASAP7_75t_L g8523 ( 
.A1(n_6744),
.A2(n_6039),
.B(n_6028),
.Y(n_8523)
);

INVx2_ASAP7_75t_L g8524 ( 
.A(n_6912),
.Y(n_8524)
);

AND2x2_ASAP7_75t_L g8525 ( 
.A(n_7422),
.B(n_6534),
.Y(n_8525)
);

BUFx3_ASAP7_75t_L g8526 ( 
.A(n_6861),
.Y(n_8526)
);

INVx1_ASAP7_75t_SL g8527 ( 
.A(n_6897),
.Y(n_8527)
);

AND2x2_ASAP7_75t_L g8528 ( 
.A(n_7422),
.B(n_6534),
.Y(n_8528)
);

INVx2_ASAP7_75t_L g8529 ( 
.A(n_6922),
.Y(n_8529)
);

INVx3_ASAP7_75t_L g8530 ( 
.A(n_6966),
.Y(n_8530)
);

BUFx3_ASAP7_75t_L g8531 ( 
.A(n_6861),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_6922),
.Y(n_8532)
);

INVx1_ASAP7_75t_L g8533 ( 
.A(n_7416),
.Y(n_8533)
);

OAI21xp5_ASAP7_75t_L g8534 ( 
.A1(n_7121),
.A2(n_6070),
.B(n_5837),
.Y(n_8534)
);

INVx1_ASAP7_75t_L g8535 ( 
.A(n_7416),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_7421),
.Y(n_8536)
);

INVx2_ASAP7_75t_SL g8537 ( 
.A(n_7070),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_7421),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_7435),
.Y(n_8539)
);

OR2x6_ASAP7_75t_L g8540 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8540)
);

AND2x2_ASAP7_75t_L g8541 ( 
.A(n_7428),
.B(n_6554),
.Y(n_8541)
);

HB1xp67_ASAP7_75t_L g8542 ( 
.A(n_7435),
.Y(n_8542)
);

INVx2_ASAP7_75t_L g8543 ( 
.A(n_6922),
.Y(n_8543)
);

BUFx2_ASAP7_75t_L g8544 ( 
.A(n_7712),
.Y(n_8544)
);

INVx2_ASAP7_75t_L g8545 ( 
.A(n_6924),
.Y(n_8545)
);

INVx3_ASAP7_75t_L g8546 ( 
.A(n_6966),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_7706),
.B(n_6475),
.Y(n_8547)
);

INVx1_ASAP7_75t_L g8548 ( 
.A(n_7440),
.Y(n_8548)
);

AOI22xp33_ASAP7_75t_SL g8549 ( 
.A1(n_6698),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8549)
);

HB1xp67_ASAP7_75t_L g8550 ( 
.A(n_7440),
.Y(n_8550)
);

AND2x4_ASAP7_75t_L g8551 ( 
.A(n_6985),
.B(n_6465),
.Y(n_8551)
);

INVx4_ASAP7_75t_L g8552 ( 
.A(n_6738),
.Y(n_8552)
);

INVx1_ASAP7_75t_L g8553 ( 
.A(n_7445),
.Y(n_8553)
);

INVx2_ASAP7_75t_L g8554 ( 
.A(n_6924),
.Y(n_8554)
);

INVx1_ASAP7_75t_L g8555 ( 
.A(n_7445),
.Y(n_8555)
);

INVx1_ASAP7_75t_L g8556 ( 
.A(n_7452),
.Y(n_8556)
);

NAND2xp5_ASAP7_75t_L g8557 ( 
.A(n_7709),
.B(n_6204),
.Y(n_8557)
);

BUFx2_ASAP7_75t_L g8558 ( 
.A(n_7539),
.Y(n_8558)
);

BUFx6f_ASAP7_75t_SL g8559 ( 
.A(n_6739),
.Y(n_8559)
);

OAI22xp5_ASAP7_75t_L g8560 ( 
.A1(n_7064),
.A2(n_6369),
.B1(n_6096),
.B2(n_6198),
.Y(n_8560)
);

INVx2_ASAP7_75t_L g8561 ( 
.A(n_6924),
.Y(n_8561)
);

OR2x2_ASAP7_75t_L g8562 ( 
.A(n_7660),
.B(n_6541),
.Y(n_8562)
);

INVx2_ASAP7_75t_L g8563 ( 
.A(n_6931),
.Y(n_8563)
);

OA21x2_ASAP7_75t_L g8564 ( 
.A1(n_7271),
.A2(n_6481),
.B(n_6463),
.Y(n_8564)
);

INVx2_ASAP7_75t_L g8565 ( 
.A(n_6931),
.Y(n_8565)
);

BUFx2_ASAP7_75t_L g8566 ( 
.A(n_7539),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7452),
.Y(n_8567)
);

INVx1_ASAP7_75t_L g8568 ( 
.A(n_7468),
.Y(n_8568)
);

CKINVDCx11_ASAP7_75t_R g8569 ( 
.A(n_6709),
.Y(n_8569)
);

HB1xp67_ASAP7_75t_SL g8570 ( 
.A(n_6861),
.Y(n_8570)
);

INVx1_ASAP7_75t_L g8571 ( 
.A(n_7468),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_7469),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_7469),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_7471),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_7471),
.Y(n_8575)
);

CKINVDCx20_ASAP7_75t_R g8576 ( 
.A(n_7028),
.Y(n_8576)
);

BUFx3_ASAP7_75t_L g8577 ( 
.A(n_6861),
.Y(n_8577)
);

INVx1_ASAP7_75t_L g8578 ( 
.A(n_7473),
.Y(n_8578)
);

HB1xp67_ASAP7_75t_L g8579 ( 
.A(n_7473),
.Y(n_8579)
);

AOI21x1_ASAP7_75t_L g8580 ( 
.A1(n_7632),
.A2(n_6380),
.B(n_6365),
.Y(n_8580)
);

INVx2_ASAP7_75t_L g8581 ( 
.A(n_6931),
.Y(n_8581)
);

INVx1_ASAP7_75t_L g8582 ( 
.A(n_7487),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_7487),
.Y(n_8583)
);

NAND2xp5_ASAP7_75t_L g8584 ( 
.A(n_7709),
.B(n_6204),
.Y(n_8584)
);

OAI21x1_ASAP7_75t_L g8585 ( 
.A1(n_6744),
.A2(n_6051),
.B(n_6028),
.Y(n_8585)
);

HB1xp67_ASAP7_75t_L g8586 ( 
.A(n_7493),
.Y(n_8586)
);

HB1xp67_ASAP7_75t_L g8587 ( 
.A(n_7493),
.Y(n_8587)
);

INVx1_ASAP7_75t_L g8588 ( 
.A(n_7501),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_6936),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_7501),
.Y(n_8590)
);

INVxp67_ASAP7_75t_SL g8591 ( 
.A(n_6688),
.Y(n_8591)
);

CKINVDCx20_ASAP7_75t_R g8592 ( 
.A(n_7037),
.Y(n_8592)
);

CKINVDCx11_ASAP7_75t_R g8593 ( 
.A(n_6762),
.Y(n_8593)
);

INVx1_ASAP7_75t_L g8594 ( 
.A(n_7505),
.Y(n_8594)
);

HB1xp67_ASAP7_75t_L g8595 ( 
.A(n_7505),
.Y(n_8595)
);

INVx2_ASAP7_75t_SL g8596 ( 
.A(n_7070),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_7514),
.Y(n_8597)
);

INVx2_ASAP7_75t_L g8598 ( 
.A(n_6936),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_7514),
.Y(n_8599)
);

OA21x2_ASAP7_75t_L g8600 ( 
.A1(n_7271),
.A2(n_6484),
.B(n_6481),
.Y(n_8600)
);

INVx2_ASAP7_75t_L g8601 ( 
.A(n_6936),
.Y(n_8601)
);

INVx3_ASAP7_75t_L g8602 ( 
.A(n_6966),
.Y(n_8602)
);

AOI21x1_ASAP7_75t_L g8603 ( 
.A1(n_7632),
.A2(n_6380),
.B(n_6365),
.Y(n_8603)
);

NAND2x1p5_ASAP7_75t_L g8604 ( 
.A(n_7070),
.B(n_5931),
.Y(n_8604)
);

INVx1_ASAP7_75t_L g8605 ( 
.A(n_7521),
.Y(n_8605)
);

INVx1_ASAP7_75t_SL g8606 ( 
.A(n_6897),
.Y(n_8606)
);

CKINVDCx5p33_ASAP7_75t_R g8607 ( 
.A(n_7038),
.Y(n_8607)
);

INVx2_ASAP7_75t_L g8608 ( 
.A(n_6963),
.Y(n_8608)
);

NAND2xp5_ASAP7_75t_L g8609 ( 
.A(n_7146),
.B(n_6228),
.Y(n_8609)
);

OAI22xp5_ASAP7_75t_L g8610 ( 
.A1(n_7064),
.A2(n_6369),
.B1(n_6096),
.B2(n_6198),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_7521),
.Y(n_8611)
);

HB1xp67_ASAP7_75t_L g8612 ( 
.A(n_7524),
.Y(n_8612)
);

INVx1_ASAP7_75t_L g8613 ( 
.A(n_7524),
.Y(n_8613)
);

NOR2xp33_ASAP7_75t_L g8614 ( 
.A(n_6743),
.B(n_6525),
.Y(n_8614)
);

AND2x2_ASAP7_75t_L g8615 ( 
.A(n_7428),
.B(n_6554),
.Y(n_8615)
);

OAI22xp5_ASAP7_75t_L g8616 ( 
.A1(n_7089),
.A2(n_6014),
.B1(n_6076),
.B2(n_6399),
.Y(n_8616)
);

CKINVDCx11_ASAP7_75t_R g8617 ( 
.A(n_6762),
.Y(n_8617)
);

INVx2_ASAP7_75t_L g8618 ( 
.A(n_6963),
.Y(n_8618)
);

AND2x2_ASAP7_75t_L g8619 ( 
.A(n_7428),
.B(n_6554),
.Y(n_8619)
);

INVx1_ASAP7_75t_L g8620 ( 
.A(n_7538),
.Y(n_8620)
);

BUFx2_ASAP7_75t_SL g8621 ( 
.A(n_6682),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_7538),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_6963),
.Y(n_8623)
);

BUFx4f_ASAP7_75t_SL g8624 ( 
.A(n_6762),
.Y(n_8624)
);

INVx2_ASAP7_75t_L g8625 ( 
.A(n_6981),
.Y(n_8625)
);

BUFx6f_ASAP7_75t_L g8626 ( 
.A(n_6732),
.Y(n_8626)
);

BUFx2_ASAP7_75t_L g8627 ( 
.A(n_7609),
.Y(n_8627)
);

AND2x2_ASAP7_75t_L g8628 ( 
.A(n_7451),
.B(n_6561),
.Y(n_8628)
);

AND2x2_ASAP7_75t_L g8629 ( 
.A(n_7451),
.B(n_6561),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_7542),
.Y(n_8630)
);

NAND2xp5_ASAP7_75t_L g8631 ( 
.A(n_7146),
.B(n_6228),
.Y(n_8631)
);

INVx1_ASAP7_75t_L g8632 ( 
.A(n_7542),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_7554),
.Y(n_8633)
);

AOI22xp33_ASAP7_75t_L g8634 ( 
.A1(n_6759),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8634)
);

INVx1_ASAP7_75t_L g8635 ( 
.A(n_7554),
.Y(n_8635)
);

INVx1_ASAP7_75t_L g8636 ( 
.A(n_7556),
.Y(n_8636)
);

INVx2_ASAP7_75t_L g8637 ( 
.A(n_6981),
.Y(n_8637)
);

BUFx3_ASAP7_75t_L g8638 ( 
.A(n_6934),
.Y(n_8638)
);

INVx1_ASAP7_75t_L g8639 ( 
.A(n_7556),
.Y(n_8639)
);

CKINVDCx11_ASAP7_75t_R g8640 ( 
.A(n_6768),
.Y(n_8640)
);

INVx1_ASAP7_75t_L g8641 ( 
.A(n_7557),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_7557),
.Y(n_8642)
);

INVx2_ASAP7_75t_L g8643 ( 
.A(n_6981),
.Y(n_8643)
);

INVx1_ASAP7_75t_L g8644 ( 
.A(n_7561),
.Y(n_8644)
);

INVx2_ASAP7_75t_L g8645 ( 
.A(n_7003),
.Y(n_8645)
);

CKINVDCx20_ASAP7_75t_R g8646 ( 
.A(n_6860),
.Y(n_8646)
);

INVx2_ASAP7_75t_L g8647 ( 
.A(n_7003),
.Y(n_8647)
);

INVxp33_ASAP7_75t_L g8648 ( 
.A(n_7273),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_7561),
.Y(n_8649)
);

AND2x2_ASAP7_75t_L g8650 ( 
.A(n_7451),
.B(n_6561),
.Y(n_8650)
);

AND2x2_ASAP7_75t_L g8651 ( 
.A(n_7613),
.B(n_6570),
.Y(n_8651)
);

AOI22xp33_ASAP7_75t_L g8652 ( 
.A1(n_6759),
.A2(n_6450),
.B1(n_6569),
.B2(n_6377),
.Y(n_8652)
);

INVx3_ASAP7_75t_L g8653 ( 
.A(n_6983),
.Y(n_8653)
);

INVx1_ASAP7_75t_L g8654 ( 
.A(n_7569),
.Y(n_8654)
);

INVx2_ASAP7_75t_L g8655 ( 
.A(n_7003),
.Y(n_8655)
);

OAI21x1_ASAP7_75t_L g8656 ( 
.A1(n_6744),
.A2(n_6053),
.B(n_6051),
.Y(n_8656)
);

INVx2_ASAP7_75t_L g8657 ( 
.A(n_7008),
.Y(n_8657)
);

CKINVDCx20_ASAP7_75t_R g8658 ( 
.A(n_6911),
.Y(n_8658)
);

CKINVDCx20_ASAP7_75t_R g8659 ( 
.A(n_6919),
.Y(n_8659)
);

AND2x4_ASAP7_75t_L g8660 ( 
.A(n_6985),
.B(n_6465),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_7008),
.Y(n_8661)
);

INVx2_ASAP7_75t_L g8662 ( 
.A(n_7008),
.Y(n_8662)
);

BUFx2_ASAP7_75t_L g8663 ( 
.A(n_7609),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_7569),
.Y(n_8664)
);

INVx1_ASAP7_75t_L g8665 ( 
.A(n_7571),
.Y(n_8665)
);

INVx2_ASAP7_75t_L g8666 ( 
.A(n_7012),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_7571),
.Y(n_8667)
);

INVx2_ASAP7_75t_L g8668 ( 
.A(n_7012),
.Y(n_8668)
);

AND2x2_ASAP7_75t_L g8669 ( 
.A(n_7613),
.B(n_6570),
.Y(n_8669)
);

INVx1_ASAP7_75t_L g8670 ( 
.A(n_7582),
.Y(n_8670)
);

AO21x1_ASAP7_75t_L g8671 ( 
.A1(n_6784),
.A2(n_6542),
.B(n_6541),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_7012),
.Y(n_8672)
);

BUFx3_ASAP7_75t_L g8673 ( 
.A(n_6934),
.Y(n_8673)
);

HB1xp67_ASAP7_75t_L g8674 ( 
.A(n_7582),
.Y(n_8674)
);

AOI22xp33_ASAP7_75t_SL g8675 ( 
.A1(n_6764),
.A2(n_6569),
.B1(n_6656),
.B2(n_6433),
.Y(n_8675)
);

OAI21x1_ASAP7_75t_L g8676 ( 
.A1(n_6744),
.A2(n_6055),
.B(n_6053),
.Y(n_8676)
);

OA21x2_ASAP7_75t_L g8677 ( 
.A1(n_7499),
.A2(n_6501),
.B(n_6484),
.Y(n_8677)
);

AND2x4_ASAP7_75t_L g8678 ( 
.A(n_6985),
.B(n_6465),
.Y(n_8678)
);

BUFx2_ASAP7_75t_R g8679 ( 
.A(n_6777),
.Y(n_8679)
);

AOI22xp33_ASAP7_75t_SL g8680 ( 
.A1(n_6764),
.A2(n_6656),
.B1(n_6433),
.B2(n_6438),
.Y(n_8680)
);

BUFx2_ASAP7_75t_L g8681 ( 
.A(n_7658),
.Y(n_8681)
);

INVx1_ASAP7_75t_L g8682 ( 
.A(n_7584),
.Y(n_8682)
);

INVx1_ASAP7_75t_L g8683 ( 
.A(n_7584),
.Y(n_8683)
);

INVx1_ASAP7_75t_L g8684 ( 
.A(n_7585),
.Y(n_8684)
);

BUFx6f_ASAP7_75t_L g8685 ( 
.A(n_6732),
.Y(n_8685)
);

INVx2_ASAP7_75t_L g8686 ( 
.A(n_7031),
.Y(n_8686)
);

INVx2_ASAP7_75t_L g8687 ( 
.A(n_7031),
.Y(n_8687)
);

OR2x2_ASAP7_75t_L g8688 ( 
.A(n_7705),
.B(n_6542),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_7585),
.Y(n_8689)
);

NAND2x1p5_ASAP7_75t_L g8690 ( 
.A(n_7070),
.B(n_5931),
.Y(n_8690)
);

INVx2_ASAP7_75t_L g8691 ( 
.A(n_7031),
.Y(n_8691)
);

INVx1_ASAP7_75t_L g8692 ( 
.A(n_7605),
.Y(n_8692)
);

HB1xp67_ASAP7_75t_L g8693 ( 
.A(n_7605),
.Y(n_8693)
);

AOI21x1_ASAP7_75t_L g8694 ( 
.A1(n_7601),
.A2(n_6212),
.B(n_5955),
.Y(n_8694)
);

INVx1_ASAP7_75t_L g8695 ( 
.A(n_7610),
.Y(n_8695)
);

INVx3_ASAP7_75t_L g8696 ( 
.A(n_6983),
.Y(n_8696)
);

OAI321xp33_ASAP7_75t_L g8697 ( 
.A1(n_6784),
.A2(n_6058),
.A3(n_6567),
.B1(n_6652),
.B2(n_6076),
.C(n_6419),
.Y(n_8697)
);

INVx2_ASAP7_75t_SL g8698 ( 
.A(n_7070),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_L g8699 ( 
.A(n_6688),
.B(n_5965),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_7610),
.Y(n_8700)
);

AOI21x1_ASAP7_75t_L g8701 ( 
.A1(n_7601),
.A2(n_6400),
.B(n_6388),
.Y(n_8701)
);

BUFx2_ASAP7_75t_L g8702 ( 
.A(n_7658),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_7612),
.Y(n_8703)
);

INVx2_ASAP7_75t_L g8704 ( 
.A(n_7058),
.Y(n_8704)
);

NAND2xp5_ASAP7_75t_L g8705 ( 
.A(n_6757),
.B(n_5965),
.Y(n_8705)
);

NAND2x1p5_ASAP7_75t_L g8706 ( 
.A(n_7083),
.B(n_5931),
.Y(n_8706)
);

AO21x1_ASAP7_75t_SL g8707 ( 
.A1(n_6883),
.A2(n_6399),
.B(n_5231),
.Y(n_8707)
);

INVx3_ASAP7_75t_L g8708 ( 
.A(n_6983),
.Y(n_8708)
);

INVx1_ASAP7_75t_L g8709 ( 
.A(n_7612),
.Y(n_8709)
);

HB1xp67_ASAP7_75t_L g8710 ( 
.A(n_7616),
.Y(n_8710)
);

INVx2_ASAP7_75t_L g8711 ( 
.A(n_7058),
.Y(n_8711)
);

HB1xp67_ASAP7_75t_L g8712 ( 
.A(n_7616),
.Y(n_8712)
);

BUFx3_ASAP7_75t_L g8713 ( 
.A(n_6934),
.Y(n_8713)
);

CKINVDCx16_ASAP7_75t_R g8714 ( 
.A(n_6682),
.Y(n_8714)
);

INVx2_ASAP7_75t_L g8715 ( 
.A(n_7058),
.Y(n_8715)
);

INVx1_ASAP7_75t_L g8716 ( 
.A(n_7620),
.Y(n_8716)
);

INVx1_ASAP7_75t_L g8717 ( 
.A(n_7620),
.Y(n_8717)
);

BUFx3_ASAP7_75t_L g8718 ( 
.A(n_6934),
.Y(n_8718)
);

NAND2xp5_ASAP7_75t_L g8719 ( 
.A(n_6757),
.B(n_5973),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_7627),
.Y(n_8720)
);

OR2x6_ASAP7_75t_L g8721 ( 
.A(n_7684),
.B(n_6455),
.Y(n_8721)
);

OAI21x1_ASAP7_75t_L g8722 ( 
.A1(n_6896),
.A2(n_6065),
.B(n_6055),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_7084),
.Y(n_8723)
);

INVx2_ASAP7_75t_L g8724 ( 
.A(n_7084),
.Y(n_8724)
);

NAND2xp5_ASAP7_75t_L g8725 ( 
.A(n_6694),
.B(n_5973),
.Y(n_8725)
);

BUFx6f_ASAP7_75t_L g8726 ( 
.A(n_6732),
.Y(n_8726)
);

INVx3_ASAP7_75t_L g8727 ( 
.A(n_6983),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_7627),
.Y(n_8728)
);

AOI22xp33_ASAP7_75t_L g8729 ( 
.A1(n_6988),
.A2(n_6363),
.B1(n_6498),
.B2(n_6168),
.Y(n_8729)
);

BUFx6f_ASAP7_75t_L g8730 ( 
.A(n_6732),
.Y(n_8730)
);

BUFx10_ASAP7_75t_L g8731 ( 
.A(n_6676),
.Y(n_8731)
);

INVx2_ASAP7_75t_L g8732 ( 
.A(n_7084),
.Y(n_8732)
);

OAI21x1_ASAP7_75t_L g8733 ( 
.A1(n_6896),
.A2(n_6082),
.B(n_6065),
.Y(n_8733)
);

CKINVDCx5p33_ASAP7_75t_R g8734 ( 
.A(n_7038),
.Y(n_8734)
);

INVx3_ASAP7_75t_L g8735 ( 
.A(n_6983),
.Y(n_8735)
);

INVx2_ASAP7_75t_L g8736 ( 
.A(n_7094),
.Y(n_8736)
);

INVx5_ASAP7_75t_L g8737 ( 
.A(n_6732),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_7647),
.Y(n_8738)
);

INVx1_ASAP7_75t_L g8739 ( 
.A(n_7647),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_7659),
.Y(n_8740)
);

AND2x2_ASAP7_75t_L g8741 ( 
.A(n_7613),
.B(n_7695),
.Y(n_8741)
);

AOI21x1_ASAP7_75t_L g8742 ( 
.A1(n_7601),
.A2(n_6400),
.B(n_6388),
.Y(n_8742)
);

INVx3_ASAP7_75t_L g8743 ( 
.A(n_6983),
.Y(n_8743)
);

INVx1_ASAP7_75t_L g8744 ( 
.A(n_7659),
.Y(n_8744)
);

AOI21x1_ASAP7_75t_L g8745 ( 
.A1(n_7765),
.A2(n_7393),
.B(n_7304),
.Y(n_8745)
);

INVxp33_ASAP7_75t_SL g8746 ( 
.A(n_7433),
.Y(n_8746)
);

INVx2_ASAP7_75t_L g8747 ( 
.A(n_7094),
.Y(n_8747)
);

INVxp67_ASAP7_75t_SL g8748 ( 
.A(n_6926),
.Y(n_8748)
);

CKINVDCx6p67_ASAP7_75t_R g8749 ( 
.A(n_6918),
.Y(n_8749)
);

INVx1_ASAP7_75t_L g8750 ( 
.A(n_7670),
.Y(n_8750)
);

BUFx3_ASAP7_75t_L g8751 ( 
.A(n_6995),
.Y(n_8751)
);

BUFx2_ASAP7_75t_L g8752 ( 
.A(n_7083),
.Y(n_8752)
);

OAI21x1_ASAP7_75t_L g8753 ( 
.A1(n_6896),
.A2(n_6129),
.B(n_6082),
.Y(n_8753)
);

AND2x4_ASAP7_75t_L g8754 ( 
.A(n_7092),
.B(n_6465),
.Y(n_8754)
);

NOR2xp33_ASAP7_75t_L g8755 ( 
.A(n_6743),
.B(n_6003),
.Y(n_8755)
);

INVx2_ASAP7_75t_L g8756 ( 
.A(n_7094),
.Y(n_8756)
);

BUFx12f_ASAP7_75t_L g8757 ( 
.A(n_7117),
.Y(n_8757)
);

BUFx3_ASAP7_75t_L g8758 ( 
.A(n_6995),
.Y(n_8758)
);

INVx1_ASAP7_75t_L g8759 ( 
.A(n_7670),
.Y(n_8759)
);

AOI21x1_ASAP7_75t_L g8760 ( 
.A1(n_7765),
.A2(n_6212),
.B(n_5955),
.Y(n_8760)
);

INVx1_ASAP7_75t_L g8761 ( 
.A(n_7679),
.Y(n_8761)
);

INVx4_ASAP7_75t_L g8762 ( 
.A(n_6739),
.Y(n_8762)
);

INVx2_ASAP7_75t_L g8763 ( 
.A(n_7112),
.Y(n_8763)
);

INVxp67_ASAP7_75t_L g8764 ( 
.A(n_7503),
.Y(n_8764)
);

INVx2_ASAP7_75t_L g8765 ( 
.A(n_7112),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_7679),
.Y(n_8766)
);

OR2x2_ASAP7_75t_L g8767 ( 
.A(n_7705),
.B(n_6567),
.Y(n_8767)
);

INVx2_ASAP7_75t_L g8768 ( 
.A(n_7112),
.Y(n_8768)
);

INVx2_ASAP7_75t_L g8769 ( 
.A(n_7132),
.Y(n_8769)
);

INVx1_ASAP7_75t_L g8770 ( 
.A(n_7687),
.Y(n_8770)
);

AO21x1_ASAP7_75t_L g8771 ( 
.A1(n_7502),
.A2(n_6567),
.B(n_6058),
.Y(n_8771)
);

INVx2_ASAP7_75t_L g8772 ( 
.A(n_7132),
.Y(n_8772)
);

INVx1_ASAP7_75t_L g8773 ( 
.A(n_7687),
.Y(n_8773)
);

INVx1_ASAP7_75t_L g8774 ( 
.A(n_7694),
.Y(n_8774)
);

AO21x1_ASAP7_75t_SL g8775 ( 
.A1(n_7105),
.A2(n_5231),
.B(n_5229),
.Y(n_8775)
);

INVx2_ASAP7_75t_L g8776 ( 
.A(n_7132),
.Y(n_8776)
);

OAI21x1_ASAP7_75t_L g8777 ( 
.A1(n_6896),
.A2(n_6129),
.B(n_6125),
.Y(n_8777)
);

INVx1_ASAP7_75t_L g8778 ( 
.A(n_7694),
.Y(n_8778)
);

INVx3_ASAP7_75t_L g8779 ( 
.A(n_6983),
.Y(n_8779)
);

INVx2_ASAP7_75t_L g8780 ( 
.A(n_7137),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_7708),
.Y(n_8781)
);

AND2x2_ASAP7_75t_L g8782 ( 
.A(n_7695),
.B(n_6570),
.Y(n_8782)
);

INVx2_ASAP7_75t_L g8783 ( 
.A(n_7137),
.Y(n_8783)
);

INVx2_ASAP7_75t_L g8784 ( 
.A(n_7137),
.Y(n_8784)
);

INVx1_ASAP7_75t_L g8785 ( 
.A(n_7708),
.Y(n_8785)
);

BUFx8_ASAP7_75t_SL g8786 ( 
.A(n_6768),
.Y(n_8786)
);

INVx2_ASAP7_75t_L g8787 ( 
.A(n_7142),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_L g8788 ( 
.A(n_6694),
.B(n_5988),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_7715),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_7715),
.Y(n_8790)
);

AND2x2_ASAP7_75t_L g8791 ( 
.A(n_7695),
.B(n_6581),
.Y(n_8791)
);

BUFx2_ASAP7_75t_L g8792 ( 
.A(n_7083),
.Y(n_8792)
);

INVx1_ASAP7_75t_L g8793 ( 
.A(n_7722),
.Y(n_8793)
);

OR2x2_ASAP7_75t_L g8794 ( 
.A(n_7549),
.B(n_6577),
.Y(n_8794)
);

INVx2_ASAP7_75t_L g8795 ( 
.A(n_7142),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_7722),
.Y(n_8796)
);

AOI222xp33_ASAP7_75t_L g8797 ( 
.A1(n_6824),
.A2(n_6332),
.B1(n_6306),
.B2(n_6296),
.C1(n_5799),
.C2(n_5813),
.Y(n_8797)
);

INVx2_ASAP7_75t_L g8798 ( 
.A(n_7142),
.Y(n_8798)
);

INVx1_ASAP7_75t_L g8799 ( 
.A(n_7723),
.Y(n_8799)
);

AND2x2_ASAP7_75t_L g8800 ( 
.A(n_7597),
.B(n_6581),
.Y(n_8800)
);

HB1xp67_ASAP7_75t_L g8801 ( 
.A(n_7723),
.Y(n_8801)
);

HB1xp67_ASAP7_75t_L g8802 ( 
.A(n_7729),
.Y(n_8802)
);

INVx1_ASAP7_75t_L g8803 ( 
.A(n_7729),
.Y(n_8803)
);

INVx3_ASAP7_75t_L g8804 ( 
.A(n_7004),
.Y(n_8804)
);

INVx2_ASAP7_75t_L g8805 ( 
.A(n_7144),
.Y(n_8805)
);

BUFx10_ASAP7_75t_L g8806 ( 
.A(n_6676),
.Y(n_8806)
);

INVx3_ASAP7_75t_L g8807 ( 
.A(n_7004),
.Y(n_8807)
);

OAI222xp33_ASAP7_75t_L g8808 ( 
.A1(n_6940),
.A2(n_6652),
.B1(n_6385),
.B2(n_6386),
.C1(n_6379),
.C2(n_6387),
.Y(n_8808)
);

INVx1_ASAP7_75t_L g8809 ( 
.A(n_7731),
.Y(n_8809)
);

INVx2_ASAP7_75t_L g8810 ( 
.A(n_7144),
.Y(n_8810)
);

HB1xp67_ASAP7_75t_L g8811 ( 
.A(n_7731),
.Y(n_8811)
);

CKINVDCx11_ASAP7_75t_R g8812 ( 
.A(n_6768),
.Y(n_8812)
);

HB1xp67_ASAP7_75t_L g8813 ( 
.A(n_7737),
.Y(n_8813)
);

BUFx3_ASAP7_75t_L g8814 ( 
.A(n_8040),
.Y(n_8814)
);

AO21x2_ASAP7_75t_L g8815 ( 
.A1(n_8771),
.A2(n_7499),
.B(n_7717),
.Y(n_8815)
);

HB1xp67_ASAP7_75t_L g8816 ( 
.A(n_8242),
.Y(n_8816)
);

INVx1_ASAP7_75t_L g8817 ( 
.A(n_7793),
.Y(n_8817)
);

AO21x2_ASAP7_75t_L g8818 ( 
.A1(n_8771),
.A2(n_7268),
.B(n_7220),
.Y(n_8818)
);

AO31x2_ASAP7_75t_L g8819 ( 
.A1(n_8771),
.A2(n_7765),
.A3(n_6956),
.B(n_6978),
.Y(n_8819)
);

OR2x2_ASAP7_75t_L g8820 ( 
.A(n_8465),
.B(n_7000),
.Y(n_8820)
);

BUFx2_ASAP7_75t_L g8821 ( 
.A(n_7884),
.Y(n_8821)
);

INVx1_ASAP7_75t_L g8822 ( 
.A(n_7793),
.Y(n_8822)
);

INVx2_ASAP7_75t_L g8823 ( 
.A(n_7847),
.Y(n_8823)
);

HB1xp67_ASAP7_75t_L g8824 ( 
.A(n_8242),
.Y(n_8824)
);

AND2x2_ASAP7_75t_L g8825 ( 
.A(n_7893),
.B(n_7016),
.Y(n_8825)
);

INVx2_ASAP7_75t_L g8826 ( 
.A(n_7847),
.Y(n_8826)
);

INVx1_ASAP7_75t_L g8827 ( 
.A(n_7797),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_7847),
.Y(n_8828)
);

HB1xp67_ASAP7_75t_L g8829 ( 
.A(n_8361),
.Y(n_8829)
);

BUFx3_ASAP7_75t_L g8830 ( 
.A(n_8040),
.Y(n_8830)
);

INVxp67_ASAP7_75t_L g8831 ( 
.A(n_8106),
.Y(n_8831)
);

HB1xp67_ASAP7_75t_L g8832 ( 
.A(n_8361),
.Y(n_8832)
);

BUFx2_ASAP7_75t_SL g8833 ( 
.A(n_8135),
.Y(n_8833)
);

INVx2_ASAP7_75t_L g8834 ( 
.A(n_7962),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_7962),
.Y(n_8835)
);

INVx1_ASAP7_75t_L g8836 ( 
.A(n_7797),
.Y(n_8836)
);

INVx1_ASAP7_75t_L g8837 ( 
.A(n_7800),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_7800),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_7802),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_7962),
.Y(n_8840)
);

OR2x2_ASAP7_75t_L g8841 ( 
.A(n_8465),
.B(n_8272),
.Y(n_8841)
);

INVx1_ASAP7_75t_L g8842 ( 
.A(n_7802),
.Y(n_8842)
);

AO21x1_ASAP7_75t_SL g8843 ( 
.A1(n_7982),
.A2(n_7046),
.B(n_7045),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_7806),
.Y(n_8844)
);

INVx2_ASAP7_75t_L g8845 ( 
.A(n_8184),
.Y(n_8845)
);

AO21x2_ASAP7_75t_L g8846 ( 
.A1(n_8507),
.A2(n_7268),
.B(n_7220),
.Y(n_8846)
);

AND2x2_ASAP7_75t_L g8847 ( 
.A(n_7893),
.B(n_7016),
.Y(n_8847)
);

INVx2_ASAP7_75t_L g8848 ( 
.A(n_8184),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_8184),
.Y(n_8849)
);

INVx1_ASAP7_75t_L g8850 ( 
.A(n_7806),
.Y(n_8850)
);

OAI21xp5_ASAP7_75t_L g8851 ( 
.A1(n_7982),
.A2(n_7121),
.B(n_6987),
.Y(n_8851)
);

INVx3_ASAP7_75t_L g8852 ( 
.A(n_7863),
.Y(n_8852)
);

AND4x1_ASAP7_75t_L g8853 ( 
.A(n_8471),
.B(n_7226),
.C(n_7552),
.D(n_7550),
.Y(n_8853)
);

OR2x2_ASAP7_75t_L g8854 ( 
.A(n_8272),
.B(n_7000),
.Y(n_8854)
);

INVx1_ASAP7_75t_L g8855 ( 
.A(n_7818),
.Y(n_8855)
);

NAND2xp5_ASAP7_75t_L g8856 ( 
.A(n_7799),
.B(n_7340),
.Y(n_8856)
);

INVx1_ASAP7_75t_L g8857 ( 
.A(n_7818),
.Y(n_8857)
);

AO21x2_ASAP7_75t_L g8858 ( 
.A1(n_8507),
.A2(n_7760),
.B(n_7211),
.Y(n_8858)
);

CKINVDCx16_ASAP7_75t_R g8859 ( 
.A(n_8246),
.Y(n_8859)
);

AND2x2_ASAP7_75t_L g8860 ( 
.A(n_7893),
.B(n_7900),
.Y(n_8860)
);

NAND2x1p5_ASAP7_75t_L g8861 ( 
.A(n_8737),
.B(n_7083),
.Y(n_8861)
);

INVx1_ASAP7_75t_L g8862 ( 
.A(n_7822),
.Y(n_8862)
);

OA21x2_ASAP7_75t_L g8863 ( 
.A1(n_8290),
.A2(n_7211),
.B(n_7136),
.Y(n_8863)
);

OR2x2_ASAP7_75t_L g8864 ( 
.A(n_8699),
.B(n_7483),
.Y(n_8864)
);

OAI21x1_ASAP7_75t_L g8865 ( 
.A1(n_8745),
.A2(n_7063),
.B(n_6968),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_7822),
.Y(n_8866)
);

INVx1_ASAP7_75t_SL g8867 ( 
.A(n_8679),
.Y(n_8867)
);

INVx2_ASAP7_75t_L g8868 ( 
.A(n_8265),
.Y(n_8868)
);

INVx2_ASAP7_75t_L g8869 ( 
.A(n_8265),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_8265),
.Y(n_8870)
);

INVx2_ASAP7_75t_L g8871 ( 
.A(n_8741),
.Y(n_8871)
);

INVx2_ASAP7_75t_L g8872 ( 
.A(n_8741),
.Y(n_8872)
);

INVx2_ASAP7_75t_SL g8873 ( 
.A(n_7863),
.Y(n_8873)
);

INVx2_ASAP7_75t_L g8874 ( 
.A(n_8741),
.Y(n_8874)
);

INVx2_ASAP7_75t_L g8875 ( 
.A(n_7965),
.Y(n_8875)
);

INVx2_ASAP7_75t_L g8876 ( 
.A(n_7965),
.Y(n_8876)
);

INVx2_ASAP7_75t_L g8877 ( 
.A(n_7965),
.Y(n_8877)
);

INVx3_ASAP7_75t_L g8878 ( 
.A(n_7863),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_7831),
.Y(n_8879)
);

INVx1_ASAP7_75t_L g8880 ( 
.A(n_7831),
.Y(n_8880)
);

CKINVDCx20_ASAP7_75t_R g8881 ( 
.A(n_8163),
.Y(n_8881)
);

AND2x4_ASAP7_75t_L g8882 ( 
.A(n_7946),
.B(n_7092),
.Y(n_8882)
);

BUFx2_ASAP7_75t_SL g8883 ( 
.A(n_8135),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_7836),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_7836),
.Y(n_8885)
);

INVx4_ASAP7_75t_L g8886 ( 
.A(n_7973),
.Y(n_8886)
);

INVx2_ASAP7_75t_L g8887 ( 
.A(n_7995),
.Y(n_8887)
);

AOI22xp33_ASAP7_75t_L g8888 ( 
.A1(n_8186),
.A2(n_7136),
.B1(n_6988),
.B2(n_7041),
.Y(n_8888)
);

INVx2_ASAP7_75t_L g8889 ( 
.A(n_7995),
.Y(n_8889)
);

OA21x2_ASAP7_75t_L g8890 ( 
.A1(n_8290),
.A2(n_8507),
.B(n_8401),
.Y(n_8890)
);

OAI21xp5_ASAP7_75t_L g8891 ( 
.A1(n_8471),
.A2(n_8159),
.B(n_7880),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_7837),
.Y(n_8892)
);

BUFx2_ASAP7_75t_L g8893 ( 
.A(n_7884),
.Y(n_8893)
);

INVx2_ASAP7_75t_SL g8894 ( 
.A(n_7863),
.Y(n_8894)
);

INVx1_ASAP7_75t_L g8895 ( 
.A(n_7837),
.Y(n_8895)
);

INVx2_ASAP7_75t_L g8896 ( 
.A(n_7995),
.Y(n_8896)
);

INVx1_ASAP7_75t_L g8897 ( 
.A(n_7842),
.Y(n_8897)
);

INVx1_ASAP7_75t_L g8898 ( 
.A(n_7842),
.Y(n_8898)
);

INVx1_ASAP7_75t_L g8899 ( 
.A(n_7846),
.Y(n_8899)
);

INVx8_ASAP7_75t_L g8900 ( 
.A(n_8040),
.Y(n_8900)
);

INVx3_ASAP7_75t_L g8901 ( 
.A(n_7863),
.Y(n_8901)
);

INVx1_ASAP7_75t_L g8902 ( 
.A(n_7846),
.Y(n_8902)
);

AND2x2_ASAP7_75t_L g8903 ( 
.A(n_7900),
.B(n_7016),
.Y(n_8903)
);

INVx2_ASAP7_75t_L g8904 ( 
.A(n_8044),
.Y(n_8904)
);

INVx1_ASAP7_75t_L g8905 ( 
.A(n_7848),
.Y(n_8905)
);

INVx2_ASAP7_75t_L g8906 ( 
.A(n_8044),
.Y(n_8906)
);

OAI21x1_ASAP7_75t_L g8907 ( 
.A1(n_8745),
.A2(n_7063),
.B(n_6968),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8044),
.Y(n_8908)
);

OR2x2_ASAP7_75t_L g8909 ( 
.A(n_8699),
.B(n_7483),
.Y(n_8909)
);

AO21x2_ASAP7_75t_L g8910 ( 
.A1(n_8671),
.A2(n_7760),
.B(n_6773),
.Y(n_8910)
);

AOI21x1_ASAP7_75t_L g8911 ( 
.A1(n_8752),
.A2(n_7157),
.B(n_7108),
.Y(n_8911)
);

INVx1_ASAP7_75t_L g8912 ( 
.A(n_7848),
.Y(n_8912)
);

AOI21xp5_ASAP7_75t_L g8913 ( 
.A1(n_7841),
.A2(n_8186),
.B(n_7880),
.Y(n_8913)
);

INVx2_ASAP7_75t_L g8914 ( 
.A(n_8118),
.Y(n_8914)
);

AND2x2_ASAP7_75t_L g8915 ( 
.A(n_7900),
.B(n_7016),
.Y(n_8915)
);

HB1xp67_ASAP7_75t_L g8916 ( 
.A(n_8527),
.Y(n_8916)
);

AOI21x1_ASAP7_75t_L g8917 ( 
.A1(n_8752),
.A2(n_7157),
.B(n_7108),
.Y(n_8917)
);

AND2x2_ASAP7_75t_L g8918 ( 
.A(n_7992),
.B(n_7275),
.Y(n_8918)
);

INVx2_ASAP7_75t_SL g8919 ( 
.A(n_8737),
.Y(n_8919)
);

BUFx2_ASAP7_75t_L g8920 ( 
.A(n_7992),
.Y(n_8920)
);

AND2x2_ASAP7_75t_L g8921 ( 
.A(n_7992),
.B(n_7275),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_7850),
.Y(n_8922)
);

HB1xp67_ASAP7_75t_L g8923 ( 
.A(n_8527),
.Y(n_8923)
);

BUFx2_ASAP7_75t_L g8924 ( 
.A(n_8025),
.Y(n_8924)
);

INVx2_ASAP7_75t_SL g8925 ( 
.A(n_8737),
.Y(n_8925)
);

OR2x2_ASAP7_75t_L g8926 ( 
.A(n_8705),
.B(n_6813),
.Y(n_8926)
);

INVx2_ASAP7_75t_L g8927 ( 
.A(n_8118),
.Y(n_8927)
);

BUFx2_ASAP7_75t_L g8928 ( 
.A(n_8025),
.Y(n_8928)
);

OA21x2_ASAP7_75t_L g8929 ( 
.A1(n_8401),
.A2(n_8301),
.B(n_8671),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_7850),
.Y(n_8930)
);

INVx1_ASAP7_75t_L g8931 ( 
.A(n_7855),
.Y(n_8931)
);

INVx3_ASAP7_75t_L g8932 ( 
.A(n_8007),
.Y(n_8932)
);

BUFx3_ASAP7_75t_L g8933 ( 
.A(n_8245),
.Y(n_8933)
);

AO21x2_ASAP7_75t_L g8934 ( 
.A1(n_8671),
.A2(n_6773),
.B(n_6906),
.Y(n_8934)
);

INVx2_ASAP7_75t_L g8935 ( 
.A(n_8118),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_7855),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_7856),
.Y(n_8937)
);

INVx2_ASAP7_75t_L g8938 ( 
.A(n_8124),
.Y(n_8938)
);

INVx2_ASAP7_75t_SL g8939 ( 
.A(n_8737),
.Y(n_8939)
);

BUFx2_ASAP7_75t_SL g8940 ( 
.A(n_8135),
.Y(n_8940)
);

NAND2xp5_ASAP7_75t_L g8941 ( 
.A(n_7799),
.B(n_7287),
.Y(n_8941)
);

INVx2_ASAP7_75t_L g8942 ( 
.A(n_8124),
.Y(n_8942)
);

NAND2xp5_ASAP7_75t_L g8943 ( 
.A(n_7824),
.B(n_7287),
.Y(n_8943)
);

INVx1_ASAP7_75t_L g8944 ( 
.A(n_7856),
.Y(n_8944)
);

AND2x2_ASAP7_75t_L g8945 ( 
.A(n_8025),
.B(n_7253),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_7860),
.Y(n_8946)
);

HB1xp67_ASAP7_75t_L g8947 ( 
.A(n_8606),
.Y(n_8947)
);

AND2x2_ASAP7_75t_L g8948 ( 
.A(n_8027),
.B(n_7253),
.Y(n_8948)
);

BUFx3_ASAP7_75t_L g8949 ( 
.A(n_8245),
.Y(n_8949)
);

INVx2_ASAP7_75t_L g8950 ( 
.A(n_8124),
.Y(n_8950)
);

INVx2_ASAP7_75t_L g8951 ( 
.A(n_8129),
.Y(n_8951)
);

AOI22xp33_ASAP7_75t_L g8952 ( 
.A1(n_8186),
.A2(n_7026),
.B1(n_7055),
.B2(n_7041),
.Y(n_8952)
);

AND2x2_ASAP7_75t_L g8953 ( 
.A(n_8027),
.B(n_7253),
.Y(n_8953)
);

INVx3_ASAP7_75t_L g8954 ( 
.A(n_8007),
.Y(n_8954)
);

OR2x2_ASAP7_75t_L g8955 ( 
.A(n_8705),
.B(n_6813),
.Y(n_8955)
);

INVx1_ASAP7_75t_L g8956 ( 
.A(n_7860),
.Y(n_8956)
);

BUFx2_ASAP7_75t_L g8957 ( 
.A(n_8027),
.Y(n_8957)
);

INVx2_ASAP7_75t_L g8958 ( 
.A(n_8129),
.Y(n_8958)
);

INVx1_ASAP7_75t_L g8959 ( 
.A(n_7862),
.Y(n_8959)
);

INVx2_ASAP7_75t_L g8960 ( 
.A(n_8129),
.Y(n_8960)
);

INVx2_ASAP7_75t_L g8961 ( 
.A(n_8141),
.Y(n_8961)
);

BUFx12f_ASAP7_75t_L g8962 ( 
.A(n_8569),
.Y(n_8962)
);

INVx2_ASAP7_75t_L g8963 ( 
.A(n_8141),
.Y(n_8963)
);

HB1xp67_ASAP7_75t_L g8964 ( 
.A(n_8606),
.Y(n_8964)
);

OAI21x1_ASAP7_75t_L g8965 ( 
.A1(n_8745),
.A2(n_7063),
.B(n_6968),
.Y(n_8965)
);

INVx1_ASAP7_75t_L g8966 ( 
.A(n_7862),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_7824),
.B(n_7443),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_7864),
.Y(n_8968)
);

INVx2_ASAP7_75t_L g8969 ( 
.A(n_8141),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_7864),
.Y(n_8970)
);

INVx1_ASAP7_75t_L g8971 ( 
.A(n_7867),
.Y(n_8971)
);

AND2x2_ASAP7_75t_L g8972 ( 
.A(n_8030),
.B(n_7253),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_7867),
.Y(n_8973)
);

INVx1_ASAP7_75t_L g8974 ( 
.A(n_7888),
.Y(n_8974)
);

NAND2xp5_ASAP7_75t_L g8975 ( 
.A(n_7945),
.B(n_7443),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_7888),
.Y(n_8976)
);

INVx1_ASAP7_75t_L g8977 ( 
.A(n_7898),
.Y(n_8977)
);

INVx3_ASAP7_75t_L g8978 ( 
.A(n_8022),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_7898),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_7906),
.Y(n_8980)
);

AND2x2_ASAP7_75t_L g8981 ( 
.A(n_8030),
.B(n_7398),
.Y(n_8981)
);

AND2x2_ASAP7_75t_L g8982 ( 
.A(n_8030),
.B(n_7398),
.Y(n_8982)
);

OR2x6_ASAP7_75t_L g8983 ( 
.A(n_7858),
.B(n_6818),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_7906),
.Y(n_8984)
);

INVx2_ASAP7_75t_L g8985 ( 
.A(n_8153),
.Y(n_8985)
);

INVx2_ASAP7_75t_L g8986 ( 
.A(n_8153),
.Y(n_8986)
);

INVx2_ASAP7_75t_L g8987 ( 
.A(n_8153),
.Y(n_8987)
);

INVx2_ASAP7_75t_SL g8988 ( 
.A(n_8737),
.Y(n_8988)
);

INVx1_ASAP7_75t_L g8989 ( 
.A(n_7907),
.Y(n_8989)
);

CKINVDCx12_ASAP7_75t_R g8990 ( 
.A(n_8041),
.Y(n_8990)
);

BUFx2_ASAP7_75t_L g8991 ( 
.A(n_8042),
.Y(n_8991)
);

HB1xp67_ASAP7_75t_L g8992 ( 
.A(n_7812),
.Y(n_8992)
);

OAI21x1_ASAP7_75t_L g8993 ( 
.A1(n_8694),
.A2(n_7063),
.B(n_6968),
.Y(n_8993)
);

INVx1_ASAP7_75t_L g8994 ( 
.A(n_7907),
.Y(n_8994)
);

OR2x2_ASAP7_75t_L g8995 ( 
.A(n_8719),
.B(n_7954),
.Y(n_8995)
);

HB1xp67_ASAP7_75t_L g8996 ( 
.A(n_7812),
.Y(n_8996)
);

INVx1_ASAP7_75t_L g8997 ( 
.A(n_7908),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_7908),
.Y(n_8998)
);

INVx2_ASAP7_75t_L g8999 ( 
.A(n_8165),
.Y(n_8999)
);

HB1xp67_ASAP7_75t_L g9000 ( 
.A(n_7823),
.Y(n_9000)
);

INVx2_ASAP7_75t_L g9001 ( 
.A(n_8165),
.Y(n_9001)
);

INVx1_ASAP7_75t_L g9002 ( 
.A(n_7910),
.Y(n_9002)
);

AND2x2_ASAP7_75t_L g9003 ( 
.A(n_8042),
.B(n_7398),
.Y(n_9003)
);

INVx1_ASAP7_75t_L g9004 ( 
.A(n_7910),
.Y(n_9004)
);

INVx1_ASAP7_75t_L g9005 ( 
.A(n_7912),
.Y(n_9005)
);

INVx2_ASAP7_75t_SL g9006 ( 
.A(n_8737),
.Y(n_9006)
);

NOR2x1_ASAP7_75t_R g9007 ( 
.A(n_8245),
.B(n_7053),
.Y(n_9007)
);

INVx2_ASAP7_75t_L g9008 ( 
.A(n_8165),
.Y(n_9008)
);

AO21x2_ASAP7_75t_L g9009 ( 
.A1(n_8131),
.A2(n_6906),
.B(n_7707),
.Y(n_9009)
);

INVx2_ASAP7_75t_L g9010 ( 
.A(n_8179),
.Y(n_9010)
);

INVx2_ASAP7_75t_L g9011 ( 
.A(n_8179),
.Y(n_9011)
);

HB1xp67_ASAP7_75t_L g9012 ( 
.A(n_7823),
.Y(n_9012)
);

INVx2_ASAP7_75t_L g9013 ( 
.A(n_8179),
.Y(n_9013)
);

BUFx3_ASAP7_75t_L g9014 ( 
.A(n_8292),
.Y(n_9014)
);

INVx2_ASAP7_75t_L g9015 ( 
.A(n_7868),
.Y(n_9015)
);

INVx2_ASAP7_75t_L g9016 ( 
.A(n_7868),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_7912),
.Y(n_9017)
);

BUFx4f_ASAP7_75t_SL g9018 ( 
.A(n_8163),
.Y(n_9018)
);

INVx1_ASAP7_75t_L g9019 ( 
.A(n_7918),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_7918),
.Y(n_9020)
);

INVx2_ASAP7_75t_L g9021 ( 
.A(n_7868),
.Y(n_9021)
);

INVx1_ASAP7_75t_L g9022 ( 
.A(n_8072),
.Y(n_9022)
);

OR2x2_ASAP7_75t_L g9023 ( 
.A(n_8719),
.B(n_7954),
.Y(n_9023)
);

INVx1_ASAP7_75t_L g9024 ( 
.A(n_8072),
.Y(n_9024)
);

INVx1_ASAP7_75t_L g9025 ( 
.A(n_8075),
.Y(n_9025)
);

INVx2_ASAP7_75t_SL g9026 ( 
.A(n_8737),
.Y(n_9026)
);

BUFx2_ASAP7_75t_L g9027 ( 
.A(n_8042),
.Y(n_9027)
);

OA21x2_ASAP7_75t_L g9028 ( 
.A1(n_8301),
.A2(n_7805),
.B(n_7795),
.Y(n_9028)
);

OAI21x1_ASAP7_75t_L g9029 ( 
.A1(n_8694),
.A2(n_7152),
.B(n_7079),
.Y(n_9029)
);

AND2x2_ASAP7_75t_L g9030 ( 
.A(n_8050),
.B(n_8104),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_8075),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8083),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_8083),
.Y(n_9033)
);

AND2x2_ASAP7_75t_L g9034 ( 
.A(n_8050),
.B(n_7398),
.Y(n_9034)
);

OAI21xp5_ASAP7_75t_L g9035 ( 
.A1(n_8159),
.A2(n_6987),
.B(n_6982),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_8096),
.Y(n_9036)
);

INVx2_ASAP7_75t_L g9037 ( 
.A(n_7894),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_8096),
.Y(n_9038)
);

NAND2x1_ASAP7_75t_L g9039 ( 
.A(n_7807),
.B(n_7587),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_8146),
.Y(n_9040)
);

INVx2_ASAP7_75t_L g9041 ( 
.A(n_7894),
.Y(n_9041)
);

AO21x2_ASAP7_75t_L g9042 ( 
.A1(n_8131),
.A2(n_7707),
.B(n_7145),
.Y(n_9042)
);

AND2x4_ASAP7_75t_L g9043 ( 
.A(n_7946),
.B(n_7092),
.Y(n_9043)
);

INVx2_ASAP7_75t_L g9044 ( 
.A(n_7894),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_8146),
.Y(n_9045)
);

INVx1_ASAP7_75t_L g9046 ( 
.A(n_8187),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8187),
.Y(n_9047)
);

INVx1_ASAP7_75t_L g9048 ( 
.A(n_8262),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_7943),
.Y(n_9049)
);

OR2x2_ASAP7_75t_L g9050 ( 
.A(n_8049),
.B(n_7549),
.Y(n_9050)
);

HB1xp67_ASAP7_75t_L g9051 ( 
.A(n_7881),
.Y(n_9051)
);

BUFx2_ASAP7_75t_SL g9052 ( 
.A(n_8737),
.Y(n_9052)
);

OR2x2_ASAP7_75t_L g9053 ( 
.A(n_8049),
.B(n_8253),
.Y(n_9053)
);

INVx1_ASAP7_75t_L g9054 ( 
.A(n_8262),
.Y(n_9054)
);

INVx1_ASAP7_75t_L g9055 ( 
.A(n_8269),
.Y(n_9055)
);

OR2x6_ASAP7_75t_L g9056 ( 
.A(n_7858),
.B(n_6818),
.Y(n_9056)
);

OR2x2_ASAP7_75t_L g9057 ( 
.A(n_8253),
.B(n_7566),
.Y(n_9057)
);

INVx2_ASAP7_75t_L g9058 ( 
.A(n_7943),
.Y(n_9058)
);

AND2x2_ASAP7_75t_L g9059 ( 
.A(n_8050),
.B(n_7432),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_8269),
.Y(n_9060)
);

AND2x2_ASAP7_75t_L g9061 ( 
.A(n_8104),
.B(n_7432),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8276),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_8276),
.Y(n_9063)
);

INVx1_ASAP7_75t_L g9064 ( 
.A(n_8279),
.Y(n_9064)
);

HB1xp67_ASAP7_75t_L g9065 ( 
.A(n_7881),
.Y(n_9065)
);

INVx2_ASAP7_75t_SL g9066 ( 
.A(n_7973),
.Y(n_9066)
);

BUFx4f_ASAP7_75t_SL g9067 ( 
.A(n_7952),
.Y(n_9067)
);

HB1xp67_ASAP7_75t_L g9068 ( 
.A(n_7882),
.Y(n_9068)
);

AND2x2_ASAP7_75t_L g9069 ( 
.A(n_8104),
.B(n_7432),
.Y(n_9069)
);

AOI22xp33_ASAP7_75t_L g9070 ( 
.A1(n_8094),
.A2(n_7026),
.B1(n_7057),
.B2(n_7055),
.Y(n_9070)
);

HB1xp67_ASAP7_75t_SL g9071 ( 
.A(n_8212),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8279),
.Y(n_9072)
);

INVx2_ASAP7_75t_L g9073 ( 
.A(n_7943),
.Y(n_9073)
);

INVx2_ASAP7_75t_SL g9074 ( 
.A(n_7973),
.Y(n_9074)
);

INVx2_ASAP7_75t_L g9075 ( 
.A(n_7794),
.Y(n_9075)
);

INVx1_ASAP7_75t_L g9076 ( 
.A(n_8297),
.Y(n_9076)
);

INVx1_ASAP7_75t_L g9077 ( 
.A(n_8297),
.Y(n_9077)
);

INVx2_ASAP7_75t_L g9078 ( 
.A(n_7794),
.Y(n_9078)
);

INVx2_ASAP7_75t_L g9079 ( 
.A(n_7794),
.Y(n_9079)
);

OR2x2_ASAP7_75t_L g9080 ( 
.A(n_8260),
.B(n_7566),
.Y(n_9080)
);

INVx2_ASAP7_75t_L g9081 ( 
.A(n_7803),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_8336),
.Y(n_9082)
);

HB1xp67_ASAP7_75t_L g9083 ( 
.A(n_7882),
.Y(n_9083)
);

OAI21x1_ASAP7_75t_L g9084 ( 
.A1(n_8760),
.A2(n_8498),
.B(n_8492),
.Y(n_9084)
);

HB1xp67_ASAP7_75t_L g9085 ( 
.A(n_7897),
.Y(n_9085)
);

AO31x2_ASAP7_75t_L g9086 ( 
.A1(n_8509),
.A2(n_8544),
.A3(n_8430),
.B(n_8752),
.Y(n_9086)
);

INVxp67_ASAP7_75t_L g9087 ( 
.A(n_8106),
.Y(n_9087)
);

INVx2_ASAP7_75t_L g9088 ( 
.A(n_7803),
.Y(n_9088)
);

INVxp67_ASAP7_75t_SL g9089 ( 
.A(n_7807),
.Y(n_9089)
);

NAND2xp5_ASAP7_75t_L g9090 ( 
.A(n_7945),
.B(n_6930),
.Y(n_9090)
);

AOI22xp33_ASAP7_75t_L g9091 ( 
.A1(n_8094),
.A2(n_7057),
.B1(n_7089),
.B2(n_6898),
.Y(n_9091)
);

INVx2_ASAP7_75t_SL g9092 ( 
.A(n_7833),
.Y(n_9092)
);

INVx1_ASAP7_75t_L g9093 ( 
.A(n_8336),
.Y(n_9093)
);

INVx1_ASAP7_75t_L g9094 ( 
.A(n_8341),
.Y(n_9094)
);

BUFx3_ASAP7_75t_L g9095 ( 
.A(n_8292),
.Y(n_9095)
);

INVx1_ASAP7_75t_L g9096 ( 
.A(n_8341),
.Y(n_9096)
);

INVx3_ASAP7_75t_L g9097 ( 
.A(n_8022),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8366),
.Y(n_9098)
);

INVx2_ASAP7_75t_SL g9099 ( 
.A(n_7833),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8366),
.Y(n_9100)
);

OAI21xp5_ASAP7_75t_L g9101 ( 
.A1(n_7841),
.A2(n_6982),
.B(n_7222),
.Y(n_9101)
);

NOR2xp33_ASAP7_75t_L g9102 ( 
.A(n_8648),
.B(n_6739),
.Y(n_9102)
);

INVx1_ASAP7_75t_L g9103 ( 
.A(n_8381),
.Y(n_9103)
);

INVx2_ASAP7_75t_L g9104 ( 
.A(n_7803),
.Y(n_9104)
);

CKINVDCx5p33_ASAP7_75t_R g9105 ( 
.A(n_8087),
.Y(n_9105)
);

CKINVDCx5p33_ASAP7_75t_R g9106 ( 
.A(n_8087),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_8381),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_8395),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_8395),
.Y(n_9109)
);

INVx2_ASAP7_75t_L g9110 ( 
.A(n_7808),
.Y(n_9110)
);

OR2x2_ASAP7_75t_L g9111 ( 
.A(n_8260),
.B(n_7591),
.Y(n_9111)
);

BUFx2_ASAP7_75t_L g9112 ( 
.A(n_8111),
.Y(n_9112)
);

INVx1_ASAP7_75t_L g9113 ( 
.A(n_8398),
.Y(n_9113)
);

INVx1_ASAP7_75t_L g9114 ( 
.A(n_8398),
.Y(n_9114)
);

BUFx3_ASAP7_75t_L g9115 ( 
.A(n_8292),
.Y(n_9115)
);

NAND2xp5_ASAP7_75t_L g9116 ( 
.A(n_7852),
.B(n_6930),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_L g9117 ( 
.A(n_7852),
.B(n_8149),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8412),
.Y(n_9118)
);

OR2x2_ASAP7_75t_L g9119 ( 
.A(n_7877),
.B(n_7591),
.Y(n_9119)
);

BUFx6f_ASAP7_75t_SL g9120 ( 
.A(n_7833),
.Y(n_9120)
);

INVx1_ASAP7_75t_L g9121 ( 
.A(n_8412),
.Y(n_9121)
);

AND2x2_ASAP7_75t_L g9122 ( 
.A(n_8111),
.B(n_7432),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_7808),
.Y(n_9123)
);

INVx1_ASAP7_75t_L g9124 ( 
.A(n_8441),
.Y(n_9124)
);

HB1xp67_ASAP7_75t_L g9125 ( 
.A(n_7897),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_8441),
.Y(n_9126)
);

INVx2_ASAP7_75t_L g9127 ( 
.A(n_7808),
.Y(n_9127)
);

BUFx3_ASAP7_75t_L g9128 ( 
.A(n_8415),
.Y(n_9128)
);

OAI21x1_ASAP7_75t_L g9129 ( 
.A1(n_8760),
.A2(n_7152),
.B(n_7079),
.Y(n_9129)
);

INVx1_ASAP7_75t_L g9130 ( 
.A(n_8473),
.Y(n_9130)
);

INVx1_ASAP7_75t_L g9131 ( 
.A(n_8473),
.Y(n_9131)
);

HB1xp67_ASAP7_75t_L g9132 ( 
.A(n_7902),
.Y(n_9132)
);

INVx2_ASAP7_75t_L g9133 ( 
.A(n_7813),
.Y(n_9133)
);

INVx2_ASAP7_75t_L g9134 ( 
.A(n_7813),
.Y(n_9134)
);

INVx1_ASAP7_75t_L g9135 ( 
.A(n_8476),
.Y(n_9135)
);

INVx8_ASAP7_75t_L g9136 ( 
.A(n_8415),
.Y(n_9136)
);

INVx11_ASAP7_75t_L g9137 ( 
.A(n_8415),
.Y(n_9137)
);

AO21x2_ASAP7_75t_L g9138 ( 
.A1(n_8131),
.A2(n_7930),
.B(n_8436),
.Y(n_9138)
);

BUFx6f_ASAP7_75t_L g9139 ( 
.A(n_7851),
.Y(n_9139)
);

INVx1_ASAP7_75t_L g9140 ( 
.A(n_8476),
.Y(n_9140)
);

OR2x6_ASAP7_75t_L g9141 ( 
.A(n_7874),
.B(n_6818),
.Y(n_9141)
);

INVx2_ASAP7_75t_L g9142 ( 
.A(n_7813),
.Y(n_9142)
);

INVx2_ASAP7_75t_L g9143 ( 
.A(n_7815),
.Y(n_9143)
);

OAI21x1_ASAP7_75t_L g9144 ( 
.A1(n_8492),
.A2(n_7152),
.B(n_7079),
.Y(n_9144)
);

INVx2_ASAP7_75t_SL g9145 ( 
.A(n_7851),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_7815),
.Y(n_9146)
);

INVx2_ASAP7_75t_L g9147 ( 
.A(n_7815),
.Y(n_9147)
);

INVx2_ASAP7_75t_L g9148 ( 
.A(n_7819),
.Y(n_9148)
);

INVx1_ASAP7_75t_L g9149 ( 
.A(n_8479),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_8479),
.Y(n_9150)
);

AND2x4_ASAP7_75t_L g9151 ( 
.A(n_7946),
.B(n_7092),
.Y(n_9151)
);

BUFx2_ASAP7_75t_L g9152 ( 
.A(n_8111),
.Y(n_9152)
);

AOI21xp5_ASAP7_75t_SL g9153 ( 
.A1(n_7825),
.A2(n_6749),
.B(n_6732),
.Y(n_9153)
);

INVxp67_ASAP7_75t_SL g9154 ( 
.A(n_7807),
.Y(n_9154)
);

AND2x2_ASAP7_75t_L g9155 ( 
.A(n_8231),
.B(n_7448),
.Y(n_9155)
);

BUFx2_ASAP7_75t_L g9156 ( 
.A(n_8231),
.Y(n_9156)
);

INVx2_ASAP7_75t_L g9157 ( 
.A(n_7819),
.Y(n_9157)
);

OR2x2_ASAP7_75t_L g9158 ( 
.A(n_7877),
.B(n_6977),
.Y(n_9158)
);

INVx1_ASAP7_75t_L g9159 ( 
.A(n_8483),
.Y(n_9159)
);

INVx1_ASAP7_75t_L g9160 ( 
.A(n_8483),
.Y(n_9160)
);

BUFx2_ASAP7_75t_L g9161 ( 
.A(n_8231),
.Y(n_9161)
);

INVx2_ASAP7_75t_L g9162 ( 
.A(n_7819),
.Y(n_9162)
);

OR2x2_ASAP7_75t_L g9163 ( 
.A(n_8591),
.B(n_7879),
.Y(n_9163)
);

OR2x2_ASAP7_75t_L g9164 ( 
.A(n_8591),
.B(n_6977),
.Y(n_9164)
);

INVx1_ASAP7_75t_L g9165 ( 
.A(n_8508),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_7843),
.Y(n_9166)
);

INVx1_ASAP7_75t_L g9167 ( 
.A(n_8508),
.Y(n_9167)
);

INVxp67_ASAP7_75t_SL g9168 ( 
.A(n_7845),
.Y(n_9168)
);

AND2x2_ASAP7_75t_L g9169 ( 
.A(n_8248),
.B(n_7448),
.Y(n_9169)
);

AND2x2_ASAP7_75t_L g9170 ( 
.A(n_8248),
.B(n_7448),
.Y(n_9170)
);

BUFx6f_ASAP7_75t_L g9171 ( 
.A(n_7851),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_8513),
.Y(n_9172)
);

OA21x2_ASAP7_75t_L g9173 ( 
.A1(n_7795),
.A2(n_6509),
.B(n_6501),
.Y(n_9173)
);

INVx1_ASAP7_75t_L g9174 ( 
.A(n_8513),
.Y(n_9174)
);

AO21x2_ASAP7_75t_L g9175 ( 
.A1(n_7930),
.A2(n_7145),
.B(n_7573),
.Y(n_9175)
);

HB1xp67_ASAP7_75t_L g9176 ( 
.A(n_7902),
.Y(n_9176)
);

OAI21xp5_ASAP7_75t_L g9177 ( 
.A1(n_7972),
.A2(n_7222),
.B(n_6940),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_8542),
.Y(n_9178)
);

INVx1_ASAP7_75t_L g9179 ( 
.A(n_8542),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_7843),
.Y(n_9180)
);

INVx1_ASAP7_75t_L g9181 ( 
.A(n_8550),
.Y(n_9181)
);

NAND2x1p5_ASAP7_75t_L g9182 ( 
.A(n_8792),
.B(n_7083),
.Y(n_9182)
);

INVx3_ASAP7_75t_L g9183 ( 
.A(n_8066),
.Y(n_9183)
);

INVx1_ASAP7_75t_L g9184 ( 
.A(n_8550),
.Y(n_9184)
);

BUFx2_ASAP7_75t_L g9185 ( 
.A(n_8248),
.Y(n_9185)
);

INVx3_ASAP7_75t_L g9186 ( 
.A(n_8066),
.Y(n_9186)
);

INVx2_ASAP7_75t_L g9187 ( 
.A(n_7843),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_8579),
.Y(n_9188)
);

INVx2_ASAP7_75t_L g9189 ( 
.A(n_7849),
.Y(n_9189)
);

INVx2_ASAP7_75t_L g9190 ( 
.A(n_7849),
.Y(n_9190)
);

INVx1_ASAP7_75t_L g9191 ( 
.A(n_8579),
.Y(n_9191)
);

INVx1_ASAP7_75t_L g9192 ( 
.A(n_8586),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_8149),
.B(n_7013),
.Y(n_9193)
);

OR2x2_ASAP7_75t_L g9194 ( 
.A(n_7879),
.B(n_7013),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_8586),
.Y(n_9195)
);

CKINVDCx5p33_ASAP7_75t_R g9196 ( 
.A(n_8212),
.Y(n_9196)
);

INVx2_ASAP7_75t_L g9197 ( 
.A(n_7849),
.Y(n_9197)
);

AND2x2_ASAP7_75t_L g9198 ( 
.A(n_8317),
.B(n_7448),
.Y(n_9198)
);

INVx2_ASAP7_75t_SL g9199 ( 
.A(n_7876),
.Y(n_9199)
);

BUFx2_ASAP7_75t_L g9200 ( 
.A(n_8317),
.Y(n_9200)
);

INVx1_ASAP7_75t_L g9201 ( 
.A(n_8587),
.Y(n_9201)
);

OR2x6_ASAP7_75t_L g9202 ( 
.A(n_7874),
.B(n_6818),
.Y(n_9202)
);

INVx2_ASAP7_75t_L g9203 ( 
.A(n_7853),
.Y(n_9203)
);

AND2x4_ASAP7_75t_L g9204 ( 
.A(n_7946),
.B(n_7092),
.Y(n_9204)
);

INVx2_ASAP7_75t_SL g9205 ( 
.A(n_7876),
.Y(n_9205)
);

AO21x2_ASAP7_75t_L g9206 ( 
.A1(n_7930),
.A2(n_7573),
.B(n_7596),
.Y(n_9206)
);

INVxp67_ASAP7_75t_L g9207 ( 
.A(n_8138),
.Y(n_9207)
);

INVx1_ASAP7_75t_L g9208 ( 
.A(n_8587),
.Y(n_9208)
);

OAI21x1_ASAP7_75t_L g9209 ( 
.A1(n_8492),
.A2(n_7152),
.B(n_7079),
.Y(n_9209)
);

AND2x2_ASAP7_75t_L g9210 ( 
.A(n_8317),
.B(n_7463),
.Y(n_9210)
);

AND2x4_ASAP7_75t_L g9211 ( 
.A(n_7946),
.B(n_7141),
.Y(n_9211)
);

INVx1_ASAP7_75t_L g9212 ( 
.A(n_8595),
.Y(n_9212)
);

AO21x2_ASAP7_75t_L g9213 ( 
.A1(n_8436),
.A2(n_7598),
.B(n_7596),
.Y(n_9213)
);

AND2x2_ASAP7_75t_L g9214 ( 
.A(n_8509),
.B(n_8544),
.Y(n_9214)
);

INVx2_ASAP7_75t_SL g9215 ( 
.A(n_7876),
.Y(n_9215)
);

BUFx12f_ASAP7_75t_L g9216 ( 
.A(n_8569),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_8595),
.Y(n_9217)
);

BUFx2_ASAP7_75t_L g9218 ( 
.A(n_8041),
.Y(n_9218)
);

INVx3_ASAP7_75t_L g9219 ( 
.A(n_8099),
.Y(n_9219)
);

INVx1_ASAP7_75t_L g9220 ( 
.A(n_8612),
.Y(n_9220)
);

INVx2_ASAP7_75t_L g9221 ( 
.A(n_7853),
.Y(n_9221)
);

AO21x2_ASAP7_75t_L g9222 ( 
.A1(n_7839),
.A2(n_7598),
.B(n_7310),
.Y(n_9222)
);

NAND2x1_ASAP7_75t_L g9223 ( 
.A(n_7845),
.B(n_7594),
.Y(n_9223)
);

OA21x2_ASAP7_75t_L g9224 ( 
.A1(n_7795),
.A2(n_6509),
.B(n_7144),
.Y(n_9224)
);

AND2x2_ASAP7_75t_L g9225 ( 
.A(n_8509),
.B(n_7463),
.Y(n_9225)
);

BUFx2_ASAP7_75t_L g9226 ( 
.A(n_8544),
.Y(n_9226)
);

INVx2_ASAP7_75t_SL g9227 ( 
.A(n_7925),
.Y(n_9227)
);

INVx2_ASAP7_75t_L g9228 ( 
.A(n_7853),
.Y(n_9228)
);

NAND3xp33_ASAP7_75t_L g9229 ( 
.A(n_7825),
.B(n_7186),
.C(n_7205),
.Y(n_9229)
);

INVx2_ASAP7_75t_L g9230 ( 
.A(n_7854),
.Y(n_9230)
);

BUFx3_ASAP7_75t_L g9231 ( 
.A(n_8757),
.Y(n_9231)
);

INVx3_ASAP7_75t_SL g9232 ( 
.A(n_7909),
.Y(n_9232)
);

INVx2_ASAP7_75t_L g9233 ( 
.A(n_7854),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8612),
.Y(n_9234)
);

HB1xp67_ASAP7_75t_L g9235 ( 
.A(n_7933),
.Y(n_9235)
);

INVx2_ASAP7_75t_L g9236 ( 
.A(n_7854),
.Y(n_9236)
);

INVx1_ASAP7_75t_L g9237 ( 
.A(n_8674),
.Y(n_9237)
);

HB1xp67_ASAP7_75t_L g9238 ( 
.A(n_7933),
.Y(n_9238)
);

BUFx3_ASAP7_75t_L g9239 ( 
.A(n_8757),
.Y(n_9239)
);

NAND2xp5_ASAP7_75t_L g9240 ( 
.A(n_8614),
.B(n_6003),
.Y(n_9240)
);

INVx1_ASAP7_75t_L g9241 ( 
.A(n_8674),
.Y(n_9241)
);

INVx2_ASAP7_75t_L g9242 ( 
.A(n_7859),
.Y(n_9242)
);

HB1xp67_ASAP7_75t_L g9243 ( 
.A(n_7949),
.Y(n_9243)
);

INVx2_ASAP7_75t_L g9244 ( 
.A(n_7859),
.Y(n_9244)
);

AOI21x1_ASAP7_75t_L g9245 ( 
.A1(n_8792),
.A2(n_7716),
.B(n_7678),
.Y(n_9245)
);

INVx2_ASAP7_75t_L g9246 ( 
.A(n_7859),
.Y(n_9246)
);

BUFx6f_ASAP7_75t_L g9247 ( 
.A(n_7925),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_8693),
.Y(n_9248)
);

INVx2_ASAP7_75t_L g9249 ( 
.A(n_7866),
.Y(n_9249)
);

AO21x2_ASAP7_75t_L g9250 ( 
.A1(n_7839),
.A2(n_7310),
.B(n_7283),
.Y(n_9250)
);

AO21x1_ASAP7_75t_SL g9251 ( 
.A1(n_8511),
.A2(n_7552),
.B(n_7550),
.Y(n_9251)
);

INVx1_ASAP7_75t_L g9252 ( 
.A(n_8693),
.Y(n_9252)
);

HB1xp67_ASAP7_75t_L g9253 ( 
.A(n_7949),
.Y(n_9253)
);

NAND2xp33_ASAP7_75t_R g9254 ( 
.A(n_8746),
.B(n_6789),
.Y(n_9254)
);

INVx2_ASAP7_75t_L g9255 ( 
.A(n_7866),
.Y(n_9255)
);

INVx1_ASAP7_75t_L g9256 ( 
.A(n_8710),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_8710),
.Y(n_9257)
);

INVx1_ASAP7_75t_L g9258 ( 
.A(n_8712),
.Y(n_9258)
);

BUFx3_ASAP7_75t_L g9259 ( 
.A(n_8757),
.Y(n_9259)
);

AO21x1_ASAP7_75t_L g9260 ( 
.A1(n_8170),
.A2(n_6739),
.B(n_6743),
.Y(n_9260)
);

INVx1_ASAP7_75t_L g9261 ( 
.A(n_8712),
.Y(n_9261)
);

INVx1_ASAP7_75t_L g9262 ( 
.A(n_8801),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_8801),
.Y(n_9263)
);

INVx1_ASAP7_75t_L g9264 ( 
.A(n_8802),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_8802),
.Y(n_9265)
);

INVx1_ASAP7_75t_L g9266 ( 
.A(n_8811),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_8811),
.Y(n_9267)
);

INVx2_ASAP7_75t_L g9268 ( 
.A(n_7866),
.Y(n_9268)
);

AND2x2_ASAP7_75t_L g9269 ( 
.A(n_7845),
.B(n_7463),
.Y(n_9269)
);

INVxp67_ASAP7_75t_SL g9270 ( 
.A(n_7920),
.Y(n_9270)
);

INVx2_ASAP7_75t_L g9271 ( 
.A(n_7869),
.Y(n_9271)
);

INVx2_ASAP7_75t_L g9272 ( 
.A(n_7869),
.Y(n_9272)
);

AOI21xp5_ASAP7_75t_SL g9273 ( 
.A1(n_7865),
.A2(n_6749),
.B(n_6724),
.Y(n_9273)
);

AOI22xp5_ASAP7_75t_L g9274 ( 
.A1(n_8430),
.A2(n_6824),
.B1(n_6978),
.B2(n_6970),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8813),
.Y(n_9275)
);

INVx4_ASAP7_75t_L g9276 ( 
.A(n_7909),
.Y(n_9276)
);

BUFx2_ASAP7_75t_L g9277 ( 
.A(n_7798),
.Y(n_9277)
);

AO21x2_ASAP7_75t_L g9278 ( 
.A1(n_7839),
.A2(n_7283),
.B(n_6769),
.Y(n_9278)
);

CKINVDCx5p33_ASAP7_75t_R g9279 ( 
.A(n_8458),
.Y(n_9279)
);

AND2x2_ASAP7_75t_L g9280 ( 
.A(n_8355),
.B(n_7463),
.Y(n_9280)
);

INVx1_ASAP7_75t_L g9281 ( 
.A(n_8813),
.Y(n_9281)
);

AOI21x1_ASAP7_75t_L g9282 ( 
.A1(n_8792),
.A2(n_7716),
.B(n_7678),
.Y(n_9282)
);

INVx1_ASAP7_75t_L g9283 ( 
.A(n_7923),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_7923),
.Y(n_9284)
);

HB1xp67_ASAP7_75t_L g9285 ( 
.A(n_7986),
.Y(n_9285)
);

INVxp33_ASAP7_75t_L g9286 ( 
.A(n_8458),
.Y(n_9286)
);

INVx2_ASAP7_75t_SL g9287 ( 
.A(n_7925),
.Y(n_9287)
);

NAND2xp5_ASAP7_75t_L g9288 ( 
.A(n_8614),
.B(n_7200),
.Y(n_9288)
);

INVx1_ASAP7_75t_L g9289 ( 
.A(n_7926),
.Y(n_9289)
);

INVx3_ASAP7_75t_L g9290 ( 
.A(n_8099),
.Y(n_9290)
);

INVx1_ASAP7_75t_L g9291 ( 
.A(n_7926),
.Y(n_9291)
);

AND2x2_ASAP7_75t_L g9292 ( 
.A(n_8355),
.B(n_7470),
.Y(n_9292)
);

OAI21x1_ASAP7_75t_L g9293 ( 
.A1(n_8498),
.A2(n_7297),
.B(n_6697),
.Y(n_9293)
);

INVx1_ASAP7_75t_L g9294 ( 
.A(n_7931),
.Y(n_9294)
);

INVx2_ASAP7_75t_L g9295 ( 
.A(n_7869),
.Y(n_9295)
);

INVx2_ASAP7_75t_L g9296 ( 
.A(n_7870),
.Y(n_9296)
);

AO21x2_ASAP7_75t_L g9297 ( 
.A1(n_7839),
.A2(n_6769),
.B(n_7475),
.Y(n_9297)
);

AND2x2_ASAP7_75t_L g9298 ( 
.A(n_8355),
.B(n_7470),
.Y(n_9298)
);

AND2x2_ASAP7_75t_L g9299 ( 
.A(n_8359),
.B(n_7470),
.Y(n_9299)
);

INVx1_ASAP7_75t_L g9300 ( 
.A(n_7931),
.Y(n_9300)
);

OR2x2_ASAP7_75t_L g9301 ( 
.A(n_7883),
.B(n_7316),
.Y(n_9301)
);

INVx1_ASAP7_75t_L g9302 ( 
.A(n_7935),
.Y(n_9302)
);

OAI21xp33_ASAP7_75t_SL g9303 ( 
.A1(n_7972),
.A2(n_6833),
.B(n_6794),
.Y(n_9303)
);

INVx1_ASAP7_75t_L g9304 ( 
.A(n_7935),
.Y(n_9304)
);

INVx2_ASAP7_75t_L g9305 ( 
.A(n_7870),
.Y(n_9305)
);

CKINVDCx5p33_ASAP7_75t_R g9306 ( 
.A(n_8786),
.Y(n_9306)
);

INVx2_ASAP7_75t_L g9307 ( 
.A(n_7870),
.Y(n_9307)
);

INVx1_ASAP7_75t_L g9308 ( 
.A(n_7936),
.Y(n_9308)
);

INVx2_ASAP7_75t_L g9309 ( 
.A(n_7872),
.Y(n_9309)
);

INVx2_ASAP7_75t_L g9310 ( 
.A(n_7872),
.Y(n_9310)
);

INVx5_ASAP7_75t_L g9311 ( 
.A(n_8786),
.Y(n_9311)
);

OR2x2_ASAP7_75t_L g9312 ( 
.A(n_7883),
.B(n_7316),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_7936),
.Y(n_9313)
);

INVx2_ASAP7_75t_SL g9314 ( 
.A(n_7967),
.Y(n_9314)
);

INVx1_ASAP7_75t_L g9315 ( 
.A(n_7937),
.Y(n_9315)
);

AND2x2_ASAP7_75t_L g9316 ( 
.A(n_8359),
.B(n_7470),
.Y(n_9316)
);

OA21x2_ASAP7_75t_L g9317 ( 
.A1(n_7805),
.A2(n_7169),
.B(n_7166),
.Y(n_9317)
);

INVx1_ASAP7_75t_L g9318 ( 
.A(n_7937),
.Y(n_9318)
);

INVx1_ASAP7_75t_L g9319 ( 
.A(n_7938),
.Y(n_9319)
);

INVx1_ASAP7_75t_L g9320 ( 
.A(n_7938),
.Y(n_9320)
);

INVx2_ASAP7_75t_L g9321 ( 
.A(n_7872),
.Y(n_9321)
);

AND2x2_ASAP7_75t_L g9322 ( 
.A(n_8359),
.B(n_7477),
.Y(n_9322)
);

OR2x6_ASAP7_75t_L g9323 ( 
.A(n_8145),
.B(n_6932),
.Y(n_9323)
);

INVx3_ASAP7_75t_L g9324 ( 
.A(n_7873),
.Y(n_9324)
);

OAI21xp5_ASAP7_75t_L g9325 ( 
.A1(n_7996),
.A2(n_6715),
.B(n_6849),
.Y(n_9325)
);

INVx1_ASAP7_75t_L g9326 ( 
.A(n_7941),
.Y(n_9326)
);

AND2x2_ASAP7_75t_L g9327 ( 
.A(n_8363),
.B(n_7477),
.Y(n_9327)
);

HB1xp67_ASAP7_75t_L g9328 ( 
.A(n_7986),
.Y(n_9328)
);

NOR2x1_ASAP7_75t_SL g9329 ( 
.A(n_8033),
.B(n_7277),
.Y(n_9329)
);

INVx2_ASAP7_75t_L g9330 ( 
.A(n_7878),
.Y(n_9330)
);

INVx1_ASAP7_75t_L g9331 ( 
.A(n_7941),
.Y(n_9331)
);

AOI22xp33_ASAP7_75t_L g9332 ( 
.A1(n_8394),
.A2(n_7323),
.B1(n_6858),
.B2(n_7186),
.Y(n_9332)
);

AO21x1_ASAP7_75t_L g9333 ( 
.A1(n_8170),
.A2(n_6795),
.B(n_6775),
.Y(n_9333)
);

OR2x2_ASAP7_75t_L g9334 ( 
.A(n_7883),
.B(n_6794),
.Y(n_9334)
);

INVx1_ASAP7_75t_L g9335 ( 
.A(n_7944),
.Y(n_9335)
);

AND2x2_ASAP7_75t_L g9336 ( 
.A(n_8363),
.B(n_7477),
.Y(n_9336)
);

AND2x4_ASAP7_75t_L g9337 ( 
.A(n_7946),
.B(n_7141),
.Y(n_9337)
);

INVx3_ASAP7_75t_L g9338 ( 
.A(n_7873),
.Y(n_9338)
);

INVx2_ASAP7_75t_SL g9339 ( 
.A(n_7967),
.Y(n_9339)
);

INVx2_ASAP7_75t_SL g9340 ( 
.A(n_7967),
.Y(n_9340)
);

INVx2_ASAP7_75t_L g9341 ( 
.A(n_7878),
.Y(n_9341)
);

AND2x2_ASAP7_75t_L g9342 ( 
.A(n_8363),
.B(n_7477),
.Y(n_9342)
);

HB1xp67_ASAP7_75t_L g9343 ( 
.A(n_7997),
.Y(n_9343)
);

NAND2xp5_ASAP7_75t_L g9344 ( 
.A(n_7939),
.B(n_7200),
.Y(n_9344)
);

INVxp67_ASAP7_75t_L g9345 ( 
.A(n_8138),
.Y(n_9345)
);

INVx2_ASAP7_75t_L g9346 ( 
.A(n_7878),
.Y(n_9346)
);

OAI21x1_ASAP7_75t_L g9347 ( 
.A1(n_8498),
.A2(n_7297),
.B(n_6697),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_7944),
.Y(n_9348)
);

INVx1_ASAP7_75t_L g9349 ( 
.A(n_7950),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_7950),
.Y(n_9350)
);

INVx1_ASAP7_75t_L g9351 ( 
.A(n_7959),
.Y(n_9351)
);

BUFx2_ASAP7_75t_L g9352 ( 
.A(n_7798),
.Y(n_9352)
);

AND2x2_ASAP7_75t_L g9353 ( 
.A(n_8383),
.B(n_7485),
.Y(n_9353)
);

BUFx6f_ASAP7_75t_L g9354 ( 
.A(n_7980),
.Y(n_9354)
);

INVx1_ASAP7_75t_L g9355 ( 
.A(n_7959),
.Y(n_9355)
);

NAND2xp5_ASAP7_75t_SL g9356 ( 
.A(n_8246),
.B(n_6785),
.Y(n_9356)
);

INVx3_ASAP7_75t_L g9357 ( 
.A(n_7873),
.Y(n_9357)
);

INVx1_ASAP7_75t_L g9358 ( 
.A(n_7960),
.Y(n_9358)
);

INVx2_ASAP7_75t_L g9359 ( 
.A(n_7889),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_7960),
.Y(n_9360)
);

INVx2_ASAP7_75t_L g9361 ( 
.A(n_7889),
.Y(n_9361)
);

INVx2_ASAP7_75t_SL g9362 ( 
.A(n_7980),
.Y(n_9362)
);

AND2x2_ASAP7_75t_L g9363 ( 
.A(n_8383),
.B(n_7485),
.Y(n_9363)
);

HB1xp67_ASAP7_75t_L g9364 ( 
.A(n_7997),
.Y(n_9364)
);

BUFx2_ASAP7_75t_L g9365 ( 
.A(n_7798),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_7961),
.Y(n_9366)
);

HB1xp67_ASAP7_75t_L g9367 ( 
.A(n_8005),
.Y(n_9367)
);

BUFx6f_ASAP7_75t_L g9368 ( 
.A(n_7980),
.Y(n_9368)
);

BUFx2_ASAP7_75t_L g9369 ( 
.A(n_7798),
.Y(n_9369)
);

INVxp67_ASAP7_75t_L g9370 ( 
.A(n_8679),
.Y(n_9370)
);

OA21x2_ASAP7_75t_L g9371 ( 
.A1(n_7805),
.A2(n_7169),
.B(n_7166),
.Y(n_9371)
);

INVx1_ASAP7_75t_L g9372 ( 
.A(n_7961),
.Y(n_9372)
);

INVx2_ASAP7_75t_L g9373 ( 
.A(n_7889),
.Y(n_9373)
);

INVx2_ASAP7_75t_L g9374 ( 
.A(n_7891),
.Y(n_9374)
);

NAND2xp5_ASAP7_75t_L g9375 ( 
.A(n_7939),
.B(n_7238),
.Y(n_9375)
);

OAI21x1_ASAP7_75t_L g9376 ( 
.A1(n_8112),
.A2(n_7297),
.B(n_6697),
.Y(n_9376)
);

AND2x2_ASAP7_75t_L g9377 ( 
.A(n_8383),
.B(n_7485),
.Y(n_9377)
);

INVx2_ASAP7_75t_L g9378 ( 
.A(n_7891),
.Y(n_9378)
);

INVx1_ASAP7_75t_L g9379 ( 
.A(n_7963),
.Y(n_9379)
);

INVx3_ASAP7_75t_L g9380 ( 
.A(n_7873),
.Y(n_9380)
);

NAND2xp5_ASAP7_75t_L g9381 ( 
.A(n_8137),
.B(n_7238),
.Y(n_9381)
);

OR2x6_ASAP7_75t_L g9382 ( 
.A(n_8145),
.B(n_6932),
.Y(n_9382)
);

AND2x2_ASAP7_75t_L g9383 ( 
.A(n_8399),
.B(n_7485),
.Y(n_9383)
);

INVx2_ASAP7_75t_L g9384 ( 
.A(n_7891),
.Y(n_9384)
);

OAI22xp5_ASAP7_75t_L g9385 ( 
.A1(n_7970),
.A2(n_6947),
.B1(n_7047),
.B2(n_6785),
.Y(n_9385)
);

OAI21x1_ASAP7_75t_L g9386 ( 
.A1(n_8112),
.A2(n_7297),
.B(n_6697),
.Y(n_9386)
);

OAI21x1_ASAP7_75t_SL g9387 ( 
.A1(n_8534),
.A2(n_6795),
.B(n_6775),
.Y(n_9387)
);

INVx2_ASAP7_75t_L g9388 ( 
.A(n_7905),
.Y(n_9388)
);

INVx3_ASAP7_75t_L g9389 ( 
.A(n_7953),
.Y(n_9389)
);

INVx2_ASAP7_75t_L g9390 ( 
.A(n_7905),
.Y(n_9390)
);

INVx1_ASAP7_75t_L g9391 ( 
.A(n_7963),
.Y(n_9391)
);

INVx1_ASAP7_75t_L g9392 ( 
.A(n_7966),
.Y(n_9392)
);

AO21x2_ASAP7_75t_L g9393 ( 
.A1(n_7839),
.A2(n_7475),
.B(n_7047),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_7966),
.Y(n_9394)
);

HB1xp67_ASAP7_75t_L g9395 ( 
.A(n_8005),
.Y(n_9395)
);

BUFx2_ASAP7_75t_L g9396 ( 
.A(n_7798),
.Y(n_9396)
);

AOI21x1_ASAP7_75t_L g9397 ( 
.A1(n_7892),
.A2(n_7761),
.B(n_7740),
.Y(n_9397)
);

INVx3_ASAP7_75t_L g9398 ( 
.A(n_7953),
.Y(n_9398)
);

BUFx6f_ASAP7_75t_SL g9399 ( 
.A(n_8016),
.Y(n_9399)
);

BUFx3_ASAP7_75t_L g9400 ( 
.A(n_8593),
.Y(n_9400)
);

INVx2_ASAP7_75t_L g9401 ( 
.A(n_7905),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_7914),
.Y(n_9402)
);

AO21x2_ASAP7_75t_L g9403 ( 
.A1(n_7903),
.A2(n_7288),
.B(n_6952),
.Y(n_9403)
);

HB1xp67_ASAP7_75t_L g9404 ( 
.A(n_8031),
.Y(n_9404)
);

INVx1_ASAP7_75t_L g9405 ( 
.A(n_7974),
.Y(n_9405)
);

BUFx4f_ASAP7_75t_SL g9406 ( 
.A(n_7952),
.Y(n_9406)
);

INVx1_ASAP7_75t_L g9407 ( 
.A(n_7974),
.Y(n_9407)
);

INVx1_ASAP7_75t_L g9408 ( 
.A(n_7975),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_7914),
.Y(n_9409)
);

BUFx6f_ASAP7_75t_L g9410 ( 
.A(n_8016),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_7975),
.Y(n_9411)
);

INVx2_ASAP7_75t_SL g9412 ( 
.A(n_8016),
.Y(n_9412)
);

HB1xp67_ASAP7_75t_L g9413 ( 
.A(n_8031),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_7984),
.Y(n_9414)
);

INVx2_ASAP7_75t_L g9415 ( 
.A(n_7914),
.Y(n_9415)
);

AND2x2_ASAP7_75t_L g9416 ( 
.A(n_8399),
.B(n_7507),
.Y(n_9416)
);

INVx1_ASAP7_75t_L g9417 ( 
.A(n_7984),
.Y(n_9417)
);

AND2x2_ASAP7_75t_L g9418 ( 
.A(n_8399),
.B(n_7507),
.Y(n_9418)
);

INVx2_ASAP7_75t_L g9419 ( 
.A(n_7922),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_7985),
.Y(n_9420)
);

INVx2_ASAP7_75t_L g9421 ( 
.A(n_7922),
.Y(n_9421)
);

INVx3_ASAP7_75t_L g9422 ( 
.A(n_7953),
.Y(n_9422)
);

AOI22xp5_ASAP7_75t_L g9423 ( 
.A1(n_7865),
.A2(n_6970),
.B1(n_7326),
.B2(n_7328),
.Y(n_9423)
);

OAI21x1_ASAP7_75t_L g9424 ( 
.A1(n_7953),
.A2(n_6723),
.B(n_6681),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_7985),
.Y(n_9425)
);

INVx1_ASAP7_75t_L g9426 ( 
.A(n_7989),
.Y(n_9426)
);

NAND2xp5_ASAP7_75t_L g9427 ( 
.A(n_8137),
.B(n_6833),
.Y(n_9427)
);

INVx2_ASAP7_75t_L g9428 ( 
.A(n_7922),
.Y(n_9428)
);

AO21x2_ASAP7_75t_L g9429 ( 
.A1(n_7903),
.A2(n_7288),
.B(n_6952),
.Y(n_9429)
);

BUFx2_ASAP7_75t_L g9430 ( 
.A(n_8482),
.Y(n_9430)
);

AND2x2_ASAP7_75t_L g9431 ( 
.A(n_8400),
.B(n_8411),
.Y(n_9431)
);

INVx2_ASAP7_75t_L g9432 ( 
.A(n_7924),
.Y(n_9432)
);

NOR2x1_ASAP7_75t_L g9433 ( 
.A(n_8175),
.B(n_6702),
.Y(n_9433)
);

AND2x2_ASAP7_75t_L g9434 ( 
.A(n_8400),
.B(n_7507),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_7989),
.Y(n_9435)
);

AND2x2_ASAP7_75t_L g9436 ( 
.A(n_8400),
.B(n_7507),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_7990),
.Y(n_9437)
);

AND2x2_ASAP7_75t_L g9438 ( 
.A(n_8411),
.B(n_7580),
.Y(n_9438)
);

AND2x2_ASAP7_75t_L g9439 ( 
.A(n_8411),
.B(n_7580),
.Y(n_9439)
);

INVx1_ASAP7_75t_L g9440 ( 
.A(n_7990),
.Y(n_9440)
);

INVx2_ASAP7_75t_L g9441 ( 
.A(n_7924),
.Y(n_9441)
);

INVx1_ASAP7_75t_L g9442 ( 
.A(n_7993),
.Y(n_9442)
);

AND2x2_ASAP7_75t_L g9443 ( 
.A(n_8426),
.B(n_8428),
.Y(n_9443)
);

INVx2_ASAP7_75t_L g9444 ( 
.A(n_7924),
.Y(n_9444)
);

INVx1_ASAP7_75t_L g9445 ( 
.A(n_7993),
.Y(n_9445)
);

INVx3_ASAP7_75t_L g9446 ( 
.A(n_8235),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_7994),
.Y(n_9447)
);

INVx1_ASAP7_75t_L g9448 ( 
.A(n_7994),
.Y(n_9448)
);

OA21x2_ASAP7_75t_L g9449 ( 
.A1(n_7835),
.A2(n_8181),
.B(n_8142),
.Y(n_9449)
);

BUFx6f_ASAP7_75t_L g9450 ( 
.A(n_8048),
.Y(n_9450)
);

INVx1_ASAP7_75t_L g9451 ( 
.A(n_7998),
.Y(n_9451)
);

INVx2_ASAP7_75t_L g9452 ( 
.A(n_7934),
.Y(n_9452)
);

AND2x2_ASAP7_75t_L g9453 ( 
.A(n_8426),
.B(n_7580),
.Y(n_9453)
);

BUFx3_ASAP7_75t_L g9454 ( 
.A(n_8593),
.Y(n_9454)
);

AND2x4_ASAP7_75t_L g9455 ( 
.A(n_8127),
.B(n_7958),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_7998),
.Y(n_9456)
);

BUFx2_ASAP7_75t_L g9457 ( 
.A(n_8482),
.Y(n_9457)
);

INVx1_ASAP7_75t_L g9458 ( 
.A(n_8000),
.Y(n_9458)
);

AOI21xp33_ASAP7_75t_SL g9459 ( 
.A1(n_7817),
.A2(n_7235),
.B(n_6986),
.Y(n_9459)
);

NAND2xp5_ASAP7_75t_L g9460 ( 
.A(n_7970),
.B(n_6196),
.Y(n_9460)
);

OAI21x1_ASAP7_75t_L g9461 ( 
.A1(n_8701),
.A2(n_6723),
.B(n_6681),
.Y(n_9461)
);

OAI21x1_ASAP7_75t_L g9462 ( 
.A1(n_8701),
.A2(n_8742),
.B(n_7892),
.Y(n_9462)
);

CKINVDCx5p33_ASAP7_75t_R g9463 ( 
.A(n_8382),
.Y(n_9463)
);

INVx2_ASAP7_75t_L g9464 ( 
.A(n_7934),
.Y(n_9464)
);

AND2x2_ASAP7_75t_L g9465 ( 
.A(n_8426),
.B(n_7580),
.Y(n_9465)
);

AND2x2_ASAP7_75t_L g9466 ( 
.A(n_8428),
.B(n_7643),
.Y(n_9466)
);

OA21x2_ASAP7_75t_L g9467 ( 
.A1(n_7835),
.A2(n_7169),
.B(n_7166),
.Y(n_9467)
);

OAI21xp5_ASAP7_75t_L g9468 ( 
.A1(n_7996),
.A2(n_6849),
.B(n_6947),
.Y(n_9468)
);

OAI21x1_ASAP7_75t_L g9469 ( 
.A1(n_8701),
.A2(n_6723),
.B(n_6681),
.Y(n_9469)
);

AND2x2_ASAP7_75t_L g9470 ( 
.A(n_8428),
.B(n_7643),
.Y(n_9470)
);

OA21x2_ASAP7_75t_L g9471 ( 
.A1(n_7835),
.A2(n_7182),
.B(n_7178),
.Y(n_9471)
);

INVx5_ASAP7_75t_L g9472 ( 
.A(n_7977),
.Y(n_9472)
);

HB1xp67_ASAP7_75t_L g9473 ( 
.A(n_8764),
.Y(n_9473)
);

BUFx6f_ASAP7_75t_L g9474 ( 
.A(n_8048),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_8000),
.Y(n_9475)
);

AND2x4_ASAP7_75t_L g9476 ( 
.A(n_8127),
.B(n_7141),
.Y(n_9476)
);

INVx3_ASAP7_75t_L g9477 ( 
.A(n_8235),
.Y(n_9477)
);

INVx2_ASAP7_75t_L g9478 ( 
.A(n_7934),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_8003),
.Y(n_9479)
);

INVx2_ASAP7_75t_L g9480 ( 
.A(n_7940),
.Y(n_9480)
);

BUFx2_ASAP7_75t_L g9481 ( 
.A(n_8482),
.Y(n_9481)
);

INVx1_ASAP7_75t_L g9482 ( 
.A(n_8003),
.Y(n_9482)
);

INVx1_ASAP7_75t_L g9483 ( 
.A(n_8006),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_8006),
.Y(n_9484)
);

OAI21x1_ASAP7_75t_L g9485 ( 
.A1(n_8742),
.A2(n_6723),
.B(n_6681),
.Y(n_9485)
);

AND2x2_ASAP7_75t_L g9486 ( 
.A(n_8437),
.B(n_7643),
.Y(n_9486)
);

OR2x2_ASAP7_75t_L g9487 ( 
.A(n_8315),
.B(n_7503),
.Y(n_9487)
);

INVx1_ASAP7_75t_L g9488 ( 
.A(n_8009),
.Y(n_9488)
);

INVx1_ASAP7_75t_L g9489 ( 
.A(n_8009),
.Y(n_9489)
);

AND2x2_ASAP7_75t_L g9490 ( 
.A(n_8437),
.B(n_7643),
.Y(n_9490)
);

INVx2_ASAP7_75t_L g9491 ( 
.A(n_7940),
.Y(n_9491)
);

INVx3_ASAP7_75t_L g9492 ( 
.A(n_8235),
.Y(n_9492)
);

HB1xp67_ASAP7_75t_L g9493 ( 
.A(n_8764),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_8010),
.Y(n_9494)
);

INVx2_ASAP7_75t_L g9495 ( 
.A(n_7940),
.Y(n_9495)
);

NAND2xp5_ASAP7_75t_L g9496 ( 
.A(n_8493),
.B(n_6196),
.Y(n_9496)
);

INVx1_ASAP7_75t_L g9497 ( 
.A(n_8010),
.Y(n_9497)
);

INVx2_ASAP7_75t_L g9498 ( 
.A(n_7942),
.Y(n_9498)
);

OA21x2_ASAP7_75t_L g9499 ( 
.A1(n_8181),
.A2(n_7182),
.B(n_7178),
.Y(n_9499)
);

AND2x2_ASAP7_75t_L g9500 ( 
.A(n_8437),
.B(n_7651),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_7942),
.Y(n_9501)
);

OA21x2_ASAP7_75t_L g9502 ( 
.A1(n_8142),
.A2(n_7182),
.B(n_7178),
.Y(n_9502)
);

AOI22xp33_ASAP7_75t_L g9503 ( 
.A1(n_8394),
.A2(n_7323),
.B1(n_6876),
.B2(n_6967),
.Y(n_9503)
);

HB1xp67_ASAP7_75t_L g9504 ( 
.A(n_8755),
.Y(n_9504)
);

INVx1_ASAP7_75t_L g9505 ( 
.A(n_8013),
.Y(n_9505)
);

INVx2_ASAP7_75t_L g9506 ( 
.A(n_7942),
.Y(n_9506)
);

INVx3_ASAP7_75t_L g9507 ( 
.A(n_8235),
.Y(n_9507)
);

INVx1_ASAP7_75t_L g9508 ( 
.A(n_8013),
.Y(n_9508)
);

AOI22xp33_ASAP7_75t_SL g9509 ( 
.A1(n_8534),
.A2(n_7124),
.B1(n_6956),
.B2(n_6785),
.Y(n_9509)
);

NOR2xp67_ASAP7_75t_R g9510 ( 
.A(n_7977),
.B(n_6749),
.Y(n_9510)
);

INVx2_ASAP7_75t_L g9511 ( 
.A(n_7947),
.Y(n_9511)
);

NAND2xp5_ASAP7_75t_L g9512 ( 
.A(n_8493),
.B(n_6201),
.Y(n_9512)
);

INVx2_ASAP7_75t_L g9513 ( 
.A(n_7947),
.Y(n_9513)
);

INVx1_ASAP7_75t_L g9514 ( 
.A(n_8014),
.Y(n_9514)
);

INVx1_ASAP7_75t_L g9515 ( 
.A(n_8014),
.Y(n_9515)
);

OAI21x1_ASAP7_75t_L g9516 ( 
.A1(n_8742),
.A2(n_6797),
.B(n_6737),
.Y(n_9516)
);

OAI21xp5_ASAP7_75t_L g9517 ( 
.A1(n_8139),
.A2(n_6937),
.B(n_6909),
.Y(n_9517)
);

INVx2_ASAP7_75t_L g9518 ( 
.A(n_7947),
.Y(n_9518)
);

BUFx3_ASAP7_75t_L g9519 ( 
.A(n_8617),
.Y(n_9519)
);

INVx2_ASAP7_75t_L g9520 ( 
.A(n_7956),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8019),
.Y(n_9521)
);

INVx1_ASAP7_75t_L g9522 ( 
.A(n_8019),
.Y(n_9522)
);

INVx3_ASAP7_75t_L g9523 ( 
.A(n_8353),
.Y(n_9523)
);

INVx2_ASAP7_75t_L g9524 ( 
.A(n_7956),
.Y(n_9524)
);

INVx2_ASAP7_75t_SL g9525 ( 
.A(n_8048),
.Y(n_9525)
);

INVx1_ASAP7_75t_SL g9526 ( 
.A(n_8617),
.Y(n_9526)
);

AND2x2_ASAP7_75t_L g9527 ( 
.A(n_8502),
.B(n_8510),
.Y(n_9527)
);

NAND2xp5_ASAP7_75t_L g9528 ( 
.A(n_8547),
.B(n_6201),
.Y(n_9528)
);

BUFx12f_ASAP7_75t_L g9529 ( 
.A(n_8640),
.Y(n_9529)
);

INVx2_ASAP7_75t_L g9530 ( 
.A(n_7956),
.Y(n_9530)
);

INVx2_ASAP7_75t_L g9531 ( 
.A(n_7957),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_8024),
.Y(n_9532)
);

INVx3_ASAP7_75t_L g9533 ( 
.A(n_8353),
.Y(n_9533)
);

CKINVDCx5p33_ASAP7_75t_R g9534 ( 
.A(n_8382),
.Y(n_9534)
);

INVx2_ASAP7_75t_L g9535 ( 
.A(n_7957),
.Y(n_9535)
);

INVx2_ASAP7_75t_L g9536 ( 
.A(n_7957),
.Y(n_9536)
);

AND2x2_ASAP7_75t_L g9537 ( 
.A(n_8502),
.B(n_8510),
.Y(n_9537)
);

INVx1_ASAP7_75t_L g9538 ( 
.A(n_8024),
.Y(n_9538)
);

OR2x2_ASAP7_75t_L g9539 ( 
.A(n_8315),
.B(n_7544),
.Y(n_9539)
);

INVx2_ASAP7_75t_L g9540 ( 
.A(n_7981),
.Y(n_9540)
);

AO21x2_ASAP7_75t_L g9541 ( 
.A1(n_7903),
.A2(n_8343),
.B(n_8480),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_8032),
.Y(n_9542)
);

AO31x2_ASAP7_75t_L g9543 ( 
.A1(n_8560),
.A2(n_7516),
.A3(n_6761),
.B(n_7345),
.Y(n_9543)
);

INVx2_ASAP7_75t_L g9544 ( 
.A(n_7981),
.Y(n_9544)
);

HB1xp67_ASAP7_75t_L g9545 ( 
.A(n_8755),
.Y(n_9545)
);

INVx2_ASAP7_75t_SL g9546 ( 
.A(n_8110),
.Y(n_9546)
);

AOI22xp33_ASAP7_75t_L g9547 ( 
.A1(n_8349),
.A2(n_6905),
.B1(n_7407),
.B2(n_6802),
.Y(n_9547)
);

INVx2_ASAP7_75t_L g9548 ( 
.A(n_7981),
.Y(n_9548)
);

INVx1_ASAP7_75t_L g9549 ( 
.A(n_8032),
.Y(n_9549)
);

OR2x2_ASAP7_75t_L g9550 ( 
.A(n_8404),
.B(n_7544),
.Y(n_9550)
);

INVx1_ASAP7_75t_L g9551 ( 
.A(n_8034),
.Y(n_9551)
);

INVx2_ASAP7_75t_L g9552 ( 
.A(n_7983),
.Y(n_9552)
);

BUFx2_ASAP7_75t_L g9553 ( 
.A(n_8482),
.Y(n_9553)
);

BUFx2_ASAP7_75t_SL g9554 ( 
.A(n_7927),
.Y(n_9554)
);

INVx1_ASAP7_75t_L g9555 ( 
.A(n_8034),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_8035),
.Y(n_9556)
);

BUFx3_ASAP7_75t_L g9557 ( 
.A(n_8640),
.Y(n_9557)
);

INVx1_ASAP7_75t_L g9558 ( 
.A(n_8035),
.Y(n_9558)
);

OAI21x1_ASAP7_75t_L g9559 ( 
.A1(n_7892),
.A2(n_6797),
.B(n_6737),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_8037),
.Y(n_9560)
);

HB1xp67_ASAP7_75t_L g9561 ( 
.A(n_8748),
.Y(n_9561)
);

AND2x2_ASAP7_75t_L g9562 ( 
.A(n_8502),
.B(n_8510),
.Y(n_9562)
);

OR2x2_ASAP7_75t_L g9563 ( 
.A(n_8404),
.B(n_7887),
.Y(n_9563)
);

OR2x6_ASAP7_75t_L g9564 ( 
.A(n_8175),
.B(n_6932),
.Y(n_9564)
);

INVx2_ASAP7_75t_L g9565 ( 
.A(n_7983),
.Y(n_9565)
);

INVx2_ASAP7_75t_L g9566 ( 
.A(n_7983),
.Y(n_9566)
);

OA21x2_ASAP7_75t_L g9567 ( 
.A1(n_7911),
.A2(n_7212),
.B(n_7198),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_8037),
.Y(n_9568)
);

INVx3_ASAP7_75t_L g9569 ( 
.A(n_8353),
.Y(n_9569)
);

INVx2_ASAP7_75t_L g9570 ( 
.A(n_7999),
.Y(n_9570)
);

BUFx2_ASAP7_75t_L g9571 ( 
.A(n_8482),
.Y(n_9571)
);

INVx1_ASAP7_75t_L g9572 ( 
.A(n_8047),
.Y(n_9572)
);

OAI21x1_ASAP7_75t_L g9573 ( 
.A1(n_8353),
.A2(n_6797),
.B(n_6737),
.Y(n_9573)
);

OAI21x1_ASAP7_75t_L g9574 ( 
.A1(n_8419),
.A2(n_8604),
.B(n_8420),
.Y(n_9574)
);

INVx2_ASAP7_75t_L g9575 ( 
.A(n_7999),
.Y(n_9575)
);

INVx1_ASAP7_75t_L g9576 ( 
.A(n_8047),
.Y(n_9576)
);

INVx1_ASAP7_75t_L g9577 ( 
.A(n_8052),
.Y(n_9577)
);

INVxp67_ASAP7_75t_SL g9578 ( 
.A(n_7920),
.Y(n_9578)
);

NAND2xp5_ASAP7_75t_L g9579 ( 
.A(n_8547),
.B(n_6775),
.Y(n_9579)
);

INVx2_ASAP7_75t_L g9580 ( 
.A(n_7999),
.Y(n_9580)
);

INVx1_ASAP7_75t_L g9581 ( 
.A(n_8052),
.Y(n_9581)
);

AND2x2_ASAP7_75t_L g9582 ( 
.A(n_7958),
.B(n_7651),
.Y(n_9582)
);

OR2x2_ASAP7_75t_L g9583 ( 
.A(n_7887),
.B(n_7583),
.Y(n_9583)
);

HB1xp67_ASAP7_75t_L g9584 ( 
.A(n_8748),
.Y(n_9584)
);

INVx2_ASAP7_75t_SL g9585 ( 
.A(n_8110),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_8054),
.Y(n_9586)
);

INVx3_ASAP7_75t_L g9587 ( 
.A(n_8419),
.Y(n_9587)
);

BUFx2_ASAP7_75t_L g9588 ( 
.A(n_8127),
.Y(n_9588)
);

OAI21x1_ASAP7_75t_L g9589 ( 
.A1(n_8419),
.A2(n_6797),
.B(n_6737),
.Y(n_9589)
);

NAND2xp5_ASAP7_75t_L g9590 ( 
.A(n_8028),
.B(n_6775),
.Y(n_9590)
);

AO21x2_ASAP7_75t_L g9591 ( 
.A1(n_7903),
.A2(n_7269),
.B(n_7236),
.Y(n_9591)
);

AND2x2_ASAP7_75t_L g9592 ( 
.A(n_7958),
.B(n_7976),
.Y(n_9592)
);

AOI22xp33_ASAP7_75t_L g9593 ( 
.A1(n_8349),
.A2(n_6905),
.B1(n_7407),
.B2(n_6855),
.Y(n_9593)
);

OAI21x1_ASAP7_75t_L g9594 ( 
.A1(n_8419),
.A2(n_6951),
.B(n_6808),
.Y(n_9594)
);

INVx2_ASAP7_75t_L g9595 ( 
.A(n_8002),
.Y(n_9595)
);

NAND2xp5_ASAP7_75t_L g9596 ( 
.A(n_8028),
.B(n_6795),
.Y(n_9596)
);

INVx1_ASAP7_75t_L g9597 ( 
.A(n_8054),
.Y(n_9597)
);

INVx1_ASAP7_75t_L g9598 ( 
.A(n_8056),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_8002),
.Y(n_9599)
);

INVx2_ASAP7_75t_L g9600 ( 
.A(n_8002),
.Y(n_9600)
);

AO21x2_ASAP7_75t_L g9601 ( 
.A1(n_7903),
.A2(n_7269),
.B(n_7236),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_8008),
.Y(n_9602)
);

AO21x2_ASAP7_75t_L g9603 ( 
.A1(n_8343),
.A2(n_6917),
.B(n_6843),
.Y(n_9603)
);

HB1xp67_ASAP7_75t_L g9604 ( 
.A(n_8725),
.Y(n_9604)
);

OR2x2_ASAP7_75t_L g9605 ( 
.A(n_7887),
.B(n_7583),
.Y(n_9605)
);

INVx1_ASAP7_75t_L g9606 ( 
.A(n_8056),
.Y(n_9606)
);

INVx2_ASAP7_75t_L g9607 ( 
.A(n_8008),
.Y(n_9607)
);

INVx1_ASAP7_75t_L g9608 ( 
.A(n_8061),
.Y(n_9608)
);

CKINVDCx20_ASAP7_75t_R g9609 ( 
.A(n_8406),
.Y(n_9609)
);

BUFx3_ASAP7_75t_L g9610 ( 
.A(n_8812),
.Y(n_9610)
);

INVxp67_ASAP7_75t_SL g9611 ( 
.A(n_8519),
.Y(n_9611)
);

BUFx3_ASAP7_75t_L g9612 ( 
.A(n_8812),
.Y(n_9612)
);

AOI21xp33_ASAP7_75t_L g9613 ( 
.A1(n_8139),
.A2(n_8797),
.B(n_8462),
.Y(n_9613)
);

INVx1_ASAP7_75t_L g9614 ( 
.A(n_8061),
.Y(n_9614)
);

AND2x2_ASAP7_75t_L g9615 ( 
.A(n_7958),
.B(n_7651),
.Y(n_9615)
);

INVx1_ASAP7_75t_L g9616 ( 
.A(n_8062),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_7958),
.B(n_7651),
.Y(n_9617)
);

AO21x2_ASAP7_75t_L g9618 ( 
.A1(n_8480),
.A2(n_6917),
.B(n_6843),
.Y(n_9618)
);

INVx2_ASAP7_75t_L g9619 ( 
.A(n_8008),
.Y(n_9619)
);

INVx2_ASAP7_75t_L g9620 ( 
.A(n_8011),
.Y(n_9620)
);

OA21x2_ASAP7_75t_L g9621 ( 
.A1(n_7911),
.A2(n_7212),
.B(n_7198),
.Y(n_9621)
);

OR2x2_ASAP7_75t_L g9622 ( 
.A(n_8255),
.B(n_6634),
.Y(n_9622)
);

INVx1_ASAP7_75t_L g9623 ( 
.A(n_8062),
.Y(n_9623)
);

OA21x2_ASAP7_75t_L g9624 ( 
.A1(n_8293),
.A2(n_7212),
.B(n_7198),
.Y(n_9624)
);

INVx1_ASAP7_75t_L g9625 ( 
.A(n_8064),
.Y(n_9625)
);

NAND2xp5_ASAP7_75t_L g9626 ( 
.A(n_8557),
.B(n_6795),
.Y(n_9626)
);

BUFx2_ASAP7_75t_L g9627 ( 
.A(n_8127),
.Y(n_9627)
);

INVx4_ASAP7_75t_L g9628 ( 
.A(n_7909),
.Y(n_9628)
);

INVx5_ASAP7_75t_L g9629 ( 
.A(n_7977),
.Y(n_9629)
);

AND2x2_ASAP7_75t_L g9630 ( 
.A(n_7976),
.B(n_7666),
.Y(n_9630)
);

AND2x2_ASAP7_75t_L g9631 ( 
.A(n_7976),
.B(n_7666),
.Y(n_9631)
);

BUFx6f_ASAP7_75t_L g9632 ( 
.A(n_8110),
.Y(n_9632)
);

NAND2xp5_ASAP7_75t_L g9633 ( 
.A(n_8557),
.B(n_8584),
.Y(n_9633)
);

INVx1_ASAP7_75t_L g9634 ( 
.A(n_8064),
.Y(n_9634)
);

INVx2_ASAP7_75t_L g9635 ( 
.A(n_8011),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_8065),
.Y(n_9636)
);

AND2x2_ASAP7_75t_L g9637 ( 
.A(n_7976),
.B(n_7666),
.Y(n_9637)
);

INVx2_ASAP7_75t_L g9638 ( 
.A(n_8011),
.Y(n_9638)
);

OAI21xp5_ASAP7_75t_L g9639 ( 
.A1(n_8408),
.A2(n_6909),
.B(n_6941),
.Y(n_9639)
);

INVx3_ASAP7_75t_L g9640 ( 
.A(n_8420),
.Y(n_9640)
);

INVx2_ASAP7_75t_L g9641 ( 
.A(n_8018),
.Y(n_9641)
);

NOR2xp33_ASAP7_75t_L g9642 ( 
.A(n_8648),
.B(n_7017),
.Y(n_9642)
);

INVx2_ASAP7_75t_L g9643 ( 
.A(n_8018),
.Y(n_9643)
);

INVx2_ASAP7_75t_L g9644 ( 
.A(n_8018),
.Y(n_9644)
);

AND2x2_ASAP7_75t_L g9645 ( 
.A(n_7976),
.B(n_7666),
.Y(n_9645)
);

AOI21x1_ASAP7_75t_L g9646 ( 
.A1(n_8580),
.A2(n_7761),
.B(n_7740),
.Y(n_9646)
);

INVx1_ASAP7_75t_L g9647 ( 
.A(n_8065),
.Y(n_9647)
);

HB1xp67_ASAP7_75t_L g9648 ( 
.A(n_8725),
.Y(n_9648)
);

INVx1_ASAP7_75t_L g9649 ( 
.A(n_8067),
.Y(n_9649)
);

AO21x2_ASAP7_75t_L g9650 ( 
.A1(n_8580),
.A2(n_7290),
.B(n_7291),
.Y(n_9650)
);

NAND2xp5_ASAP7_75t_L g9651 ( 
.A(n_8584),
.B(n_6857),
.Y(n_9651)
);

OA21x2_ASAP7_75t_L g9652 ( 
.A1(n_8293),
.A2(n_7218),
.B(n_7216),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_8023),
.Y(n_9653)
);

INVx2_ASAP7_75t_L g9654 ( 
.A(n_8023),
.Y(n_9654)
);

AND2x2_ASAP7_75t_L g9655 ( 
.A(n_8051),
.B(n_7719),
.Y(n_9655)
);

HB1xp67_ASAP7_75t_L g9656 ( 
.A(n_8788),
.Y(n_9656)
);

INVx2_ASAP7_75t_SL g9657 ( 
.A(n_8147),
.Y(n_9657)
);

INVx2_ASAP7_75t_SL g9658 ( 
.A(n_8147),
.Y(n_9658)
);

INVx2_ASAP7_75t_L g9659 ( 
.A(n_8023),
.Y(n_9659)
);

AND2x2_ASAP7_75t_L g9660 ( 
.A(n_8051),
.B(n_7719),
.Y(n_9660)
);

AND2x4_ASAP7_75t_SL g9661 ( 
.A(n_8806),
.B(n_7150),
.Y(n_9661)
);

AND2x2_ASAP7_75t_L g9662 ( 
.A(n_8051),
.B(n_7719),
.Y(n_9662)
);

BUFx2_ASAP7_75t_L g9663 ( 
.A(n_8127),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_8067),
.Y(n_9664)
);

INVx3_ASAP7_75t_L g9665 ( 
.A(n_8420),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8068),
.Y(n_9666)
);

INVx2_ASAP7_75t_L g9667 ( 
.A(n_8026),
.Y(n_9667)
);

AND2x2_ASAP7_75t_L g9668 ( 
.A(n_8051),
.B(n_7719),
.Y(n_9668)
);

INVx2_ASAP7_75t_SL g9669 ( 
.A(n_8147),
.Y(n_9669)
);

INVx2_ASAP7_75t_L g9670 ( 
.A(n_8026),
.Y(n_9670)
);

HB1xp67_ASAP7_75t_L g9671 ( 
.A(n_8788),
.Y(n_9671)
);

BUFx2_ASAP7_75t_L g9672 ( 
.A(n_8127),
.Y(n_9672)
);

AO21x2_ASAP7_75t_L g9673 ( 
.A1(n_8580),
.A2(n_7290),
.B(n_7291),
.Y(n_9673)
);

OA21x2_ASAP7_75t_L g9674 ( 
.A1(n_8295),
.A2(n_7218),
.B(n_7216),
.Y(n_9674)
);

INVx2_ASAP7_75t_L g9675 ( 
.A(n_8026),
.Y(n_9675)
);

INVx8_ASAP7_75t_L g9676 ( 
.A(n_8409),
.Y(n_9676)
);

AND2x2_ASAP7_75t_L g9677 ( 
.A(n_8051),
.B(n_6722),
.Y(n_9677)
);

BUFx2_ASAP7_75t_SL g9678 ( 
.A(n_7927),
.Y(n_9678)
);

INVx2_ASAP7_75t_L g9679 ( 
.A(n_8029),
.Y(n_9679)
);

OA21x2_ASAP7_75t_L g9680 ( 
.A1(n_8295),
.A2(n_7218),
.B(n_7216),
.Y(n_9680)
);

NAND2xp5_ASAP7_75t_L g9681 ( 
.A(n_8455),
.B(n_6857),
.Y(n_9681)
);

AND2x4_ASAP7_75t_L g9682 ( 
.A(n_8346),
.B(n_7141),
.Y(n_9682)
);

OAI21xp5_ASAP7_75t_L g9683 ( 
.A1(n_8408),
.A2(n_6879),
.B(n_7205),
.Y(n_9683)
);

AND2x2_ASAP7_75t_L g9684 ( 
.A(n_8346),
.B(n_6722),
.Y(n_9684)
);

OA21x2_ASAP7_75t_L g9685 ( 
.A1(n_7827),
.A2(n_7232),
.B(n_7224),
.Y(n_9685)
);

INVx1_ASAP7_75t_L g9686 ( 
.A(n_8068),
.Y(n_9686)
);

INVx1_ASAP7_75t_L g9687 ( 
.A(n_8071),
.Y(n_9687)
);

NOR2xp33_ASAP7_75t_L g9688 ( 
.A(n_8427),
.B(n_7017),
.Y(n_9688)
);

INVx1_ASAP7_75t_L g9689 ( 
.A(n_8071),
.Y(n_9689)
);

HB1xp67_ASAP7_75t_L g9690 ( 
.A(n_7978),
.Y(n_9690)
);

INVx1_ASAP7_75t_L g9691 ( 
.A(n_8073),
.Y(n_9691)
);

OR2x2_ASAP7_75t_L g9692 ( 
.A(n_8255),
.B(n_6634),
.Y(n_9692)
);

OAI21x1_ASAP7_75t_L g9693 ( 
.A1(n_8420),
.A2(n_6951),
.B(n_6808),
.Y(n_9693)
);

INVx1_ASAP7_75t_L g9694 ( 
.A(n_8073),
.Y(n_9694)
);

INVx2_ASAP7_75t_L g9695 ( 
.A(n_8029),
.Y(n_9695)
);

INVx2_ASAP7_75t_L g9696 ( 
.A(n_9139),
.Y(n_9696)
);

AND2x4_ASAP7_75t_L g9697 ( 
.A(n_9433),
.B(n_7816),
.Y(n_9697)
);

OAI21xp5_ASAP7_75t_L g9698 ( 
.A1(n_8913),
.A2(n_7811),
.B(n_8697),
.Y(n_9698)
);

INVx1_ASAP7_75t_L g9699 ( 
.A(n_8817),
.Y(n_9699)
);

INVx1_ASAP7_75t_L g9700 ( 
.A(n_8992),
.Y(n_9700)
);

NOR2xp33_ASAP7_75t_L g9701 ( 
.A(n_9071),
.B(n_8151),
.Y(n_9701)
);

INVx1_ASAP7_75t_L g9702 ( 
.A(n_8996),
.Y(n_9702)
);

INVxp67_ASAP7_75t_SL g9703 ( 
.A(n_8821),
.Y(n_9703)
);

AND2x2_ASAP7_75t_L g9704 ( 
.A(n_8859),
.B(n_7817),
.Y(n_9704)
);

AOI21xp5_ASAP7_75t_SL g9705 ( 
.A1(n_8851),
.A2(n_8559),
.B(n_7927),
.Y(n_9705)
);

INVx2_ASAP7_75t_L g9706 ( 
.A(n_9139),
.Y(n_9706)
);

AOI22xp33_ASAP7_75t_L g9707 ( 
.A1(n_9035),
.A2(n_9613),
.B1(n_8891),
.B2(n_9101),
.Y(n_9707)
);

AOI21xp5_ASAP7_75t_L g9708 ( 
.A1(n_9273),
.A2(n_8697),
.B(n_8012),
.Y(n_9708)
);

NAND2xp5_ASAP7_75t_L g9709 ( 
.A(n_8859),
.B(n_8166),
.Y(n_9709)
);

AND2x4_ASAP7_75t_L g9710 ( 
.A(n_8821),
.B(n_7816),
.Y(n_9710)
);

AOI221xp5_ASAP7_75t_L g9711 ( 
.A1(n_9229),
.A2(n_8226),
.B1(n_7811),
.B2(n_7875),
.C(n_7890),
.Y(n_9711)
);

AOI22xp5_ASAP7_75t_L g9712 ( 
.A1(n_9274),
.A2(n_8171),
.B1(n_8190),
.B2(n_8560),
.Y(n_9712)
);

A2O1A1Ixp33_ASAP7_75t_L g9713 ( 
.A1(n_9177),
.A2(n_8457),
.B(n_8229),
.C(n_8190),
.Y(n_9713)
);

NAND2xp5_ASAP7_75t_L g9714 ( 
.A(n_8831),
.B(n_8166),
.Y(n_9714)
);

AND2x4_ASAP7_75t_SL g9715 ( 
.A(n_8881),
.B(n_6677),
.Y(n_9715)
);

O2A1O1Ixp33_ASAP7_75t_L g9716 ( 
.A1(n_9270),
.A2(n_8226),
.B(n_8808),
.C(n_8193),
.Y(n_9716)
);

AND2x4_ASAP7_75t_L g9717 ( 
.A(n_8893),
.B(n_7816),
.Y(n_9717)
);

AND2x2_ASAP7_75t_L g9718 ( 
.A(n_8893),
.B(n_7817),
.Y(n_9718)
);

OR2x2_ASAP7_75t_L g9719 ( 
.A(n_9087),
.B(n_8255),
.Y(n_9719)
);

AND2x2_ASAP7_75t_L g9720 ( 
.A(n_8860),
.B(n_7817),
.Y(n_9720)
);

INVx3_ASAP7_75t_L g9721 ( 
.A(n_8861),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_8817),
.Y(n_9722)
);

INVxp67_ASAP7_75t_L g9723 ( 
.A(n_9226),
.Y(n_9723)
);

INVx1_ASAP7_75t_L g9724 ( 
.A(n_8822),
.Y(n_9724)
);

AND2x2_ASAP7_75t_L g9725 ( 
.A(n_8860),
.B(n_8377),
.Y(n_9725)
);

NAND2xp5_ASAP7_75t_L g9726 ( 
.A(n_9207),
.B(n_8193),
.Y(n_9726)
);

AND2x4_ASAP7_75t_L g9727 ( 
.A(n_9030),
.B(n_7816),
.Y(n_9727)
);

OA21x2_ASAP7_75t_L g9728 ( 
.A1(n_9578),
.A2(n_7844),
.B(n_7827),
.Y(n_9728)
);

AOI21x1_ASAP7_75t_L g9729 ( 
.A1(n_9226),
.A2(n_8566),
.B(n_8558),
.Y(n_9729)
);

AOI221xp5_ASAP7_75t_L g9730 ( 
.A1(n_9683),
.A2(n_7875),
.B1(n_7890),
.B2(n_8808),
.C(n_8055),
.Y(n_9730)
);

AND2x2_ASAP7_75t_L g9731 ( 
.A(n_9030),
.B(n_8377),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_8822),
.Y(n_9732)
);

AND2x2_ASAP7_75t_L g9733 ( 
.A(n_9214),
.B(n_8377),
.Y(n_9733)
);

OAI21xp5_ASAP7_75t_L g9734 ( 
.A1(n_9423),
.A2(n_8229),
.B(n_7844),
.Y(n_9734)
);

AND2x2_ASAP7_75t_SL g9735 ( 
.A(n_9218),
.B(n_7801),
.Y(n_9735)
);

AND2x4_ASAP7_75t_L g9736 ( 
.A(n_8920),
.B(n_7816),
.Y(n_9736)
);

AND2x6_ASAP7_75t_L g9737 ( 
.A(n_8814),
.B(n_8830),
.Y(n_9737)
);

OAI21xp5_ASAP7_75t_L g9738 ( 
.A1(n_9273),
.A2(n_7885),
.B(n_8015),
.Y(n_9738)
);

NAND4xp25_ASAP7_75t_L g9739 ( 
.A(n_9214),
.B(n_8888),
.C(n_8952),
.D(n_9070),
.Y(n_9739)
);

AND2x2_ASAP7_75t_L g9740 ( 
.A(n_8918),
.B(n_8377),
.Y(n_9740)
);

OAI21xp5_ASAP7_75t_L g9741 ( 
.A1(n_9153),
.A2(n_7885),
.B(n_8015),
.Y(n_9741)
);

AOI21xp5_ASAP7_75t_L g9742 ( 
.A1(n_9153),
.A2(n_8012),
.B(n_7801),
.Y(n_9742)
);

OAI21xp5_ASAP7_75t_L g9743 ( 
.A1(n_9385),
.A2(n_8729),
.B(n_8330),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9000),
.Y(n_9744)
);

NOR2xp33_ASAP7_75t_L g9745 ( 
.A(n_9286),
.B(n_8151),
.Y(n_9745)
);

AND2x2_ASAP7_75t_L g9746 ( 
.A(n_8918),
.B(n_8519),
.Y(n_9746)
);

NOR2xp33_ASAP7_75t_L g9747 ( 
.A(n_9196),
.B(n_8151),
.Y(n_9747)
);

OR2x2_ASAP7_75t_L g9748 ( 
.A(n_9345),
.B(n_8275),
.Y(n_9748)
);

OR2x2_ASAP7_75t_L g9749 ( 
.A(n_9117),
.B(n_8275),
.Y(n_9749)
);

INVx1_ASAP7_75t_SL g9750 ( 
.A(n_9018),
.Y(n_9750)
);

AND2x2_ASAP7_75t_L g9751 ( 
.A(n_8921),
.B(n_8714),
.Y(n_9751)
);

OR2x6_ASAP7_75t_L g9752 ( 
.A(n_8833),
.B(n_7977),
.Y(n_9752)
);

AND2x2_ASAP7_75t_L g9753 ( 
.A(n_8921),
.B(n_8714),
.Y(n_9753)
);

A2O1A1Ixp33_ASAP7_75t_L g9754 ( 
.A1(n_9468),
.A2(n_8457),
.B(n_8055),
.C(n_8238),
.Y(n_9754)
);

AND2x4_ASAP7_75t_L g9755 ( 
.A(n_8920),
.B(n_7886),
.Y(n_9755)
);

AO21x2_ASAP7_75t_L g9756 ( 
.A1(n_9089),
.A2(n_8330),
.B(n_8468),
.Y(n_9756)
);

AND2x4_ASAP7_75t_L g9757 ( 
.A(n_8924),
.B(n_7886),
.Y(n_9757)
);

CKINVDCx6p67_ASAP7_75t_R g9758 ( 
.A(n_9311),
.Y(n_9758)
);

AND2x2_ASAP7_75t_L g9759 ( 
.A(n_9592),
.B(n_8621),
.Y(n_9759)
);

BUFx3_ASAP7_75t_L g9760 ( 
.A(n_8962),
.Y(n_9760)
);

OR2x2_ASAP7_75t_L g9761 ( 
.A(n_8941),
.B(n_8275),
.Y(n_9761)
);

A2O1A1Ixp33_ASAP7_75t_L g9762 ( 
.A1(n_9639),
.A2(n_8238),
.B(n_7857),
.C(n_7968),
.Y(n_9762)
);

AND2x4_ASAP7_75t_L g9763 ( 
.A(n_8924),
.B(n_7886),
.Y(n_9763)
);

NAND3xp33_ASAP7_75t_L g9764 ( 
.A(n_8929),
.B(n_8288),
.C(n_8797),
.Y(n_9764)
);

OA21x2_ASAP7_75t_L g9765 ( 
.A1(n_9154),
.A2(n_9168),
.B(n_9559),
.Y(n_9765)
);

O2A1O1Ixp33_ASAP7_75t_SL g9766 ( 
.A1(n_9370),
.A2(n_8746),
.B(n_7231),
.C(n_7242),
.Y(n_9766)
);

AND2x2_ASAP7_75t_L g9767 ( 
.A(n_9592),
.B(n_8621),
.Y(n_9767)
);

NOR2x1p5_ASAP7_75t_L g9768 ( 
.A(n_8962),
.B(n_8749),
.Y(n_9768)
);

AND2x2_ASAP7_75t_L g9769 ( 
.A(n_8833),
.B(n_8883),
.Y(n_9769)
);

BUFx6f_ASAP7_75t_L g9770 ( 
.A(n_8900),
.Y(n_9770)
);

AND2x2_ASAP7_75t_L g9771 ( 
.A(n_8883),
.B(n_8178),
.Y(n_9771)
);

INVx2_ASAP7_75t_L g9772 ( 
.A(n_9139),
.Y(n_9772)
);

AND2x4_ASAP7_75t_L g9773 ( 
.A(n_8928),
.B(n_8957),
.Y(n_9773)
);

NAND2xp5_ASAP7_75t_L g9774 ( 
.A(n_8928),
.B(n_8957),
.Y(n_9774)
);

NOR2xp33_ASAP7_75t_L g9775 ( 
.A(n_9196),
.B(n_8749),
.Y(n_9775)
);

AO32x2_ASAP7_75t_L g9776 ( 
.A1(n_8873),
.A2(n_7929),
.A3(n_8488),
.B1(n_8610),
.B2(n_8616),
.Y(n_9776)
);

HB1xp67_ASAP7_75t_L g9777 ( 
.A(n_8816),
.Y(n_9777)
);

AND2x4_ASAP7_75t_L g9778 ( 
.A(n_8991),
.B(n_7886),
.Y(n_9778)
);

INVxp67_ASAP7_75t_L g9779 ( 
.A(n_8940),
.Y(n_9779)
);

AND2x2_ASAP7_75t_L g9780 ( 
.A(n_8940),
.B(n_8178),
.Y(n_9780)
);

INVx1_ASAP7_75t_L g9781 ( 
.A(n_9012),
.Y(n_9781)
);

OR2x2_ASAP7_75t_L g9782 ( 
.A(n_8943),
.B(n_8344),
.Y(n_9782)
);

NOR2xp33_ASAP7_75t_L g9783 ( 
.A(n_9216),
.B(n_8749),
.Y(n_9783)
);

HB1xp67_ASAP7_75t_L g9784 ( 
.A(n_8824),
.Y(n_9784)
);

NOR2x1_ASAP7_75t_SL g9785 ( 
.A(n_8818),
.B(n_8815),
.Y(n_9785)
);

OA21x2_ASAP7_75t_L g9786 ( 
.A1(n_9559),
.A2(n_8053),
.B(n_8029),
.Y(n_9786)
);

AND2x4_ASAP7_75t_L g9787 ( 
.A(n_8991),
.B(n_7886),
.Y(n_9787)
);

NOR2xp33_ASAP7_75t_L g9788 ( 
.A(n_9216),
.B(n_8157),
.Y(n_9788)
);

AND2x2_ASAP7_75t_L g9789 ( 
.A(n_8825),
.B(n_8178),
.Y(n_9789)
);

AND2x2_ASAP7_75t_L g9790 ( 
.A(n_8825),
.B(n_8202),
.Y(n_9790)
);

INVx1_ASAP7_75t_L g9791 ( 
.A(n_8827),
.Y(n_9791)
);

AND2x2_ASAP7_75t_L g9792 ( 
.A(n_8847),
.B(n_8202),
.Y(n_9792)
);

A2O1A1Ixp33_ASAP7_75t_L g9793 ( 
.A1(n_9517),
.A2(n_7857),
.B(n_7968),
.C(n_8511),
.Y(n_9793)
);

OR2x2_ASAP7_75t_L g9794 ( 
.A(n_8967),
.B(n_8344),
.Y(n_9794)
);

OAI22xp5_ASAP7_75t_L g9795 ( 
.A1(n_9091),
.A2(n_8043),
.B1(n_8327),
.B2(n_8001),
.Y(n_9795)
);

OAI21x1_ASAP7_75t_L g9796 ( 
.A1(n_9039),
.A2(n_8690),
.B(n_8604),
.Y(n_9796)
);

NOR2xp33_ASAP7_75t_L g9797 ( 
.A(n_9529),
.B(n_8157),
.Y(n_9797)
);

BUFx6f_ASAP7_75t_L g9798 ( 
.A(n_8900),
.Y(n_9798)
);

INVx2_ASAP7_75t_L g9799 ( 
.A(n_9139),
.Y(n_9799)
);

AO21x1_ASAP7_75t_SL g9800 ( 
.A1(n_9681),
.A2(n_7830),
.B(n_8455),
.Y(n_9800)
);

OAI21xp5_ASAP7_75t_L g9801 ( 
.A1(n_9325),
.A2(n_8729),
.B(n_8043),
.Y(n_9801)
);

AOI221xp5_ASAP7_75t_L g9802 ( 
.A1(n_9611),
.A2(n_8224),
.B1(n_8001),
.B2(n_8466),
.C(n_8321),
.Y(n_9802)
);

A2O1A1Ixp33_ASAP7_75t_L g9803 ( 
.A1(n_9303),
.A2(n_7801),
.B(n_8012),
.C(n_8273),
.Y(n_9803)
);

NAND2xp5_ASAP7_75t_L g9804 ( 
.A(n_9027),
.B(n_7978),
.Y(n_9804)
);

AO32x2_ASAP7_75t_L g9805 ( 
.A1(n_8873),
.A2(n_7929),
.A3(n_8488),
.B1(n_8610),
.B2(n_8616),
.Y(n_9805)
);

AND2x2_ASAP7_75t_L g9806 ( 
.A(n_8847),
.B(n_8202),
.Y(n_9806)
);

INVx2_ASAP7_75t_L g9807 ( 
.A(n_9139),
.Y(n_9807)
);

OAI22xp5_ASAP7_75t_L g9808 ( 
.A1(n_9509),
.A2(n_8327),
.B1(n_8466),
.B2(n_8273),
.Y(n_9808)
);

AOI21xp5_ASAP7_75t_L g9809 ( 
.A1(n_9007),
.A2(n_8012),
.B(n_7801),
.Y(n_9809)
);

AOI22xp5_ASAP7_75t_L g9810 ( 
.A1(n_8990),
.A2(n_8462),
.B1(n_8288),
.B2(n_7830),
.Y(n_9810)
);

OR2x2_ASAP7_75t_L g9811 ( 
.A(n_9590),
.B(n_8344),
.Y(n_9811)
);

CKINVDCx11_ASAP7_75t_R g9812 ( 
.A(n_9529),
.Y(n_9812)
);

HB1xp67_ASAP7_75t_L g9813 ( 
.A(n_8829),
.Y(n_9813)
);

OAI21xp5_ASAP7_75t_L g9814 ( 
.A1(n_8929),
.A2(n_8371),
.B(n_8298),
.Y(n_9814)
);

AND2x2_ASAP7_75t_L g9815 ( 
.A(n_8903),
.B(n_8278),
.Y(n_9815)
);

INVx2_ASAP7_75t_SL g9816 ( 
.A(n_8900),
.Y(n_9816)
);

A2O1A1Ixp33_ASAP7_75t_L g9817 ( 
.A1(n_9459),
.A2(n_7801),
.B(n_8012),
.C(n_8298),
.Y(n_9817)
);

NOR2xp33_ASAP7_75t_L g9818 ( 
.A(n_9137),
.B(n_8570),
.Y(n_9818)
);

AND2x2_ASAP7_75t_L g9819 ( 
.A(n_8903),
.B(n_8278),
.Y(n_9819)
);

AO21x2_ASAP7_75t_L g9820 ( 
.A1(n_9541),
.A2(n_8468),
.B(n_8497),
.Y(n_9820)
);

INVx2_ASAP7_75t_SL g9821 ( 
.A(n_8900),
.Y(n_9821)
);

INVx5_ASAP7_75t_L g9822 ( 
.A(n_8900),
.Y(n_9822)
);

OR2x2_ASAP7_75t_L g9823 ( 
.A(n_9596),
.B(n_8841),
.Y(n_9823)
);

BUFx3_ASAP7_75t_L g9824 ( 
.A(n_9067),
.Y(n_9824)
);

AND2x2_ASAP7_75t_L g9825 ( 
.A(n_8915),
.B(n_8278),
.Y(n_9825)
);

BUFx12f_ASAP7_75t_L g9826 ( 
.A(n_9105),
.Y(n_9826)
);

OA21x2_ASAP7_75t_L g9827 ( 
.A1(n_9424),
.A2(n_8059),
.B(n_8053),
.Y(n_9827)
);

AND2x2_ASAP7_75t_L g9828 ( 
.A(n_8915),
.B(n_8294),
.Y(n_9828)
);

INVx3_ASAP7_75t_L g9829 ( 
.A(n_8861),
.Y(n_9829)
);

BUFx2_ASAP7_75t_L g9830 ( 
.A(n_9400),
.Y(n_9830)
);

BUFx2_ASAP7_75t_L g9831 ( 
.A(n_9400),
.Y(n_9831)
);

INVx2_ASAP7_75t_SL g9832 ( 
.A(n_9136),
.Y(n_9832)
);

OAI21xp5_ASAP7_75t_L g9833 ( 
.A1(n_8929),
.A2(n_8371),
.B(n_7979),
.Y(n_9833)
);

INVx2_ASAP7_75t_L g9834 ( 
.A(n_9171),
.Y(n_9834)
);

INVx3_ASAP7_75t_L g9835 ( 
.A(n_8861),
.Y(n_9835)
);

AND2x2_ASAP7_75t_L g9836 ( 
.A(n_8882),
.B(n_8294),
.Y(n_9836)
);

INVx1_ASAP7_75t_L g9837 ( 
.A(n_9051),
.Y(n_9837)
);

AND2x4_ASAP7_75t_L g9838 ( 
.A(n_9027),
.B(n_9112),
.Y(n_9838)
);

OR2x2_ASAP7_75t_L g9839 ( 
.A(n_8841),
.B(n_8357),
.Y(n_9839)
);

OAI211xp5_ASAP7_75t_SL g9840 ( 
.A1(n_9332),
.A2(n_8321),
.B(n_8085),
.C(n_8405),
.Y(n_9840)
);

AOI211xp5_ASAP7_75t_L g9841 ( 
.A1(n_9260),
.A2(n_8224),
.B(n_8497),
.C(n_8196),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_9065),
.Y(n_9842)
);

CKINVDCx6p67_ASAP7_75t_R g9843 ( 
.A(n_9311),
.Y(n_9843)
);

AND2x4_ASAP7_75t_L g9844 ( 
.A(n_9112),
.B(n_8076),
.Y(n_9844)
);

A2O1A1Ixp33_ASAP7_75t_L g9845 ( 
.A1(n_9218),
.A2(n_9547),
.B(n_9311),
.C(n_9503),
.Y(n_9845)
);

INVx4_ASAP7_75t_SL g9846 ( 
.A(n_9232),
.Y(n_9846)
);

OAI21x1_ASAP7_75t_L g9847 ( 
.A1(n_9039),
.A2(n_8690),
.B(n_8604),
.Y(n_9847)
);

NAND2xp5_ASAP7_75t_L g9848 ( 
.A(n_9152),
.B(n_8289),
.Y(n_9848)
);

AO21x2_ASAP7_75t_L g9849 ( 
.A1(n_9541),
.A2(n_8603),
.B(n_7861),
.Y(n_9849)
);

AOI22xp5_ASAP7_75t_L g9850 ( 
.A1(n_8990),
.A2(n_7871),
.B1(n_7979),
.B2(n_8675),
.Y(n_9850)
);

A2O1A1Ixp33_ASAP7_75t_L g9851 ( 
.A1(n_9311),
.A2(n_7871),
.B(n_8680),
.C(n_8675),
.Y(n_9851)
);

AND2x2_ASAP7_75t_L g9852 ( 
.A(n_8882),
.B(n_8294),
.Y(n_9852)
);

NOR2xp33_ASAP7_75t_L g9853 ( 
.A(n_9137),
.B(n_8570),
.Y(n_9853)
);

AND2x4_ASAP7_75t_L g9854 ( 
.A(n_9152),
.B(n_8076),
.Y(n_9854)
);

A2O1A1Ixp33_ASAP7_75t_L g9855 ( 
.A1(n_9311),
.A2(n_8680),
.B(n_8549),
.C(n_8405),
.Y(n_9855)
);

INVxp67_ASAP7_75t_L g9856 ( 
.A(n_9156),
.Y(n_9856)
);

AND2x2_ASAP7_75t_L g9857 ( 
.A(n_8882),
.B(n_8303),
.Y(n_9857)
);

AOI21xp5_ASAP7_75t_L g9858 ( 
.A1(n_9136),
.A2(n_7235),
.B(n_8020),
.Y(n_9858)
);

INVx1_ASAP7_75t_L g9859 ( 
.A(n_8827),
.Y(n_9859)
);

HB1xp67_ASAP7_75t_L g9860 ( 
.A(n_8832),
.Y(n_9860)
);

INVxp67_ASAP7_75t_L g9861 ( 
.A(n_9156),
.Y(n_9861)
);

AOI22xp5_ASAP7_75t_L g9862 ( 
.A1(n_9138),
.A2(n_8486),
.B1(n_8600),
.B2(n_8564),
.Y(n_9862)
);

AND2x2_ASAP7_75t_L g9863 ( 
.A(n_9043),
.B(n_8303),
.Y(n_9863)
);

AOI22xp5_ASAP7_75t_L g9864 ( 
.A1(n_9138),
.A2(n_8486),
.B1(n_8600),
.B2(n_8564),
.Y(n_9864)
);

AND2x2_ASAP7_75t_L g9865 ( 
.A(n_9043),
.B(n_8303),
.Y(n_9865)
);

AND2x2_ASAP7_75t_L g9866 ( 
.A(n_9043),
.B(n_8342),
.Y(n_9866)
);

OAI21xp5_ASAP7_75t_L g9867 ( 
.A1(n_8929),
.A2(n_8549),
.B(n_8487),
.Y(n_9867)
);

A2O1A1Ixp33_ASAP7_75t_L g9868 ( 
.A1(n_9311),
.A2(n_6785),
.B(n_8487),
.C(n_8634),
.Y(n_9868)
);

INVx4_ASAP7_75t_SL g9869 ( 
.A(n_9232),
.Y(n_9869)
);

AND2x2_ASAP7_75t_L g9870 ( 
.A(n_9151),
.B(n_8342),
.Y(n_9870)
);

AND2x2_ASAP7_75t_L g9871 ( 
.A(n_9151),
.B(n_8342),
.Y(n_9871)
);

NAND2xp5_ASAP7_75t_L g9872 ( 
.A(n_9161),
.B(n_8289),
.Y(n_9872)
);

INVx4_ASAP7_75t_L g9873 ( 
.A(n_9136),
.Y(n_9873)
);

AND2x2_ASAP7_75t_L g9874 ( 
.A(n_9151),
.B(n_8374),
.Y(n_9874)
);

OAI22xp5_ASAP7_75t_L g9875 ( 
.A1(n_9593),
.A2(n_8108),
.B1(n_6920),
.B2(n_6921),
.Y(n_9875)
);

OAI22xp5_ASAP7_75t_L g9876 ( 
.A1(n_9460),
.A2(n_8108),
.B1(n_6920),
.B2(n_6921),
.Y(n_9876)
);

AOI22xp5_ASAP7_75t_L g9877 ( 
.A1(n_9138),
.A2(n_8486),
.B1(n_8600),
.B2(n_8564),
.Y(n_9877)
);

AND2x2_ASAP7_75t_L g9878 ( 
.A(n_9204),
.B(n_8374),
.Y(n_9878)
);

AND2x4_ASAP7_75t_L g9879 ( 
.A(n_9161),
.B(n_8076),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_8836),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_8836),
.Y(n_9881)
);

NOR2x1_ASAP7_75t_L g9882 ( 
.A(n_9454),
.B(n_6702),
.Y(n_9882)
);

INVx3_ASAP7_75t_L g9883 ( 
.A(n_9204),
.Y(n_9883)
);

A2O1A1Ixp33_ASAP7_75t_L g9884 ( 
.A1(n_8867),
.A2(n_8634),
.B(n_8652),
.C(n_7568),
.Y(n_9884)
);

INVx2_ASAP7_75t_L g9885 ( 
.A(n_9171),
.Y(n_9885)
);

A2O1A1Ixp33_ASAP7_75t_L g9886 ( 
.A1(n_9454),
.A2(n_8652),
.B(n_7568),
.C(n_8388),
.Y(n_9886)
);

CKINVDCx5p33_ASAP7_75t_R g9887 ( 
.A(n_9105),
.Y(n_9887)
);

AND2x2_ASAP7_75t_L g9888 ( 
.A(n_9204),
.B(n_9211),
.Y(n_9888)
);

CKINVDCx20_ASAP7_75t_R g9889 ( 
.A(n_9609),
.Y(n_9889)
);

O2A1O1Ixp33_ASAP7_75t_SL g9890 ( 
.A1(n_9223),
.A2(n_7215),
.B(n_8576),
.C(n_8406),
.Y(n_9890)
);

OR2x2_ASAP7_75t_L g9891 ( 
.A(n_8916),
.B(n_8357),
.Y(n_9891)
);

HB1xp67_ASAP7_75t_L g9892 ( 
.A(n_8923),
.Y(n_9892)
);

INVx2_ASAP7_75t_L g9893 ( 
.A(n_9171),
.Y(n_9893)
);

AND2x2_ASAP7_75t_L g9894 ( 
.A(n_9211),
.B(n_8374),
.Y(n_9894)
);

NAND2xp5_ASAP7_75t_L g9895 ( 
.A(n_9185),
.B(n_8300),
.Y(n_9895)
);

AOI22xp5_ASAP7_75t_L g9896 ( 
.A1(n_8934),
.A2(n_8486),
.B1(n_8600),
.B2(n_8564),
.Y(n_9896)
);

O2A1O1Ixp33_ASAP7_75t_L g9897 ( 
.A1(n_9541),
.A2(n_8196),
.B(n_7124),
.C(n_8677),
.Y(n_9897)
);

AND2x2_ASAP7_75t_L g9898 ( 
.A(n_9211),
.B(n_8388),
.Y(n_9898)
);

INVx1_ASAP7_75t_L g9899 ( 
.A(n_9068),
.Y(n_9899)
);

INVxp67_ASAP7_75t_L g9900 ( 
.A(n_9185),
.Y(n_9900)
);

INVx2_ASAP7_75t_SL g9901 ( 
.A(n_9136),
.Y(n_9901)
);

AOI22xp33_ASAP7_75t_L g9902 ( 
.A1(n_8843),
.A2(n_8136),
.B1(n_8033),
.B2(n_7971),
.Y(n_9902)
);

A2O1A1Ixp33_ASAP7_75t_L g9903 ( 
.A1(n_9519),
.A2(n_8423),
.B(n_8445),
.C(n_8388),
.Y(n_9903)
);

HB1xp67_ASAP7_75t_L g9904 ( 
.A(n_8947),
.Y(n_9904)
);

AND2x2_ASAP7_75t_L g9905 ( 
.A(n_9200),
.B(n_8423),
.Y(n_9905)
);

INVx2_ASAP7_75t_L g9906 ( 
.A(n_9171),
.Y(n_9906)
);

AND2x4_ASAP7_75t_L g9907 ( 
.A(n_9200),
.B(n_9472),
.Y(n_9907)
);

INVx1_ASAP7_75t_L g9908 ( 
.A(n_8837),
.Y(n_9908)
);

AND2x4_ASAP7_75t_L g9909 ( 
.A(n_9472),
.B(n_8076),
.Y(n_9909)
);

INVx1_ASAP7_75t_L g9910 ( 
.A(n_8837),
.Y(n_9910)
);

AOI221xp5_ASAP7_75t_L g9911 ( 
.A1(n_8818),
.A2(n_8085),
.B1(n_7516),
.B2(n_8039),
.C(n_8020),
.Y(n_9911)
);

OA21x2_ASAP7_75t_L g9912 ( 
.A1(n_9424),
.A2(n_8059),
.B(n_8053),
.Y(n_9912)
);

NOR2x1_ASAP7_75t_SL g9913 ( 
.A(n_8818),
.B(n_8033),
.Y(n_9913)
);

NAND2xp5_ASAP7_75t_SL g9914 ( 
.A(n_9472),
.B(n_8076),
.Y(n_9914)
);

AO32x2_ASAP7_75t_L g9915 ( 
.A1(n_8894),
.A2(n_7690),
.A3(n_7517),
.B1(n_8274),
.B2(n_8077),
.Y(n_9915)
);

AOI221xp5_ASAP7_75t_L g9916 ( 
.A1(n_8934),
.A2(n_8039),
.B1(n_8020),
.B2(n_8512),
.C(n_8499),
.Y(n_9916)
);

NAND2xp5_ASAP7_75t_L g9917 ( 
.A(n_8975),
.B(n_8300),
.Y(n_9917)
);

AND2x2_ASAP7_75t_SL g9918 ( 
.A(n_8853),
.B(n_6960),
.Y(n_9918)
);

OAI22xp5_ASAP7_75t_SL g9919 ( 
.A1(n_9232),
.A2(n_7113),
.B1(n_7018),
.B2(n_7035),
.Y(n_9919)
);

AND2x2_ASAP7_75t_L g9920 ( 
.A(n_9337),
.B(n_9455),
.Y(n_9920)
);

INVx2_ASAP7_75t_L g9921 ( 
.A(n_9171),
.Y(n_9921)
);

NOR2x1_ASAP7_75t_SL g9922 ( 
.A(n_8815),
.B(n_8136),
.Y(n_9922)
);

AND2x2_ASAP7_75t_L g9923 ( 
.A(n_9337),
.B(n_8423),
.Y(n_9923)
);

BUFx6f_ASAP7_75t_L g9924 ( 
.A(n_9136),
.Y(n_9924)
);

OAI22xp5_ASAP7_75t_L g9925 ( 
.A1(n_9356),
.A2(n_6788),
.B1(n_7243),
.B2(n_6991),
.Y(n_9925)
);

INVx1_ASAP7_75t_L g9926 ( 
.A(n_9083),
.Y(n_9926)
);

OA21x2_ASAP7_75t_L g9927 ( 
.A1(n_9084),
.A2(n_8069),
.B(n_8059),
.Y(n_9927)
);

OAI22xp5_ASAP7_75t_L g9928 ( 
.A1(n_8983),
.A2(n_6788),
.B1(n_7243),
.B2(n_6913),
.Y(n_9928)
);

INVx2_ASAP7_75t_L g9929 ( 
.A(n_9247),
.Y(n_9929)
);

AND2x2_ASAP7_75t_L g9930 ( 
.A(n_9337),
.B(n_8445),
.Y(n_9930)
);

OAI22xp5_ASAP7_75t_L g9931 ( 
.A1(n_8983),
.A2(n_6901),
.B1(n_6913),
.B2(n_7150),
.Y(n_9931)
);

OAI22xp5_ASAP7_75t_L g9932 ( 
.A1(n_8983),
.A2(n_6901),
.B1(n_7219),
.B2(n_7183),
.Y(n_9932)
);

NOR2xp33_ASAP7_75t_L g9933 ( 
.A(n_9463),
.B(n_8427),
.Y(n_9933)
);

OAI22xp33_ASAP7_75t_SL g9934 ( 
.A1(n_9223),
.A2(n_7977),
.B1(n_8252),
.B2(n_8058),
.Y(n_9934)
);

AND2x2_ASAP7_75t_L g9935 ( 
.A(n_9337),
.B(n_8445),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_9085),
.Y(n_9936)
);

NOR2xp33_ASAP7_75t_L g9937 ( 
.A(n_9463),
.B(n_8624),
.Y(n_9937)
);

AND2x2_ASAP7_75t_L g9938 ( 
.A(n_9455),
.B(n_8469),
.Y(n_9938)
);

OR2x2_ASAP7_75t_L g9939 ( 
.A(n_8964),
.B(n_8357),
.Y(n_9939)
);

INVx1_ASAP7_75t_L g9940 ( 
.A(n_8838),
.Y(n_9940)
);

AO32x2_ASAP7_75t_L g9941 ( 
.A1(n_8894),
.A2(n_7690),
.A3(n_7517),
.B1(n_8274),
.B2(n_8077),
.Y(n_9941)
);

INVx1_ASAP7_75t_L g9942 ( 
.A(n_8838),
.Y(n_9942)
);

INVxp67_ASAP7_75t_SL g9943 ( 
.A(n_9329),
.Y(n_9943)
);

NAND3xp33_ASAP7_75t_L g9944 ( 
.A(n_8890),
.B(n_8677),
.C(n_8393),
.Y(n_9944)
);

AND2x2_ASAP7_75t_L g9945 ( 
.A(n_9455),
.B(n_8469),
.Y(n_9945)
);

BUFx2_ASAP7_75t_L g9946 ( 
.A(n_9519),
.Y(n_9946)
);

INVx2_ASAP7_75t_L g9947 ( 
.A(n_9247),
.Y(n_9947)
);

INVxp67_ASAP7_75t_L g9948 ( 
.A(n_9247),
.Y(n_9948)
);

AO21x2_ASAP7_75t_L g9949 ( 
.A1(n_9329),
.A2(n_8603),
.B(n_7861),
.Y(n_9949)
);

BUFx2_ASAP7_75t_L g9950 ( 
.A(n_9557),
.Y(n_9950)
);

INVxp33_ASAP7_75t_L g9951 ( 
.A(n_9642),
.Y(n_9951)
);

HB1xp67_ASAP7_75t_L g9952 ( 
.A(n_9125),
.Y(n_9952)
);

AO32x2_ASAP7_75t_L g9953 ( 
.A1(n_9092),
.A2(n_8447),
.A3(n_8552),
.B1(n_8274),
.B2(n_8077),
.Y(n_9953)
);

NAND2xp5_ASAP7_75t_L g9954 ( 
.A(n_9090),
.B(n_8432),
.Y(n_9954)
);

AND2x2_ASAP7_75t_L g9955 ( 
.A(n_9677),
.B(n_8469),
.Y(n_9955)
);

NAND2xp5_ASAP7_75t_L g9956 ( 
.A(n_9504),
.B(n_8432),
.Y(n_9956)
);

AO21x1_ASAP7_75t_L g9957 ( 
.A1(n_9182),
.A2(n_8274),
.B(n_8077),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_9247),
.Y(n_9958)
);

OA21x2_ASAP7_75t_L g9959 ( 
.A1(n_9084),
.A2(n_8070),
.B(n_8069),
.Y(n_9959)
);

OAI22xp5_ASAP7_75t_L g9960 ( 
.A1(n_8983),
.A2(n_7219),
.B1(n_7244),
.B2(n_7183),
.Y(n_9960)
);

AOI221xp5_ASAP7_75t_L g9961 ( 
.A1(n_8934),
.A2(n_9403),
.B1(n_9429),
.B2(n_8910),
.C(n_8846),
.Y(n_9961)
);

INVx3_ASAP7_75t_L g9962 ( 
.A(n_9682),
.Y(n_9962)
);

INVx2_ASAP7_75t_L g9963 ( 
.A(n_9247),
.Y(n_9963)
);

NOR2xp33_ASAP7_75t_L g9964 ( 
.A(n_9534),
.B(n_8624),
.Y(n_9964)
);

INVx4_ASAP7_75t_L g9965 ( 
.A(n_9106),
.Y(n_9965)
);

A2O1A1Ixp33_ASAP7_75t_L g9966 ( 
.A1(n_9557),
.A2(n_8531),
.B(n_8577),
.C(n_8526),
.Y(n_9966)
);

AOI22xp5_ASAP7_75t_L g9967 ( 
.A1(n_9120),
.A2(n_8564),
.B1(n_8600),
.B2(n_8486),
.Y(n_9967)
);

INVx2_ASAP7_75t_L g9968 ( 
.A(n_9354),
.Y(n_9968)
);

A2O1A1Ixp33_ASAP7_75t_L g9969 ( 
.A1(n_9610),
.A2(n_8531),
.B(n_8577),
.C(n_8526),
.Y(n_9969)
);

O2A1O1Ixp33_ASAP7_75t_L g9970 ( 
.A1(n_9260),
.A2(n_8890),
.B(n_9333),
.C(n_9403),
.Y(n_9970)
);

NAND2xp5_ASAP7_75t_L g9971 ( 
.A(n_9545),
.B(n_8609),
.Y(n_9971)
);

AND2x2_ASAP7_75t_L g9972 ( 
.A(n_9677),
.B(n_8526),
.Y(n_9972)
);

A2O1A1Ixp33_ASAP7_75t_L g9973 ( 
.A1(n_9610),
.A2(n_8577),
.B(n_8638),
.C(n_8531),
.Y(n_9973)
);

AND2x2_ASAP7_75t_L g9974 ( 
.A(n_9684),
.B(n_8638),
.Y(n_9974)
);

AOI22xp33_ASAP7_75t_L g9975 ( 
.A1(n_8843),
.A2(n_8136),
.B1(n_7971),
.B2(n_7828),
.Y(n_9975)
);

BUFx4f_ASAP7_75t_L g9976 ( 
.A(n_9354),
.Y(n_9976)
);

AND2x2_ASAP7_75t_L g9977 ( 
.A(n_9684),
.B(n_9661),
.Y(n_9977)
);

OAI21xp5_ASAP7_75t_L g9978 ( 
.A1(n_8890),
.A2(n_8677),
.B(n_8603),
.Y(n_9978)
);

AND2x2_ASAP7_75t_L g9979 ( 
.A(n_9661),
.B(n_8638),
.Y(n_9979)
);

OA21x2_ASAP7_75t_L g9980 ( 
.A1(n_9462),
.A2(n_8070),
.B(n_8069),
.Y(n_9980)
);

INVx6_ASAP7_75t_SL g9981 ( 
.A(n_9056),
.Y(n_9981)
);

O2A1O1Ixp33_ASAP7_75t_L g9982 ( 
.A1(n_8890),
.A2(n_8677),
.B(n_7832),
.C(n_7932),
.Y(n_9982)
);

NOR2xp33_ASAP7_75t_R g9983 ( 
.A(n_9106),
.B(n_9534),
.Y(n_9983)
);

OR2x2_ASAP7_75t_L g9984 ( 
.A(n_9193),
.B(n_8609),
.Y(n_9984)
);

OR2x6_ASAP7_75t_L g9985 ( 
.A(n_9277),
.B(n_7977),
.Y(n_9985)
);

AND2x2_ASAP7_75t_L g9986 ( 
.A(n_9682),
.B(n_8673),
.Y(n_9986)
);

OAI21x1_ASAP7_75t_L g9987 ( 
.A1(n_8865),
.A2(n_8690),
.B(n_8604),
.Y(n_9987)
);

AND2x2_ASAP7_75t_L g9988 ( 
.A(n_9682),
.B(n_8673),
.Y(n_9988)
);

OA21x2_ASAP7_75t_L g9989 ( 
.A1(n_9462),
.A2(n_8074),
.B(n_8070),
.Y(n_9989)
);

INVx4_ASAP7_75t_L g9990 ( 
.A(n_9279),
.Y(n_9990)
);

OAI22xp5_ASAP7_75t_L g9991 ( 
.A1(n_9056),
.A2(n_7219),
.B1(n_7244),
.B2(n_7183),
.Y(n_9991)
);

INVx1_ASAP7_75t_L g9992 ( 
.A(n_9132),
.Y(n_9992)
);

OAI21xp5_ASAP7_75t_L g9993 ( 
.A1(n_8863),
.A2(n_8677),
.B(n_8585),
.Y(n_9993)
);

NAND2xp5_ASAP7_75t_L g9994 ( 
.A(n_9690),
.B(n_8631),
.Y(n_9994)
);

INVx1_ASAP7_75t_L g9995 ( 
.A(n_8839),
.Y(n_9995)
);

NAND4xp25_ASAP7_75t_L g9996 ( 
.A(n_9102),
.B(n_8434),
.C(n_8376),
.D(n_6879),
.Y(n_9996)
);

OR2x6_ASAP7_75t_L g9997 ( 
.A(n_9277),
.B(n_8058),
.Y(n_9997)
);

INVx2_ASAP7_75t_L g9998 ( 
.A(n_9354),
.Y(n_9998)
);

AND2x2_ASAP7_75t_L g9999 ( 
.A(n_9225),
.B(n_8673),
.Y(n_9999)
);

AND2x2_ASAP7_75t_L g10000 ( 
.A(n_9225),
.B(n_8713),
.Y(n_10000)
);

INVx2_ASAP7_75t_L g10001 ( 
.A(n_9354),
.Y(n_10001)
);

A2O1A1Ixp33_ASAP7_75t_L g10002 ( 
.A1(n_9612),
.A2(n_8718),
.B(n_8751),
.C(n_8713),
.Y(n_10002)
);

A2O1A1Ixp33_ASAP7_75t_L g10003 ( 
.A1(n_9612),
.A2(n_8718),
.B(n_8751),
.C(n_8713),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_8839),
.Y(n_10004)
);

AO32x2_ASAP7_75t_L g10005 ( 
.A1(n_9092),
.A2(n_8447),
.A3(n_8552),
.B1(n_8274),
.B2(n_8077),
.Y(n_10005)
);

OR2x2_ASAP7_75t_L g10006 ( 
.A(n_9158),
.B(n_8631),
.Y(n_10006)
);

OAI21xp5_ASAP7_75t_L g10007 ( 
.A1(n_8863),
.A2(n_8585),
.B(n_8523),
.Y(n_10007)
);

OAI22xp5_ASAP7_75t_L g10008 ( 
.A1(n_9056),
.A2(n_7244),
.B1(n_6908),
.B2(n_7426),
.Y(n_10008)
);

AND2x2_ASAP7_75t_L g10009 ( 
.A(n_9588),
.B(n_8718),
.Y(n_10009)
);

AO21x2_ASAP7_75t_L g10010 ( 
.A1(n_9333),
.A2(n_7861),
.B(n_8198),
.Y(n_10010)
);

AND2x2_ASAP7_75t_L g10011 ( 
.A(n_9588),
.B(n_9627),
.Y(n_10011)
);

OAI21x1_ASAP7_75t_L g10012 ( 
.A1(n_8865),
.A2(n_8706),
.B(n_8690),
.Y(n_10012)
);

INVxp67_ASAP7_75t_SL g10013 ( 
.A(n_9182),
.Y(n_10013)
);

AO32x1_ASAP7_75t_L g10014 ( 
.A1(n_9099),
.A2(n_8447),
.A3(n_8762),
.B1(n_8552),
.B2(n_6867),
.Y(n_10014)
);

AND2x4_ASAP7_75t_L g10015 ( 
.A(n_9472),
.B(n_8447),
.Y(n_10015)
);

NAND4xp25_ASAP7_75t_L g10016 ( 
.A(n_9276),
.B(n_8376),
.C(n_8434),
.D(n_7202),
.Y(n_10016)
);

BUFx3_ASAP7_75t_L g10017 ( 
.A(n_9406),
.Y(n_10017)
);

OAI22xp5_ASAP7_75t_L g10018 ( 
.A1(n_9056),
.A2(n_7426),
.B1(n_7172),
.B2(n_7199),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_8842),
.Y(n_10019)
);

CKINVDCx11_ASAP7_75t_R g10020 ( 
.A(n_9526),
.Y(n_10020)
);

AOI22xp5_ASAP7_75t_L g10021 ( 
.A1(n_9120),
.A2(n_7927),
.B1(n_8559),
.B2(n_6761),
.Y(n_10021)
);

OAI21xp5_ASAP7_75t_L g10022 ( 
.A1(n_8863),
.A2(n_8585),
.B(n_8523),
.Y(n_10022)
);

AOI22xp5_ASAP7_75t_L g10023 ( 
.A1(n_9120),
.A2(n_8559),
.B1(n_7927),
.B2(n_7326),
.Y(n_10023)
);

INVx2_ASAP7_75t_L g10024 ( 
.A(n_9354),
.Y(n_10024)
);

AO32x2_ASAP7_75t_L g10025 ( 
.A1(n_9099),
.A2(n_8762),
.A3(n_8552),
.B1(n_8447),
.B2(n_7821),
.Y(n_10025)
);

AND2x2_ASAP7_75t_L g10026 ( 
.A(n_9627),
.B(n_8751),
.Y(n_10026)
);

HB1xp67_ASAP7_75t_L g10027 ( 
.A(n_9176),
.Y(n_10027)
);

BUFx2_ASAP7_75t_L g10028 ( 
.A(n_8814),
.Y(n_10028)
);

NAND2xp5_ASAP7_75t_L g10029 ( 
.A(n_9145),
.B(n_8552),
.Y(n_10029)
);

O2A1O1Ixp33_ASAP7_75t_SL g10030 ( 
.A1(n_9145),
.A2(n_8592),
.B(n_8576),
.C(n_7832),
.Y(n_10030)
);

AO21x2_ASAP7_75t_L g10031 ( 
.A1(n_8815),
.A2(n_8199),
.B(n_8198),
.Y(n_10031)
);

OR2x2_ASAP7_75t_L g10032 ( 
.A(n_9158),
.B(n_8794),
.Y(n_10032)
);

AND2x2_ASAP7_75t_L g10033 ( 
.A(n_9663),
.B(n_8758),
.Y(n_10033)
);

AND2x4_ASAP7_75t_L g10034 ( 
.A(n_9472),
.B(n_8762),
.Y(n_10034)
);

AND2x2_ASAP7_75t_L g10035 ( 
.A(n_9663),
.B(n_8758),
.Y(n_10035)
);

INVx1_ASAP7_75t_L g10036 ( 
.A(n_9235),
.Y(n_10036)
);

AOI22xp5_ASAP7_75t_L g10037 ( 
.A1(n_9399),
.A2(n_8559),
.B1(n_7361),
.B2(n_7380),
.Y(n_10037)
);

INVx1_ASAP7_75t_L g10038 ( 
.A(n_8842),
.Y(n_10038)
);

AOI221xp5_ASAP7_75t_L g10039 ( 
.A1(n_9403),
.A2(n_8039),
.B1(n_8020),
.B2(n_8512),
.C(n_8499),
.Y(n_10039)
);

AND2x2_ASAP7_75t_L g10040 ( 
.A(n_9672),
.B(n_8758),
.Y(n_10040)
);

O2A1O1Ixp33_ASAP7_75t_L g10041 ( 
.A1(n_9429),
.A2(n_7821),
.B(n_7932),
.C(n_7832),
.Y(n_10041)
);

AND2x2_ASAP7_75t_L g10042 ( 
.A(n_9672),
.B(n_8221),
.Y(n_10042)
);

INVx1_ASAP7_75t_L g10043 ( 
.A(n_9238),
.Y(n_10043)
);

AOI22xp5_ASAP7_75t_L g10044 ( 
.A1(n_9399),
.A2(n_8559),
.B1(n_7361),
.B2(n_7380),
.Y(n_10044)
);

OA21x2_ASAP7_75t_L g10045 ( 
.A1(n_9573),
.A2(n_8080),
.B(n_8074),
.Y(n_10045)
);

A2O1A1Ixp33_ASAP7_75t_L g10046 ( 
.A1(n_8830),
.A2(n_6702),
.B(n_6724),
.C(n_7202),
.Y(n_10046)
);

AND2x2_ASAP7_75t_L g10047 ( 
.A(n_9141),
.B(n_8221),
.Y(n_10047)
);

INVx1_ASAP7_75t_L g10048 ( 
.A(n_9243),
.Y(n_10048)
);

AND2x6_ASAP7_75t_L g10049 ( 
.A(n_8933),
.B(n_6724),
.Y(n_10049)
);

HB1xp67_ASAP7_75t_L g10050 ( 
.A(n_9253),
.Y(n_10050)
);

INVx4_ASAP7_75t_L g10051 ( 
.A(n_9279),
.Y(n_10051)
);

INVxp67_ASAP7_75t_L g10052 ( 
.A(n_9368),
.Y(n_10052)
);

AOI22xp33_ASAP7_75t_SL g10053 ( 
.A1(n_8910),
.A2(n_8858),
.B1(n_8846),
.B2(n_8863),
.Y(n_10053)
);

AO32x1_ASAP7_75t_L g10054 ( 
.A1(n_9199),
.A2(n_8762),
.A3(n_6867),
.B1(n_6857),
.B2(n_7932),
.Y(n_10054)
);

O2A1O1Ixp33_ASAP7_75t_SL g10055 ( 
.A1(n_9199),
.A2(n_8592),
.B(n_7955),
.C(n_7987),
.Y(n_10055)
);

INVx2_ASAP7_75t_L g10056 ( 
.A(n_9368),
.Y(n_10056)
);

AND2x4_ASAP7_75t_L g10057 ( 
.A(n_9472),
.B(n_9629),
.Y(n_10057)
);

AND2x2_ASAP7_75t_L g10058 ( 
.A(n_9141),
.B(n_8221),
.Y(n_10058)
);

INVx1_ASAP7_75t_L g10059 ( 
.A(n_8844),
.Y(n_10059)
);

NOR2x1_ASAP7_75t_R g10060 ( 
.A(n_9306),
.B(n_7072),
.Y(n_10060)
);

NAND2x1_ASAP7_75t_L g10061 ( 
.A(n_8932),
.B(n_7820),
.Y(n_10061)
);

AOI22xp5_ASAP7_75t_L g10062 ( 
.A1(n_9399),
.A2(n_8910),
.B1(n_9042),
.B2(n_9009),
.Y(n_10062)
);

OA21x2_ASAP7_75t_L g10063 ( 
.A1(n_9573),
.A2(n_8080),
.B(n_8074),
.Y(n_10063)
);

NAND2xp5_ASAP7_75t_SL g10064 ( 
.A(n_9629),
.B(n_8762),
.Y(n_10064)
);

OAI21xp5_ASAP7_75t_L g10065 ( 
.A1(n_9449),
.A2(n_8656),
.B(n_8523),
.Y(n_10065)
);

AND2x2_ASAP7_75t_L g10066 ( 
.A(n_9141),
.B(n_7901),
.Y(n_10066)
);

INVx1_ASAP7_75t_L g10067 ( 
.A(n_8844),
.Y(n_10067)
);

INVx1_ASAP7_75t_L g10068 ( 
.A(n_8850),
.Y(n_10068)
);

AND2x2_ASAP7_75t_L g10069 ( 
.A(n_9141),
.B(n_7901),
.Y(n_10069)
);

OA21x2_ASAP7_75t_L g10070 ( 
.A1(n_9589),
.A2(n_8084),
.B(n_8080),
.Y(n_10070)
);

OAI21x1_ASAP7_75t_L g10071 ( 
.A1(n_8907),
.A2(n_8706),
.B(n_7829),
.Y(n_10071)
);

OR2x6_ASAP7_75t_L g10072 ( 
.A(n_9352),
.B(n_8058),
.Y(n_10072)
);

A2O1A1Ixp33_ASAP7_75t_L g10073 ( 
.A1(n_8933),
.A2(n_8676),
.B(n_8656),
.C(n_8800),
.Y(n_10073)
);

O2A1O1Ixp33_ASAP7_75t_SL g10074 ( 
.A1(n_9205),
.A2(n_9227),
.B(n_9287),
.C(n_9215),
.Y(n_10074)
);

OR2x2_ASAP7_75t_L g10075 ( 
.A(n_9579),
.B(n_8794),
.Y(n_10075)
);

NOR2xp33_ASAP7_75t_L g10076 ( 
.A(n_8949),
.B(n_8607),
.Y(n_10076)
);

NAND2xp5_ASAP7_75t_SL g10077 ( 
.A(n_9629),
.B(n_9276),
.Y(n_10077)
);

AND2x2_ASAP7_75t_L g10078 ( 
.A(n_9202),
.B(n_7901),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9285),
.Y(n_10079)
);

AND2x2_ASAP7_75t_L g10080 ( 
.A(n_9202),
.B(n_7901),
.Y(n_10080)
);

AND2x2_ASAP7_75t_L g10081 ( 
.A(n_9202),
.B(n_7901),
.Y(n_10081)
);

OR2x2_ASAP7_75t_L g10082 ( 
.A(n_9626),
.B(n_8794),
.Y(n_10082)
);

INVxp67_ASAP7_75t_L g10083 ( 
.A(n_9368),
.Y(n_10083)
);

AND2x2_ASAP7_75t_L g10084 ( 
.A(n_9202),
.B(n_7904),
.Y(n_10084)
);

OAI22xp5_ASAP7_75t_SL g10085 ( 
.A1(n_9306),
.A2(n_7113),
.B1(n_7018),
.B2(n_7035),
.Y(n_10085)
);

NOR2x1p5_ASAP7_75t_L g10086 ( 
.A(n_8949),
.B(n_8734),
.Y(n_10086)
);

INVx1_ASAP7_75t_L g10087 ( 
.A(n_8850),
.Y(n_10087)
);

INVx1_ASAP7_75t_L g10088 ( 
.A(n_8855),
.Y(n_10088)
);

AND2x2_ASAP7_75t_L g10089 ( 
.A(n_9323),
.B(n_7904),
.Y(n_10089)
);

OAI21xp5_ASAP7_75t_L g10090 ( 
.A1(n_9449),
.A2(n_8676),
.B(n_8656),
.Y(n_10090)
);

A2O1A1Ixp33_ASAP7_75t_L g10091 ( 
.A1(n_9014),
.A2(n_8676),
.B(n_8800),
.C(n_7049),
.Y(n_10091)
);

OAI22xp5_ASAP7_75t_L g10092 ( 
.A1(n_9323),
.A2(n_9382),
.B1(n_7171),
.B2(n_7518),
.Y(n_10092)
);

AO32x2_ASAP7_75t_L g10093 ( 
.A1(n_9205),
.A2(n_7821),
.A3(n_8017),
.B1(n_7987),
.B2(n_7955),
.Y(n_10093)
);

INVx2_ASAP7_75t_L g10094 ( 
.A(n_9368),
.Y(n_10094)
);

NAND2xp33_ASAP7_75t_L g10095 ( 
.A(n_9368),
.B(n_8285),
.Y(n_10095)
);

INVx2_ASAP7_75t_L g10096 ( 
.A(n_9410),
.Y(n_10096)
);

HB1xp67_ASAP7_75t_L g10097 ( 
.A(n_9328),
.Y(n_10097)
);

OA21x2_ASAP7_75t_L g10098 ( 
.A1(n_9589),
.A2(n_8088),
.B(n_8084),
.Y(n_10098)
);

HB1xp67_ASAP7_75t_L g10099 ( 
.A(n_9343),
.Y(n_10099)
);

OAI21xp5_ASAP7_75t_L g10100 ( 
.A1(n_9449),
.A2(n_8733),
.B(n_8722),
.Y(n_10100)
);

OR2x6_ASAP7_75t_L g10101 ( 
.A(n_9352),
.B(n_8058),
.Y(n_10101)
);

NOR2xp33_ASAP7_75t_L g10102 ( 
.A(n_9014),
.B(n_6866),
.Y(n_10102)
);

HB1xp67_ASAP7_75t_L g10103 ( 
.A(n_9364),
.Y(n_10103)
);

INVx1_ASAP7_75t_L g10104 ( 
.A(n_9367),
.Y(n_10104)
);

OAI21xp5_ASAP7_75t_L g10105 ( 
.A1(n_9449),
.A2(n_8733),
.B(n_8722),
.Y(n_10105)
);

NOR2x1_ASAP7_75t_SL g10106 ( 
.A(n_8846),
.B(n_7828),
.Y(n_10106)
);

INVx2_ASAP7_75t_L g10107 ( 
.A(n_9410),
.Y(n_10107)
);

AOI22xp33_ASAP7_75t_L g10108 ( 
.A1(n_9251),
.A2(n_7971),
.B1(n_7828),
.B2(n_8020),
.Y(n_10108)
);

INVxp33_ASAP7_75t_SL g10109 ( 
.A(n_9095),
.Y(n_10109)
);

AND2x2_ASAP7_75t_L g10110 ( 
.A(n_9323),
.B(n_7904),
.Y(n_10110)
);

AND2x2_ASAP7_75t_L g10111 ( 
.A(n_9323),
.B(n_9382),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_8855),
.Y(n_10112)
);

OA21x2_ASAP7_75t_L g10113 ( 
.A1(n_9594),
.A2(n_8088),
.B(n_8084),
.Y(n_10113)
);

CKINVDCx6p67_ASAP7_75t_R g10114 ( 
.A(n_9095),
.Y(n_10114)
);

OAI21x1_ASAP7_75t_SL g10115 ( 
.A1(n_9387),
.A2(n_6971),
.B(n_6960),
.Y(n_10115)
);

BUFx4f_ASAP7_75t_L g10116 ( 
.A(n_9410),
.Y(n_10116)
);

BUFx3_ASAP7_75t_L g10117 ( 
.A(n_9115),
.Y(n_10117)
);

AOI21x1_ASAP7_75t_L g10118 ( 
.A1(n_9245),
.A2(n_8566),
.B(n_8558),
.Y(n_10118)
);

OAI22xp5_ASAP7_75t_L g10119 ( 
.A1(n_9382),
.A2(n_7518),
.B1(n_7217),
.B2(n_7492),
.Y(n_10119)
);

AND2x2_ASAP7_75t_L g10120 ( 
.A(n_9382),
.B(n_7904),
.Y(n_10120)
);

NOR2x1_ASAP7_75t_SL g10121 ( 
.A(n_9052),
.B(n_8448),
.Y(n_10121)
);

AND2x4_ASAP7_75t_L g10122 ( 
.A(n_9629),
.B(n_8346),
.Y(n_10122)
);

AOI21xp5_ASAP7_75t_L g10123 ( 
.A1(n_9429),
.A2(n_8039),
.B(n_8413),
.Y(n_10123)
);

OR2x2_ASAP7_75t_L g10124 ( 
.A(n_9651),
.B(n_5956),
.Y(n_10124)
);

AND2x4_ASAP7_75t_L g10125 ( 
.A(n_9629),
.B(n_8346),
.Y(n_10125)
);

AND2x2_ASAP7_75t_L g10126 ( 
.A(n_9476),
.B(n_7904),
.Y(n_10126)
);

BUFx6f_ASAP7_75t_L g10127 ( 
.A(n_9115),
.Y(n_10127)
);

AND2x2_ASAP7_75t_L g10128 ( 
.A(n_9476),
.B(n_7913),
.Y(n_10128)
);

OAI21x1_ASAP7_75t_L g10129 ( 
.A1(n_8907),
.A2(n_8706),
.B(n_7829),
.Y(n_10129)
);

AND2x2_ASAP7_75t_L g10130 ( 
.A(n_9476),
.B(n_7913),
.Y(n_10130)
);

INVx1_ASAP7_75t_L g10131 ( 
.A(n_8857),
.Y(n_10131)
);

AOI21xp5_ASAP7_75t_SL g10132 ( 
.A1(n_9128),
.A2(n_7050),
.B(n_7049),
.Y(n_10132)
);

AOI21x1_ASAP7_75t_L g10133 ( 
.A1(n_9245),
.A2(n_8566),
.B(n_8558),
.Y(n_10133)
);

AND2x2_ASAP7_75t_L g10134 ( 
.A(n_9629),
.B(n_7913),
.Y(n_10134)
);

AND2x2_ASAP7_75t_L g10135 ( 
.A(n_9365),
.B(n_9369),
.Y(n_10135)
);

AND2x2_ASAP7_75t_L g10136 ( 
.A(n_9365),
.B(n_9369),
.Y(n_10136)
);

INVx2_ASAP7_75t_L g10137 ( 
.A(n_9410),
.Y(n_10137)
);

INVx2_ASAP7_75t_L g10138 ( 
.A(n_9410),
.Y(n_10138)
);

AND2x2_ASAP7_75t_L g10139 ( 
.A(n_9396),
.B(n_7913),
.Y(n_10139)
);

AND2x2_ASAP7_75t_L g10140 ( 
.A(n_9396),
.B(n_7913),
.Y(n_10140)
);

AND2x2_ASAP7_75t_L g10141 ( 
.A(n_9430),
.B(n_7919),
.Y(n_10141)
);

BUFx2_ASAP7_75t_L g10142 ( 
.A(n_9128),
.Y(n_10142)
);

BUFx12f_ASAP7_75t_L g10143 ( 
.A(n_9231),
.Y(n_10143)
);

OAI22xp5_ASAP7_75t_L g10144 ( 
.A1(n_9564),
.A2(n_7518),
.B1(n_7217),
.B2(n_7492),
.Y(n_10144)
);

OR2x2_ASAP7_75t_L g10145 ( 
.A(n_9194),
.B(n_5956),
.Y(n_10145)
);

AOI221xp5_ASAP7_75t_L g10146 ( 
.A1(n_9278),
.A2(n_8039),
.B1(n_8512),
.B2(n_8499),
.C(n_8413),
.Y(n_10146)
);

NAND3xp33_ASAP7_75t_L g10147 ( 
.A(n_9473),
.B(n_8393),
.C(n_8261),
.Y(n_10147)
);

OA21x2_ASAP7_75t_L g10148 ( 
.A1(n_9594),
.A2(n_8089),
.B(n_8088),
.Y(n_10148)
);

CKINVDCx5p33_ASAP7_75t_R g10149 ( 
.A(n_9254),
.Y(n_10149)
);

NAND2xp5_ASAP7_75t_L g10150 ( 
.A(n_9215),
.B(n_6857),
.Y(n_10150)
);

A2O1A1Ixp33_ASAP7_75t_L g10151 ( 
.A1(n_9231),
.A2(n_8800),
.B(n_7049),
.C(n_7088),
.Y(n_10151)
);

OA21x2_ASAP7_75t_L g10152 ( 
.A1(n_9693),
.A2(n_8097),
.B(n_8089),
.Y(n_10152)
);

AOI22xp33_ASAP7_75t_L g10153 ( 
.A1(n_9251),
.A2(n_8448),
.B1(n_8393),
.B2(n_8413),
.Y(n_10153)
);

AND2x2_ASAP7_75t_L g10154 ( 
.A(n_9430),
.B(n_7919),
.Y(n_10154)
);

BUFx6f_ASAP7_75t_L g10155 ( 
.A(n_9239),
.Y(n_10155)
);

AND2x2_ASAP7_75t_L g10156 ( 
.A(n_9457),
.B(n_7919),
.Y(n_10156)
);

INVx1_ASAP7_75t_L g10157 ( 
.A(n_9395),
.Y(n_10157)
);

AND2x2_ASAP7_75t_L g10158 ( 
.A(n_9457),
.B(n_7919),
.Y(n_10158)
);

AO21x2_ASAP7_75t_L g10159 ( 
.A1(n_9387),
.A2(n_9282),
.B(n_9393),
.Y(n_10159)
);

OR2x2_ASAP7_75t_L g10160 ( 
.A(n_9194),
.B(n_8562),
.Y(n_10160)
);

INVx1_ASAP7_75t_L g10161 ( 
.A(n_8857),
.Y(n_10161)
);

NOR2x1_ASAP7_75t_SL g10162 ( 
.A(n_9052),
.B(n_8448),
.Y(n_10162)
);

NAND2xp5_ASAP7_75t_L g10163 ( 
.A(n_9227),
.B(n_6867),
.Y(n_10163)
);

AND2x2_ASAP7_75t_L g10164 ( 
.A(n_9481),
.B(n_7919),
.Y(n_10164)
);

A2O1A1Ixp33_ASAP7_75t_L g10165 ( 
.A1(n_9239),
.A2(n_7050),
.B(n_7100),
.C(n_7088),
.Y(n_10165)
);

OR2x6_ASAP7_75t_L g10166 ( 
.A(n_9481),
.B(n_8058),
.Y(n_10166)
);

OAI22xp5_ASAP7_75t_L g10167 ( 
.A1(n_9564),
.A2(n_7217),
.B1(n_7482),
.B2(n_6812),
.Y(n_10167)
);

AND2x4_ASAP7_75t_L g10168 ( 
.A(n_9287),
.B(n_8346),
.Y(n_10168)
);

AND2x2_ASAP7_75t_L g10169 ( 
.A(n_9553),
.B(n_9571),
.Y(n_10169)
);

AND2x2_ASAP7_75t_L g10170 ( 
.A(n_9553),
.B(n_7921),
.Y(n_10170)
);

OAI22xp5_ASAP7_75t_L g10171 ( 
.A1(n_9564),
.A2(n_7482),
.B1(n_6826),
.B2(n_6810),
.Y(n_10171)
);

OAI22xp5_ASAP7_75t_L g10172 ( 
.A1(n_9564),
.A2(n_6975),
.B1(n_7170),
.B2(n_7274),
.Y(n_10172)
);

INVxp67_ASAP7_75t_L g10173 ( 
.A(n_9450),
.Y(n_10173)
);

AND2x2_ASAP7_75t_L g10174 ( 
.A(n_9571),
.B(n_8945),
.Y(n_10174)
);

AOI22xp5_ASAP7_75t_L g10175 ( 
.A1(n_9042),
.A2(n_7476),
.B1(n_6929),
.B2(n_8393),
.Y(n_10175)
);

AND2x2_ASAP7_75t_L g10176 ( 
.A(n_8945),
.B(n_7921),
.Y(n_10176)
);

INVx2_ASAP7_75t_L g10177 ( 
.A(n_9450),
.Y(n_10177)
);

OR2x2_ASAP7_75t_L g10178 ( 
.A(n_9053),
.B(n_8562),
.Y(n_10178)
);

OAI21x1_ASAP7_75t_L g10179 ( 
.A1(n_8965),
.A2(n_9574),
.B(n_9386),
.Y(n_10179)
);

OA21x2_ASAP7_75t_L g10180 ( 
.A1(n_9693),
.A2(n_8097),
.B(n_8089),
.Y(n_10180)
);

INVx1_ASAP7_75t_L g10181 ( 
.A(n_8862),
.Y(n_10181)
);

A2O1A1Ixp33_ASAP7_75t_L g10182 ( 
.A1(n_9259),
.A2(n_9053),
.B(n_9688),
.C(n_8909),
.Y(n_10182)
);

OAI21x1_ASAP7_75t_SL g10183 ( 
.A1(n_9282),
.A2(n_6971),
.B(n_6960),
.Y(n_10183)
);

AND2x4_ASAP7_75t_L g10184 ( 
.A(n_9314),
.B(n_8407),
.Y(n_10184)
);

INVx4_ASAP7_75t_L g10185 ( 
.A(n_9259),
.Y(n_10185)
);

CKINVDCx5p33_ASAP7_75t_R g10186 ( 
.A(n_9276),
.Y(n_10186)
);

AND2x2_ASAP7_75t_L g10187 ( 
.A(n_8948),
.B(n_7921),
.Y(n_10187)
);

AND2x2_ASAP7_75t_L g10188 ( 
.A(n_8948),
.B(n_7921),
.Y(n_10188)
);

HB1xp67_ASAP7_75t_L g10189 ( 
.A(n_9404),
.Y(n_10189)
);

INVx1_ASAP7_75t_L g10190 ( 
.A(n_8862),
.Y(n_10190)
);

NAND2xp33_ASAP7_75t_L g10191 ( 
.A(n_9450),
.B(n_7809),
.Y(n_10191)
);

OA21x2_ASAP7_75t_L g10192 ( 
.A1(n_9574),
.A2(n_8109),
.B(n_8097),
.Y(n_10192)
);

NAND2xp5_ASAP7_75t_L g10193 ( 
.A(n_9314),
.B(n_6867),
.Y(n_10193)
);

NOR2xp33_ASAP7_75t_L g10194 ( 
.A(n_9628),
.B(n_6866),
.Y(n_10194)
);

OR2x2_ASAP7_75t_L g10195 ( 
.A(n_9288),
.B(n_8562),
.Y(n_10195)
);

NAND2xp5_ASAP7_75t_L g10196 ( 
.A(n_9339),
.B(n_8522),
.Y(n_10196)
);

OR2x2_ASAP7_75t_L g10197 ( 
.A(n_8820),
.B(n_8688),
.Y(n_10197)
);

AOI221xp5_ASAP7_75t_L g10198 ( 
.A1(n_9278),
.A2(n_8512),
.B1(n_8413),
.B2(n_8499),
.C(n_7023),
.Y(n_10198)
);

AND2x4_ASAP7_75t_L g10199 ( 
.A(n_9339),
.B(n_8407),
.Y(n_10199)
);

A2O1A1Ixp33_ASAP7_75t_L g10200 ( 
.A1(n_8864),
.A2(n_7050),
.B(n_7100),
.C(n_7088),
.Y(n_10200)
);

INVx2_ASAP7_75t_L g10201 ( 
.A(n_9450),
.Y(n_10201)
);

NAND2xp5_ASAP7_75t_L g10202 ( 
.A(n_9340),
.B(n_8522),
.Y(n_10202)
);

A2O1A1Ixp33_ASAP7_75t_L g10203 ( 
.A1(n_8864),
.A2(n_7100),
.B(n_8520),
.C(n_8517),
.Y(n_10203)
);

AOI221xp5_ASAP7_75t_L g10204 ( 
.A1(n_9278),
.A2(n_9393),
.B1(n_9297),
.B2(n_9601),
.C(n_9591),
.Y(n_10204)
);

OAI21xp5_ASAP7_75t_L g10205 ( 
.A1(n_9340),
.A2(n_8733),
.B(n_8722),
.Y(n_10205)
);

NAND2xp5_ASAP7_75t_L g10206 ( 
.A(n_9362),
.B(n_8522),
.Y(n_10206)
);

CKINVDCx20_ASAP7_75t_R g10207 ( 
.A(n_9676),
.Y(n_10207)
);

OAI21xp5_ASAP7_75t_L g10208 ( 
.A1(n_9362),
.A2(n_8753),
.B(n_8517),
.Y(n_10208)
);

INVx3_ASAP7_75t_L g10209 ( 
.A(n_8932),
.Y(n_10209)
);

NAND2xp5_ASAP7_75t_L g10210 ( 
.A(n_9412),
.B(n_9525),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_9450),
.Y(n_10211)
);

OR2x2_ASAP7_75t_L g10212 ( 
.A(n_8820),
.B(n_8688),
.Y(n_10212)
);

AO21x2_ASAP7_75t_L g10213 ( 
.A1(n_9393),
.A2(n_8199),
.B(n_8198),
.Y(n_10213)
);

AND2x2_ASAP7_75t_L g10214 ( 
.A(n_8953),
.B(n_8972),
.Y(n_10214)
);

OAI21xp5_ASAP7_75t_L g10215 ( 
.A1(n_9412),
.A2(n_8753),
.B(n_8517),
.Y(n_10215)
);

AOI221xp5_ASAP7_75t_L g10216 ( 
.A1(n_9297),
.A2(n_8512),
.B1(n_8413),
.B2(n_8499),
.C(n_7023),
.Y(n_10216)
);

OAI211xp5_ASAP7_75t_SL g10217 ( 
.A1(n_8856),
.A2(n_7076),
.B(n_7131),
.C(n_7119),
.Y(n_10217)
);

BUFx8_ASAP7_75t_SL g10218 ( 
.A(n_9474),
.Y(n_10218)
);

AND2x2_ASAP7_75t_L g10219 ( 
.A(n_8953),
.B(n_7921),
.Y(n_10219)
);

INVx4_ASAP7_75t_SL g10220 ( 
.A(n_9474),
.Y(n_10220)
);

A2O1A1Ixp33_ASAP7_75t_L g10221 ( 
.A1(n_8909),
.A2(n_8520),
.B(n_8485),
.C(n_8500),
.Y(n_10221)
);

AND2x2_ASAP7_75t_L g10222 ( 
.A(n_8972),
.B(n_7948),
.Y(n_10222)
);

OR2x2_ASAP7_75t_L g10223 ( 
.A(n_8854),
.B(n_8688),
.Y(n_10223)
);

AND2x4_ASAP7_75t_L g10224 ( 
.A(n_9525),
.B(n_8407),
.Y(n_10224)
);

AND2x2_ASAP7_75t_L g10225 ( 
.A(n_8981),
.B(n_7948),
.Y(n_10225)
);

OAI21xp5_ASAP7_75t_L g10226 ( 
.A1(n_9546),
.A2(n_8753),
.B(n_8520),
.Y(n_10226)
);

AND2x2_ASAP7_75t_L g10227 ( 
.A(n_8981),
.B(n_7948),
.Y(n_10227)
);

AOI22xp5_ASAP7_75t_L g10228 ( 
.A1(n_9042),
.A2(n_7476),
.B1(n_6929),
.B2(n_8393),
.Y(n_10228)
);

AND2x2_ASAP7_75t_L g10229 ( 
.A(n_8982),
.B(n_7948),
.Y(n_10229)
);

A2O1A1Ixp33_ASAP7_75t_L g10230 ( 
.A1(n_9676),
.A2(n_8485),
.B(n_8500),
.C(n_8477),
.Y(n_10230)
);

INVx2_ASAP7_75t_L g10231 ( 
.A(n_9474),
.Y(n_10231)
);

AND2x4_ASAP7_75t_L g10232 ( 
.A(n_9546),
.B(n_8407),
.Y(n_10232)
);

NAND2xp5_ASAP7_75t_L g10233 ( 
.A(n_9585),
.B(n_8525),
.Y(n_10233)
);

AOI22xp5_ASAP7_75t_L g10234 ( 
.A1(n_9009),
.A2(n_7352),
.B1(n_7328),
.B2(n_8058),
.Y(n_10234)
);

OAI211xp5_ASAP7_75t_L g10235 ( 
.A1(n_9685),
.A2(n_8261),
.B(n_8209),
.C(n_8216),
.Y(n_10235)
);

NOR2xp33_ASAP7_75t_L g10236 ( 
.A(n_9628),
.B(n_8886),
.Y(n_10236)
);

AOI21x1_ASAP7_75t_L g10237 ( 
.A1(n_8911),
.A2(n_8663),
.B(n_8627),
.Y(n_10237)
);

INVx2_ASAP7_75t_L g10238 ( 
.A(n_9474),
.Y(n_10238)
);

AND2x4_ASAP7_75t_L g10239 ( 
.A(n_9585),
.B(n_9657),
.Y(n_10239)
);

BUFx3_ASAP7_75t_L g10240 ( 
.A(n_9474),
.Y(n_10240)
);

AND2x2_ASAP7_75t_L g10241 ( 
.A(n_8982),
.B(n_7948),
.Y(n_10241)
);

BUFx12f_ASAP7_75t_L g10242 ( 
.A(n_9628),
.Y(n_10242)
);

INVx2_ASAP7_75t_L g10243 ( 
.A(n_9632),
.Y(n_10243)
);

AND2x6_ASAP7_75t_L g10244 ( 
.A(n_9632),
.B(n_7122),
.Y(n_10244)
);

OAI22xp5_ASAP7_75t_L g10245 ( 
.A1(n_9554),
.A2(n_7274),
.B1(n_6916),
.B2(n_6893),
.Y(n_10245)
);

AND2x2_ASAP7_75t_L g10246 ( 
.A(n_9003),
.B(n_7969),
.Y(n_10246)
);

INVx1_ASAP7_75t_L g10247 ( 
.A(n_8866),
.Y(n_10247)
);

NAND2xp5_ASAP7_75t_L g10248 ( 
.A(n_9657),
.B(n_8525),
.Y(n_10248)
);

AND2x4_ASAP7_75t_L g10249 ( 
.A(n_9658),
.B(n_8407),
.Y(n_10249)
);

NOR2x1_ASAP7_75t_SL g10250 ( 
.A(n_9009),
.B(n_8707),
.Y(n_10250)
);

BUFx3_ASAP7_75t_L g10251 ( 
.A(n_9632),
.Y(n_10251)
);

AO32x2_ASAP7_75t_L g10252 ( 
.A1(n_9658),
.A2(n_8017),
.A3(n_8063),
.B1(n_7987),
.B2(n_7955),
.Y(n_10252)
);

NAND2xp5_ASAP7_75t_L g10253 ( 
.A(n_9669),
.B(n_8525),
.Y(n_10253)
);

OA21x2_ASAP7_75t_L g10254 ( 
.A1(n_8965),
.A2(n_8116),
.B(n_8109),
.Y(n_10254)
);

AND2x4_ASAP7_75t_L g10255 ( 
.A(n_9669),
.B(n_8551),
.Y(n_10255)
);

NOR2xp33_ASAP7_75t_L g10256 ( 
.A(n_8886),
.B(n_6961),
.Y(n_10256)
);

OR2x2_ASAP7_75t_L g10257 ( 
.A(n_8854),
.B(n_8767),
.Y(n_10257)
);

NOR2xp33_ASAP7_75t_L g10258 ( 
.A(n_8886),
.B(n_6961),
.Y(n_10258)
);

NAND2xp5_ASAP7_75t_SL g10259 ( 
.A(n_9632),
.B(n_8324),
.Y(n_10259)
);

AOI221xp5_ASAP7_75t_L g10260 ( 
.A1(n_9297),
.A2(n_7916),
.B1(n_7022),
.B2(n_7014),
.C(n_7036),
.Y(n_10260)
);

OAI21x1_ASAP7_75t_L g10261 ( 
.A1(n_9376),
.A2(n_8706),
.B(n_7829),
.Y(n_10261)
);

OAI22xp33_ASAP7_75t_SL g10262 ( 
.A1(n_9182),
.A2(n_8252),
.B1(n_8063),
.B2(n_8095),
.Y(n_10262)
);

OAI21xp5_ASAP7_75t_L g10263 ( 
.A1(n_9493),
.A2(n_8500),
.B(n_8485),
.Y(n_10263)
);

OR2x2_ASAP7_75t_L g10264 ( 
.A(n_8995),
.B(n_9023),
.Y(n_10264)
);

AND2x4_ASAP7_75t_L g10265 ( 
.A(n_8852),
.B(n_8551),
.Y(n_10265)
);

AOI22xp33_ASAP7_75t_L g10266 ( 
.A1(n_9603),
.A2(n_8281),
.B1(n_7916),
.B2(n_7282),
.Y(n_10266)
);

A2O1A1Ixp33_ASAP7_75t_L g10267 ( 
.A1(n_9676),
.A2(n_9163),
.B(n_9074),
.C(n_9066),
.Y(n_10267)
);

AND2x2_ASAP7_75t_L g10268 ( 
.A(n_9003),
.B(n_7969),
.Y(n_10268)
);

A2O1A1Ixp33_ASAP7_75t_L g10269 ( 
.A1(n_9676),
.A2(n_8477),
.B(n_7122),
.C(n_7135),
.Y(n_10269)
);

HB1xp67_ASAP7_75t_L g10270 ( 
.A(n_9413),
.Y(n_10270)
);

OAI21xp5_ASAP7_75t_L g10271 ( 
.A1(n_9685),
.A2(n_8477),
.B(n_8261),
.Y(n_10271)
);

AND2x2_ASAP7_75t_L g10272 ( 
.A(n_9034),
.B(n_7969),
.Y(n_10272)
);

INVx4_ASAP7_75t_L g10273 ( 
.A(n_9632),
.Y(n_10273)
);

AND2x4_ASAP7_75t_L g10274 ( 
.A(n_8852),
.B(n_8551),
.Y(n_10274)
);

OAI21xp5_ASAP7_75t_L g10275 ( 
.A1(n_9685),
.A2(n_8261),
.B(n_8506),
.Y(n_10275)
);

INVx4_ASAP7_75t_L g10276 ( 
.A(n_9676),
.Y(n_10276)
);

NAND2xp5_ASAP7_75t_L g10277 ( 
.A(n_9086),
.B(n_9240),
.Y(n_10277)
);

INVx1_ASAP7_75t_L g10278 ( 
.A(n_8866),
.Y(n_10278)
);

OR2x6_ASAP7_75t_L g10279 ( 
.A(n_9554),
.B(n_8252),
.Y(n_10279)
);

A2O1A1Ixp33_ASAP7_75t_L g10280 ( 
.A1(n_9163),
.A2(n_7122),
.B(n_7135),
.C(n_8506),
.Y(n_10280)
);

AND2x2_ASAP7_75t_L g10281 ( 
.A(n_9034),
.B(n_7969),
.Y(n_10281)
);

NAND2xp5_ASAP7_75t_L g10282 ( 
.A(n_9086),
.B(n_8528),
.Y(n_10282)
);

NOR2xp33_ASAP7_75t_SL g10283 ( 
.A(n_9066),
.B(n_6822),
.Y(n_10283)
);

OR2x2_ASAP7_75t_L g10284 ( 
.A(n_8995),
.B(n_8767),
.Y(n_10284)
);

OR2x2_ASAP7_75t_L g10285 ( 
.A(n_9023),
.B(n_8767),
.Y(n_10285)
);

NOR2xp33_ASAP7_75t_L g10286 ( 
.A(n_9074),
.B(n_6961),
.Y(n_10286)
);

O2A1O1Ixp33_ASAP7_75t_L g10287 ( 
.A1(n_9561),
.A2(n_8063),
.B(n_8095),
.C(n_8017),
.Y(n_10287)
);

AOI221xp5_ASAP7_75t_L g10288 ( 
.A1(n_9591),
.A2(n_7916),
.B1(n_7022),
.B2(n_7014),
.C(n_7036),
.Y(n_10288)
);

OAI22xp5_ASAP7_75t_L g10289 ( 
.A1(n_9678),
.A2(n_6893),
.B1(n_7414),
.B2(n_8252),
.Y(n_10289)
);

AND2x2_ASAP7_75t_L g10290 ( 
.A(n_9059),
.B(n_7969),
.Y(n_10290)
);

NAND2xp5_ASAP7_75t_L g10291 ( 
.A(n_9086),
.B(n_8528),
.Y(n_10291)
);

NAND2xp5_ASAP7_75t_L g10292 ( 
.A(n_9086),
.B(n_8528),
.Y(n_10292)
);

OR2x2_ASAP7_75t_L g10293 ( 
.A(n_9344),
.B(n_6634),
.Y(n_10293)
);

OAI22xp5_ASAP7_75t_SL g10294 ( 
.A1(n_9678),
.A2(n_7095),
.B1(n_6989),
.B2(n_7056),
.Y(n_10294)
);

AND2x2_ASAP7_75t_L g10295 ( 
.A(n_9059),
.B(n_7988),
.Y(n_10295)
);

NOR2xp33_ASAP7_75t_L g10296 ( 
.A(n_9633),
.B(n_6965),
.Y(n_10296)
);

AO21x2_ASAP7_75t_L g10297 ( 
.A1(n_9222),
.A2(n_8200),
.B(n_8199),
.Y(n_10297)
);

INVx2_ASAP7_75t_L g10298 ( 
.A(n_8852),
.Y(n_10298)
);

OAI22xp5_ASAP7_75t_L g10299 ( 
.A1(n_9119),
.A2(n_7414),
.B1(n_8252),
.B2(n_7479),
.Y(n_10299)
);

AND2x4_ASAP7_75t_L g10300 ( 
.A(n_8878),
.B(n_8901),
.Y(n_10300)
);

AND2x2_ASAP7_75t_L g10301 ( 
.A(n_9061),
.B(n_7988),
.Y(n_10301)
);

INVx3_ASAP7_75t_L g10302 ( 
.A(n_8932),
.Y(n_10302)
);

INVxp67_ASAP7_75t_L g10303 ( 
.A(n_9584),
.Y(n_10303)
);

OAI21xp5_ASAP7_75t_L g10304 ( 
.A1(n_9685),
.A2(n_8261),
.B(n_8506),
.Y(n_10304)
);

OAI21xp5_ASAP7_75t_L g10305 ( 
.A1(n_9461),
.A2(n_8503),
.B(n_8216),
.Y(n_10305)
);

INVx1_ASAP7_75t_L g10306 ( 
.A(n_9691),
.Y(n_10306)
);

AOI221x1_ASAP7_75t_SL g10307 ( 
.A1(n_9427),
.A2(n_7039),
.B1(n_7065),
.B2(n_7201),
.C(n_7286),
.Y(n_10307)
);

AND2x2_ASAP7_75t_L g10308 ( 
.A(n_9061),
.B(n_7988),
.Y(n_10308)
);

AOI21xp5_ASAP7_75t_L g10309 ( 
.A1(n_9510),
.A2(n_7804),
.B(n_7810),
.Y(n_10309)
);

AND2x2_ASAP7_75t_L g10310 ( 
.A(n_9069),
.B(n_7988),
.Y(n_10310)
);

AND2x2_ASAP7_75t_L g10311 ( 
.A(n_9069),
.B(n_7988),
.Y(n_10311)
);

NAND2xp5_ASAP7_75t_L g10312 ( 
.A(n_9086),
.B(n_8541),
.Y(n_10312)
);

INVx1_ASAP7_75t_L g10313 ( 
.A(n_9686),
.Y(n_10313)
);

AND2x2_ASAP7_75t_L g10314 ( 
.A(n_9122),
.B(n_8004),
.Y(n_10314)
);

NOR2xp33_ASAP7_75t_L g10315 ( 
.A(n_9496),
.B(n_6965),
.Y(n_10315)
);

AND2x2_ASAP7_75t_L g10316 ( 
.A(n_9122),
.B(n_8004),
.Y(n_10316)
);

OAI21xp5_ASAP7_75t_L g10317 ( 
.A1(n_9461),
.A2(n_8503),
.B(n_8216),
.Y(n_10317)
);

OR2x2_ASAP7_75t_L g10318 ( 
.A(n_9375),
.B(n_5992),
.Y(n_10318)
);

AND2x4_ASAP7_75t_L g10319 ( 
.A(n_8878),
.B(n_8551),
.Y(n_10319)
);

AND2x4_ASAP7_75t_L g10320 ( 
.A(n_8878),
.B(n_8551),
.Y(n_10320)
);

AND2x2_ASAP7_75t_L g10321 ( 
.A(n_9155),
.B(n_9169),
.Y(n_10321)
);

AND2x4_ASAP7_75t_L g10322 ( 
.A(n_8901),
.B(n_8660),
.Y(n_10322)
);

OA21x2_ASAP7_75t_L g10323 ( 
.A1(n_9293),
.A2(n_8116),
.B(n_8109),
.Y(n_10323)
);

NOR4xp25_ASAP7_75t_SL g10324 ( 
.A(n_9022),
.B(n_7256),
.C(n_7281),
.D(n_7187),
.Y(n_10324)
);

AO32x2_ASAP7_75t_L g10325 ( 
.A1(n_8919),
.A2(n_8095),
.A3(n_8126),
.B1(n_8105),
.B2(n_8101),
.Y(n_10325)
);

AND2x4_ASAP7_75t_L g10326 ( 
.A(n_8901),
.B(n_8660),
.Y(n_10326)
);

OR2x2_ASAP7_75t_L g10327 ( 
.A(n_9381),
.B(n_5992),
.Y(n_10327)
);

AND2x6_ASAP7_75t_L g10328 ( 
.A(n_9446),
.B(n_7135),
.Y(n_10328)
);

NAND2xp33_ASAP7_75t_SL g10329 ( 
.A(n_8858),
.B(n_6683),
.Y(n_10329)
);

OAI21xp5_ASAP7_75t_L g10330 ( 
.A1(n_9469),
.A2(n_8503),
.B(n_9485),
.Y(n_10330)
);

OR2x2_ASAP7_75t_L g10331 ( 
.A(n_9116),
.B(n_5992),
.Y(n_10331)
);

A2O1A1Ixp33_ASAP7_75t_L g10332 ( 
.A1(n_9119),
.A2(n_8036),
.B(n_8046),
.C(n_7991),
.Y(n_10332)
);

BUFx2_ASAP7_75t_L g10333 ( 
.A(n_9269),
.Y(n_10333)
);

AND2x2_ASAP7_75t_L g10334 ( 
.A(n_9155),
.B(n_8004),
.Y(n_10334)
);

INVx2_ASAP7_75t_L g10335 ( 
.A(n_8919),
.Y(n_10335)
);

OAI21xp5_ASAP7_75t_L g10336 ( 
.A1(n_9469),
.A2(n_8216),
.B(n_8209),
.Y(n_10336)
);

INVx4_ASAP7_75t_L g10337 ( 
.A(n_8925),
.Y(n_10337)
);

INVx1_ASAP7_75t_L g10338 ( 
.A(n_9694),
.Y(n_10338)
);

AND2x2_ASAP7_75t_L g10339 ( 
.A(n_9169),
.B(n_8004),
.Y(n_10339)
);

AOI21xp5_ASAP7_75t_L g10340 ( 
.A1(n_8858),
.A2(n_8281),
.B(n_7916),
.Y(n_10340)
);

INVx1_ASAP7_75t_L g10341 ( 
.A(n_8879),
.Y(n_10341)
);

OAI21xp5_ASAP7_75t_L g10342 ( 
.A1(n_9485),
.A2(n_8216),
.B(n_8209),
.Y(n_10342)
);

OR2x2_ASAP7_75t_L g10343 ( 
.A(n_9563),
.B(n_6011),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_8925),
.Y(n_10344)
);

OAI21xp5_ASAP7_75t_L g10345 ( 
.A1(n_9516),
.A2(n_8209),
.B(n_8105),
.Y(n_10345)
);

AND2x2_ASAP7_75t_L g10346 ( 
.A(n_9170),
.B(n_8004),
.Y(n_10346)
);

AO32x1_ASAP7_75t_L g10347 ( 
.A1(n_8939),
.A2(n_8126),
.A3(n_8150),
.B1(n_8105),
.B2(n_8101),
.Y(n_10347)
);

A2O1A1Ixp33_ASAP7_75t_L g10348 ( 
.A1(n_9050),
.A2(n_9080),
.B(n_9111),
.C(n_9057),
.Y(n_10348)
);

OA21x2_ASAP7_75t_L g10349 ( 
.A1(n_9293),
.A2(n_8120),
.B(n_8116),
.Y(n_10349)
);

INVx5_ASAP7_75t_SL g10350 ( 
.A(n_9603),
.Y(n_10350)
);

O2A1O1Ixp33_ASAP7_75t_L g10351 ( 
.A1(n_9250),
.A2(n_8126),
.B(n_8150),
.C(n_8101),
.Y(n_10351)
);

AO32x2_ASAP7_75t_L g10352 ( 
.A1(n_8939),
.A2(n_8150),
.A3(n_8433),
.B1(n_8282),
.B2(n_8180),
.Y(n_10352)
);

OAI21xp5_ASAP7_75t_L g10353 ( 
.A1(n_9516),
.A2(n_8917),
.B(n_8911),
.Y(n_10353)
);

AND2x2_ASAP7_75t_L g10354 ( 
.A(n_9170),
.B(n_9198),
.Y(n_10354)
);

AND2x2_ASAP7_75t_L g10355 ( 
.A(n_9198),
.B(n_8021),
.Y(n_10355)
);

AND2x2_ASAP7_75t_L g10356 ( 
.A(n_9210),
.B(n_8021),
.Y(n_10356)
);

NOR2x1_ASAP7_75t_SL g10357 ( 
.A(n_9603),
.B(n_8707),
.Y(n_10357)
);

BUFx3_ASAP7_75t_L g10358 ( 
.A(n_9210),
.Y(n_10358)
);

AOI211xp5_ASAP7_75t_L g10359 ( 
.A1(n_9050),
.A2(n_7306),
.B(n_7307),
.C(n_6902),
.Y(n_10359)
);

AND2x2_ASAP7_75t_L g10360 ( 
.A(n_9431),
.B(n_8021),
.Y(n_10360)
);

AND2x2_ASAP7_75t_L g10361 ( 
.A(n_9431),
.B(n_8021),
.Y(n_10361)
);

NOR2x1_ASAP7_75t_SL g10362 ( 
.A(n_8917),
.B(n_8707),
.Y(n_10362)
);

INVx1_ASAP7_75t_L g10363 ( 
.A(n_8879),
.Y(n_10363)
);

OR2x2_ASAP7_75t_L g10364 ( 
.A(n_9563),
.B(n_6011),
.Y(n_10364)
);

AND2x2_ASAP7_75t_L g10365 ( 
.A(n_9443),
.B(n_8021),
.Y(n_10365)
);

INVxp67_ASAP7_75t_L g10366 ( 
.A(n_9604),
.Y(n_10366)
);

OR2x2_ASAP7_75t_L g10367 ( 
.A(n_9512),
.B(n_6011),
.Y(n_10367)
);

AND2x4_ASAP7_75t_L g10368 ( 
.A(n_9443),
.B(n_8660),
.Y(n_10368)
);

NAND2x1_ASAP7_75t_L g10369 ( 
.A(n_8954),
.B(n_7820),
.Y(n_10369)
);

NAND3xp33_ASAP7_75t_L g10370 ( 
.A(n_9648),
.B(n_8209),
.C(n_8368),
.Y(n_10370)
);

AND2x4_ASAP7_75t_L g10371 ( 
.A(n_9527),
.B(n_8660),
.Y(n_10371)
);

OAI22xp5_ASAP7_75t_L g10372 ( 
.A1(n_9057),
.A2(n_8252),
.B1(n_7479),
.B2(n_7454),
.Y(n_10372)
);

OR2x2_ASAP7_75t_L g10373 ( 
.A(n_9528),
.B(n_9080),
.Y(n_10373)
);

NAND2xp5_ASAP7_75t_L g10374 ( 
.A(n_9656),
.B(n_8541),
.Y(n_10374)
);

NAND2xp5_ASAP7_75t_L g10375 ( 
.A(n_9671),
.B(n_8541),
.Y(n_10375)
);

INVx2_ASAP7_75t_L g10376 ( 
.A(n_8988),
.Y(n_10376)
);

INVx2_ASAP7_75t_L g10377 ( 
.A(n_8988),
.Y(n_10377)
);

AOI21x1_ASAP7_75t_L g10378 ( 
.A1(n_9397),
.A2(n_8663),
.B(n_8627),
.Y(n_10378)
);

AOI221xp5_ASAP7_75t_L g10379 ( 
.A1(n_9591),
.A2(n_7916),
.B1(n_7899),
.B2(n_8281),
.C(n_7201),
.Y(n_10379)
);

CKINVDCx5p33_ASAP7_75t_R g10380 ( 
.A(n_9006),
.Y(n_10380)
);

INVx2_ASAP7_75t_L g10381 ( 
.A(n_9006),
.Y(n_10381)
);

NAND2xp5_ASAP7_75t_L g10382 ( 
.A(n_9543),
.B(n_8615),
.Y(n_10382)
);

INVx2_ASAP7_75t_L g10383 ( 
.A(n_9026),
.Y(n_10383)
);

AND2x2_ASAP7_75t_L g10384 ( 
.A(n_9527),
.B(n_8045),
.Y(n_10384)
);

OR2x2_ASAP7_75t_L g10385 ( 
.A(n_9111),
.B(n_6073),
.Y(n_10385)
);

AND2x2_ASAP7_75t_L g10386 ( 
.A(n_9537),
.B(n_8045),
.Y(n_10386)
);

A2O1A1Ixp33_ASAP7_75t_L g10387 ( 
.A1(n_9376),
.A2(n_8036),
.B(n_8046),
.C(n_7991),
.Y(n_10387)
);

NAND2xp5_ASAP7_75t_L g10388 ( 
.A(n_9543),
.B(n_8615),
.Y(n_10388)
);

HB1xp67_ASAP7_75t_L g10389 ( 
.A(n_9022),
.Y(n_10389)
);

NAND2xp5_ASAP7_75t_L g10390 ( 
.A(n_9543),
.B(n_8615),
.Y(n_10390)
);

AO21x2_ASAP7_75t_L g10391 ( 
.A1(n_9222),
.A2(n_8211),
.B(n_8200),
.Y(n_10391)
);

AND2x2_ASAP7_75t_L g10392 ( 
.A(n_9537),
.B(n_8045),
.Y(n_10392)
);

A2O1A1Ixp33_ASAP7_75t_L g10393 ( 
.A1(n_9386),
.A2(n_8036),
.B(n_8046),
.C(n_7991),
.Y(n_10393)
);

A2O1A1Ixp33_ASAP7_75t_L g10394 ( 
.A1(n_8993),
.A2(n_8090),
.B(n_8091),
.C(n_8081),
.Y(n_10394)
);

INVx1_ASAP7_75t_L g10395 ( 
.A(n_8880),
.Y(n_10395)
);

INVx2_ASAP7_75t_L g10396 ( 
.A(n_9026),
.Y(n_10396)
);

OR2x2_ASAP7_75t_L g10397 ( 
.A(n_9583),
.B(n_6073),
.Y(n_10397)
);

NOR2x1_ASAP7_75t_SL g10398 ( 
.A(n_9206),
.B(n_7277),
.Y(n_10398)
);

AND2x2_ASAP7_75t_L g10399 ( 
.A(n_9562),
.B(n_8045),
.Y(n_10399)
);

AOI21xp5_ASAP7_75t_L g10400 ( 
.A1(n_9601),
.A2(n_8281),
.B(n_7917),
.Y(n_10400)
);

A2O1A1Ixp33_ASAP7_75t_L g10401 ( 
.A1(n_8993),
.A2(n_8090),
.B(n_8091),
.C(n_8081),
.Y(n_10401)
);

NAND2xp5_ASAP7_75t_L g10402 ( 
.A(n_9543),
.B(n_8619),
.Y(n_10402)
);

BUFx2_ASAP7_75t_L g10403 ( 
.A(n_9269),
.Y(n_10403)
);

OR2x2_ASAP7_75t_L g10404 ( 
.A(n_9583),
.B(n_6073),
.Y(n_10404)
);

AND2x2_ASAP7_75t_L g10405 ( 
.A(n_9562),
.B(n_8045),
.Y(n_10405)
);

OR2x2_ASAP7_75t_L g10406 ( 
.A(n_9605),
.B(n_6505),
.Y(n_10406)
);

INVx1_ASAP7_75t_L g10407 ( 
.A(n_8880),
.Y(n_10407)
);

AO21x2_ASAP7_75t_L g10408 ( 
.A1(n_9222),
.A2(n_8211),
.B(n_8200),
.Y(n_10408)
);

AND2x2_ASAP7_75t_L g10409 ( 
.A(n_9582),
.B(n_8057),
.Y(n_10409)
);

OA21x2_ASAP7_75t_L g10410 ( 
.A1(n_9347),
.A2(n_8123),
.B(n_8120),
.Y(n_10410)
);

AND2x2_ASAP7_75t_L g10411 ( 
.A(n_9582),
.B(n_8057),
.Y(n_10411)
);

INVx1_ASAP7_75t_L g10412 ( 
.A(n_8884),
.Y(n_10412)
);

AND2x2_ASAP7_75t_L g10413 ( 
.A(n_9615),
.B(n_8057),
.Y(n_10413)
);

AND2x2_ASAP7_75t_L g10414 ( 
.A(n_9615),
.B(n_8057),
.Y(n_10414)
);

OAI22xp5_ASAP7_75t_L g10415 ( 
.A1(n_9015),
.A2(n_7454),
.B1(n_7734),
.B2(n_7693),
.Y(n_10415)
);

AOI22xp5_ASAP7_75t_L g10416 ( 
.A1(n_9213),
.A2(n_7352),
.B1(n_7917),
.B2(n_7796),
.Y(n_10416)
);

NAND2xp5_ASAP7_75t_L g10417 ( 
.A(n_9543),
.B(n_8619),
.Y(n_10417)
);

AND2x2_ASAP7_75t_L g10418 ( 
.A(n_9617),
.B(n_8057),
.Y(n_10418)
);

OA21x2_ASAP7_75t_L g10419 ( 
.A1(n_9347),
.A2(n_8123),
.B(n_8120),
.Y(n_10419)
);

OAI22xp5_ASAP7_75t_L g10420 ( 
.A1(n_9015),
.A2(n_7734),
.B1(n_7693),
.B2(n_7156),
.Y(n_10420)
);

AO32x1_ASAP7_75t_L g10421 ( 
.A1(n_9024),
.A2(n_8433),
.A3(n_8450),
.B1(n_8282),
.B2(n_8180),
.Y(n_10421)
);

OR2x2_ASAP7_75t_L g10422 ( 
.A(n_9605),
.B(n_9487),
.Y(n_10422)
);

AO21x2_ASAP7_75t_L g10423 ( 
.A1(n_9250),
.A2(n_8218),
.B(n_8211),
.Y(n_10423)
);

OAI22xp5_ASAP7_75t_L g10424 ( 
.A1(n_9016),
.A2(n_7156),
.B1(n_7917),
.B2(n_7796),
.Y(n_10424)
);

A2O1A1Ixp33_ASAP7_75t_L g10425 ( 
.A1(n_9029),
.A2(n_8090),
.B(n_8091),
.C(n_8081),
.Y(n_10425)
);

A2O1A1Ixp33_ASAP7_75t_L g10426 ( 
.A1(n_9029),
.A2(n_8167),
.B(n_8206),
.C(n_8148),
.Y(n_10426)
);

NAND2xp5_ASAP7_75t_L g10427 ( 
.A(n_9487),
.B(n_8619),
.Y(n_10427)
);

OAI22xp5_ASAP7_75t_L g10428 ( 
.A1(n_9016),
.A2(n_7917),
.B1(n_7796),
.B2(n_7589),
.Y(n_10428)
);

OAI21xp5_ASAP7_75t_L g10429 ( 
.A1(n_9397),
.A2(n_8282),
.B(n_8180),
.Y(n_10429)
);

OAI211xp5_ASAP7_75t_L g10430 ( 
.A1(n_9502),
.A2(n_8368),
.B(n_8312),
.C(n_7951),
.Y(n_10430)
);

AND2x2_ASAP7_75t_L g10431 ( 
.A(n_9617),
.B(n_8107),
.Y(n_10431)
);

OAI211xp5_ASAP7_75t_L g10432 ( 
.A1(n_9502),
.A2(n_8368),
.B(n_9652),
.C(n_9624),
.Y(n_10432)
);

AOI21xp5_ASAP7_75t_L g10433 ( 
.A1(n_9601),
.A2(n_8281),
.B(n_7917),
.Y(n_10433)
);

AND2x2_ASAP7_75t_L g10434 ( 
.A(n_9630),
.B(n_8107),
.Y(n_10434)
);

OA21x2_ASAP7_75t_L g10435 ( 
.A1(n_9144),
.A2(n_9209),
.B(n_9129),
.Y(n_10435)
);

A2O1A1Ixp33_ASAP7_75t_L g10436 ( 
.A1(n_9129),
.A2(n_8167),
.B(n_8206),
.C(n_8148),
.Y(n_10436)
);

INVx1_ASAP7_75t_L g10437 ( 
.A(n_8884),
.Y(n_10437)
);

NAND2xp5_ASAP7_75t_SL g10438 ( 
.A(n_8954),
.B(n_8324),
.Y(n_10438)
);

NOR2xp33_ASAP7_75t_L g10439 ( 
.A(n_9539),
.B(n_6965),
.Y(n_10439)
);

AOI221xp5_ASAP7_75t_L g10440 ( 
.A1(n_9250),
.A2(n_7899),
.B1(n_7039),
.B2(n_7189),
.C(n_8103),
.Y(n_10440)
);

INVx1_ASAP7_75t_L g10441 ( 
.A(n_8885),
.Y(n_10441)
);

NAND2xp5_ASAP7_75t_L g10442 ( 
.A(n_9539),
.B(n_8628),
.Y(n_10442)
);

INVx2_ASAP7_75t_L g10443 ( 
.A(n_9446),
.Y(n_10443)
);

NAND2xp5_ASAP7_75t_L g10444 ( 
.A(n_9550),
.B(n_8628),
.Y(n_10444)
);

AND2x2_ASAP7_75t_L g10445 ( 
.A(n_9704),
.B(n_9630),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_9718),
.B(n_9631),
.Y(n_10446)
);

HB1xp67_ASAP7_75t_L g10447 ( 
.A(n_9777),
.Y(n_10447)
);

INVx2_ASAP7_75t_L g10448 ( 
.A(n_9830),
.Y(n_10448)
);

AND2x2_ASAP7_75t_L g10449 ( 
.A(n_9703),
.B(n_9631),
.Y(n_10449)
);

OR2x2_ASAP7_75t_L g10450 ( 
.A(n_9714),
.B(n_9550),
.Y(n_10450)
);

INVx3_ASAP7_75t_L g10451 ( 
.A(n_9773),
.Y(n_10451)
);

HB1xp67_ASAP7_75t_L g10452 ( 
.A(n_9784),
.Y(n_10452)
);

NAND2xp5_ASAP7_75t_L g10453 ( 
.A(n_9707),
.B(n_9024),
.Y(n_10453)
);

INVx2_ASAP7_75t_L g10454 ( 
.A(n_9831),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_9813),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_9860),
.Y(n_10456)
);

BUFx6f_ASAP7_75t_L g10457 ( 
.A(n_9812),
.Y(n_10457)
);

NAND2xp5_ASAP7_75t_L g10458 ( 
.A(n_9698),
.B(n_9025),
.Y(n_10458)
);

INVx1_ASAP7_75t_L g10459 ( 
.A(n_9892),
.Y(n_10459)
);

OAI21x1_ASAP7_75t_SL g10460 ( 
.A1(n_9785),
.A2(n_6971),
.B(n_6960),
.Y(n_10460)
);

AOI21x1_ASAP7_75t_L g10461 ( 
.A1(n_10118),
.A2(n_9031),
.B(n_9025),
.Y(n_10461)
);

INVx2_ASAP7_75t_L g10462 ( 
.A(n_9946),
.Y(n_10462)
);

INVx5_ASAP7_75t_L g10463 ( 
.A(n_9737),
.Y(n_10463)
);

INVx1_ASAP7_75t_L g10464 ( 
.A(n_9904),
.Y(n_10464)
);

AND2x4_ASAP7_75t_L g10465 ( 
.A(n_9882),
.B(n_8954),
.Y(n_10465)
);

AND2x2_ASAP7_75t_L g10466 ( 
.A(n_9769),
.B(n_9637),
.Y(n_10466)
);

AOI22xp33_ASAP7_75t_L g10467 ( 
.A1(n_9764),
.A2(n_9618),
.B1(n_9213),
.B2(n_9175),
.Y(n_10467)
);

NAND2xp5_ASAP7_75t_L g10468 ( 
.A(n_9711),
.B(n_9031),
.Y(n_10468)
);

OR2x2_ASAP7_75t_L g10469 ( 
.A(n_9726),
.B(n_8926),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_9699),
.Y(n_10470)
);

INVx1_ASAP7_75t_L g10471 ( 
.A(n_9699),
.Y(n_10471)
);

NOR2xp33_ASAP7_75t_L g10472 ( 
.A(n_9965),
.B(n_6986),
.Y(n_10472)
);

INVx2_ASAP7_75t_L g10473 ( 
.A(n_9950),
.Y(n_10473)
);

AND2x4_ASAP7_75t_L g10474 ( 
.A(n_9773),
.B(n_8978),
.Y(n_10474)
);

INVx1_ASAP7_75t_L g10475 ( 
.A(n_9722),
.Y(n_10475)
);

NAND2xp5_ASAP7_75t_L g10476 ( 
.A(n_9754),
.B(n_9032),
.Y(n_10476)
);

INVx2_ASAP7_75t_L g10477 ( 
.A(n_9838),
.Y(n_10477)
);

INVx2_ASAP7_75t_L g10478 ( 
.A(n_9838),
.Y(n_10478)
);

INVx2_ASAP7_75t_L g10479 ( 
.A(n_10127),
.Y(n_10479)
);

INVx1_ASAP7_75t_L g10480 ( 
.A(n_9722),
.Y(n_10480)
);

BUFx2_ASAP7_75t_L g10481 ( 
.A(n_9981),
.Y(n_10481)
);

INVx2_ASAP7_75t_L g10482 ( 
.A(n_10127),
.Y(n_10482)
);

AND2x2_ASAP7_75t_L g10483 ( 
.A(n_9751),
.B(n_9637),
.Y(n_10483)
);

INVx2_ASAP7_75t_L g10484 ( 
.A(n_10127),
.Y(n_10484)
);

AND2x2_ASAP7_75t_L g10485 ( 
.A(n_9753),
.B(n_9645),
.Y(n_10485)
);

NAND2xp5_ASAP7_75t_L g10486 ( 
.A(n_9723),
.B(n_9032),
.Y(n_10486)
);

INVx2_ASAP7_75t_L g10487 ( 
.A(n_10155),
.Y(n_10487)
);

BUFx2_ASAP7_75t_L g10488 ( 
.A(n_9981),
.Y(n_10488)
);

HB1xp67_ASAP7_75t_L g10489 ( 
.A(n_9952),
.Y(n_10489)
);

INVx1_ASAP7_75t_L g10490 ( 
.A(n_9724),
.Y(n_10490)
);

INVxp67_ASAP7_75t_L g10491 ( 
.A(n_9774),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_9724),
.Y(n_10492)
);

INVxp67_ASAP7_75t_SL g10493 ( 
.A(n_9785),
.Y(n_10493)
);

INVx2_ASAP7_75t_L g10494 ( 
.A(n_10155),
.Y(n_10494)
);

INVx2_ASAP7_75t_SL g10495 ( 
.A(n_9976),
.Y(n_10495)
);

NOR2x1_ASAP7_75t_SL g10496 ( 
.A(n_9752),
.B(n_7095),
.Y(n_10496)
);

OAI22xp5_ASAP7_75t_L g10497 ( 
.A1(n_9810),
.A2(n_7259),
.B1(n_7917),
.B2(n_7796),
.Y(n_10497)
);

BUFx3_ASAP7_75t_L g10498 ( 
.A(n_9826),
.Y(n_10498)
);

AO21x2_ASAP7_75t_L g10499 ( 
.A1(n_10062),
.A2(n_9036),
.B(n_9033),
.Y(n_10499)
);

INVx2_ASAP7_75t_L g10500 ( 
.A(n_10155),
.Y(n_10500)
);

AND2x2_ASAP7_75t_L g10501 ( 
.A(n_9733),
.B(n_9645),
.Y(n_10501)
);

NAND2xp5_ASAP7_75t_L g10502 ( 
.A(n_10027),
.B(n_9033),
.Y(n_10502)
);

NAND2xp5_ASAP7_75t_L g10503 ( 
.A(n_10050),
.B(n_9036),
.Y(n_10503)
);

INVx2_ASAP7_75t_L g10504 ( 
.A(n_10093),
.Y(n_10504)
);

INVx4_ASAP7_75t_L g10505 ( 
.A(n_10143),
.Y(n_10505)
);

HB1xp67_ASAP7_75t_L g10506 ( 
.A(n_10097),
.Y(n_10506)
);

INVx2_ASAP7_75t_L g10507 ( 
.A(n_10093),
.Y(n_10507)
);

AND2x2_ASAP7_75t_L g10508 ( 
.A(n_9771),
.B(n_9655),
.Y(n_10508)
);

AND2x2_ASAP7_75t_L g10509 ( 
.A(n_9780),
.B(n_9655),
.Y(n_10509)
);

NAND2xp5_ASAP7_75t_L g10510 ( 
.A(n_10099),
.B(n_9038),
.Y(n_10510)
);

AND2x2_ASAP7_75t_L g10511 ( 
.A(n_9720),
.B(n_9660),
.Y(n_10511)
);

AND2x2_ASAP7_75t_L g10512 ( 
.A(n_9725),
.B(n_9660),
.Y(n_10512)
);

INVx2_ASAP7_75t_L g10513 ( 
.A(n_10093),
.Y(n_10513)
);

AND2x2_ASAP7_75t_L g10514 ( 
.A(n_9731),
.B(n_9662),
.Y(n_10514)
);

AOI22xp33_ASAP7_75t_L g10515 ( 
.A1(n_9739),
.A2(n_9618),
.B1(n_9213),
.B2(n_9175),
.Y(n_10515)
);

INVx1_ASAP7_75t_L g10516 ( 
.A(n_9732),
.Y(n_10516)
);

AND2x2_ASAP7_75t_L g10517 ( 
.A(n_9888),
.B(n_9662),
.Y(n_10517)
);

INVx1_ASAP7_75t_L g10518 ( 
.A(n_9732),
.Y(n_10518)
);

INVx1_ASAP7_75t_L g10519 ( 
.A(n_9791),
.Y(n_10519)
);

AOI33xp33_ASAP7_75t_L g10520 ( 
.A1(n_10053),
.A2(n_7259),
.A3(n_9038),
.B1(n_9046),
.B2(n_9045),
.B3(n_9040),
.Y(n_10520)
);

INVx1_ASAP7_75t_L g10521 ( 
.A(n_9791),
.Y(n_10521)
);

HB1xp67_ASAP7_75t_L g10522 ( 
.A(n_10103),
.Y(n_10522)
);

AND2x2_ASAP7_75t_L g10523 ( 
.A(n_9999),
.B(n_9668),
.Y(n_10523)
);

AND2x2_ASAP7_75t_L g10524 ( 
.A(n_10000),
.B(n_10174),
.Y(n_10524)
);

AND2x2_ASAP7_75t_L g10525 ( 
.A(n_10135),
.B(n_9668),
.Y(n_10525)
);

INVx2_ASAP7_75t_L g10526 ( 
.A(n_10252),
.Y(n_10526)
);

INVx4_ASAP7_75t_R g10527 ( 
.A(n_9760),
.Y(n_10527)
);

AND2x2_ASAP7_75t_L g10528 ( 
.A(n_10136),
.B(n_8107),
.Y(n_10528)
);

BUFx2_ASAP7_75t_L g10529 ( 
.A(n_10218),
.Y(n_10529)
);

HB1xp67_ASAP7_75t_L g10530 ( 
.A(n_10189),
.Y(n_10530)
);

NAND2xp5_ASAP7_75t_L g10531 ( 
.A(n_10270),
.B(n_9040),
.Y(n_10531)
);

AND2x4_ASAP7_75t_SL g10532 ( 
.A(n_9752),
.B(n_6677),
.Y(n_10532)
);

OR2x2_ASAP7_75t_L g10533 ( 
.A(n_9709),
.B(n_8926),
.Y(n_10533)
);

INVx3_ASAP7_75t_L g10534 ( 
.A(n_10300),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_9859),
.Y(n_10535)
);

BUFx6f_ASAP7_75t_L g10536 ( 
.A(n_10020),
.Y(n_10536)
);

NAND2xp5_ASAP7_75t_L g10537 ( 
.A(n_10307),
.B(n_9045),
.Y(n_10537)
);

OR2x2_ASAP7_75t_L g10538 ( 
.A(n_10373),
.B(n_8955),
.Y(n_10538)
);

AND2x2_ASAP7_75t_L g10539 ( 
.A(n_10169),
.B(n_8107),
.Y(n_10539)
);

INVx1_ASAP7_75t_L g10540 ( 
.A(n_9859),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9880),
.Y(n_10541)
);

INVx3_ASAP7_75t_L g10542 ( 
.A(n_10300),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_9880),
.Y(n_10543)
);

INVx2_ASAP7_75t_L g10544 ( 
.A(n_10252),
.Y(n_10544)
);

HB1xp67_ASAP7_75t_L g10545 ( 
.A(n_9856),
.Y(n_10545)
);

AND2x2_ASAP7_75t_L g10546 ( 
.A(n_9789),
.B(n_8107),
.Y(n_10546)
);

INVx1_ASAP7_75t_L g10547 ( 
.A(n_9881),
.Y(n_10547)
);

INVx2_ASAP7_75t_SL g10548 ( 
.A(n_9976),
.Y(n_10548)
);

INVx1_ASAP7_75t_L g10549 ( 
.A(n_9881),
.Y(n_10549)
);

INVx1_ASAP7_75t_L g10550 ( 
.A(n_9908),
.Y(n_10550)
);

AND2x2_ASAP7_75t_SL g10551 ( 
.A(n_9918),
.B(n_6971),
.Y(n_10551)
);

NAND2xp5_ASAP7_75t_L g10552 ( 
.A(n_9861),
.B(n_9046),
.Y(n_10552)
);

AND2x2_ASAP7_75t_L g10553 ( 
.A(n_9790),
.B(n_8113),
.Y(n_10553)
);

INVx2_ASAP7_75t_L g10554 ( 
.A(n_10252),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_9792),
.B(n_8113),
.Y(n_10555)
);

NOR2xp67_ASAP7_75t_L g10556 ( 
.A(n_9990),
.B(n_8978),
.Y(n_10556)
);

INVx2_ASAP7_75t_L g10557 ( 
.A(n_10220),
.Y(n_10557)
);

HB1xp67_ASAP7_75t_L g10558 ( 
.A(n_9900),
.Y(n_10558)
);

NAND2xp5_ASAP7_75t_L g10559 ( 
.A(n_10303),
.B(n_9047),
.Y(n_10559)
);

OR2x2_ASAP7_75t_L g10560 ( 
.A(n_9804),
.B(n_8955),
.Y(n_10560)
);

AND2x2_ASAP7_75t_L g10561 ( 
.A(n_9806),
.B(n_8113),
.Y(n_10561)
);

OR2x2_ASAP7_75t_L g10562 ( 
.A(n_10264),
.B(n_9334),
.Y(n_10562)
);

INVx1_ASAP7_75t_L g10563 ( 
.A(n_9908),
.Y(n_10563)
);

HB1xp67_ASAP7_75t_L g10564 ( 
.A(n_10333),
.Y(n_10564)
);

AND2x4_ASAP7_75t_L g10565 ( 
.A(n_10220),
.B(n_8978),
.Y(n_10565)
);

NAND2xp5_ASAP7_75t_L g10566 ( 
.A(n_9734),
.B(n_9047),
.Y(n_10566)
);

NAND2xp5_ASAP7_75t_L g10567 ( 
.A(n_9700),
.B(n_9048),
.Y(n_10567)
);

AOI22xp33_ASAP7_75t_L g10568 ( 
.A1(n_9801),
.A2(n_9618),
.B1(n_9175),
.B2(n_8103),
.Y(n_10568)
);

AND2x2_ASAP7_75t_L g10569 ( 
.A(n_9815),
.B(n_8113),
.Y(n_10569)
);

INVx2_ASAP7_75t_L g10570 ( 
.A(n_10265),
.Y(n_10570)
);

NAND2xp5_ASAP7_75t_SL g10571 ( 
.A(n_9961),
.B(n_6691),
.Y(n_10571)
);

INVx1_ASAP7_75t_L g10572 ( 
.A(n_9910),
.Y(n_10572)
);

BUFx3_ASAP7_75t_L g10573 ( 
.A(n_9824),
.Y(n_10573)
);

AND2x2_ASAP7_75t_L g10574 ( 
.A(n_9819),
.B(n_8113),
.Y(n_10574)
);

AND2x2_ASAP7_75t_L g10575 ( 
.A(n_9825),
.B(n_8117),
.Y(n_10575)
);

INVx2_ASAP7_75t_L g10576 ( 
.A(n_10265),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_9910),
.Y(n_10577)
);

AND2x4_ASAP7_75t_L g10578 ( 
.A(n_10273),
.B(n_9097),
.Y(n_10578)
);

BUFx2_ASAP7_75t_L g10579 ( 
.A(n_10242),
.Y(n_10579)
);

CKINVDCx11_ASAP7_75t_R g10580 ( 
.A(n_10114),
.Y(n_10580)
);

BUFx6f_ASAP7_75t_L g10581 ( 
.A(n_9770),
.Y(n_10581)
);

AND2x4_ASAP7_75t_L g10582 ( 
.A(n_10273),
.B(n_9097),
.Y(n_10582)
);

HB1xp67_ASAP7_75t_L g10583 ( 
.A(n_10403),
.Y(n_10583)
);

AND2x2_ASAP7_75t_L g10584 ( 
.A(n_9828),
.B(n_8117),
.Y(n_10584)
);

INVx1_ASAP7_75t_SL g10585 ( 
.A(n_10028),
.Y(n_10585)
);

HB1xp67_ASAP7_75t_L g10586 ( 
.A(n_9729),
.Y(n_10586)
);

HB1xp67_ASAP7_75t_L g10587 ( 
.A(n_10389),
.Y(n_10587)
);

OR2x2_ASAP7_75t_L g10588 ( 
.A(n_9891),
.B(n_9334),
.Y(n_10588)
);

BUFx6f_ASAP7_75t_L g10589 ( 
.A(n_9770),
.Y(n_10589)
);

AND2x2_ASAP7_75t_L g10590 ( 
.A(n_9740),
.B(n_8117),
.Y(n_10590)
);

INVx2_ASAP7_75t_L g10591 ( 
.A(n_10325),
.Y(n_10591)
);

INVx1_ASAP7_75t_L g10592 ( 
.A(n_9940),
.Y(n_10592)
);

AND2x2_ASAP7_75t_L g10593 ( 
.A(n_9746),
.B(n_9955),
.Y(n_10593)
);

AND2x2_ASAP7_75t_L g10594 ( 
.A(n_9972),
.B(n_8117),
.Y(n_10594)
);

BUFx2_ASAP7_75t_L g10595 ( 
.A(n_9983),
.Y(n_10595)
);

NOR2x1_ASAP7_75t_SL g10596 ( 
.A(n_10279),
.B(n_7095),
.Y(n_10596)
);

INVx2_ASAP7_75t_L g10597 ( 
.A(n_10325),
.Y(n_10597)
);

CKINVDCx5p33_ASAP7_75t_R g10598 ( 
.A(n_9887),
.Y(n_10598)
);

INVxp67_ASAP7_75t_SL g10599 ( 
.A(n_9970),
.Y(n_10599)
);

NAND2xp5_ASAP7_75t_L g10600 ( 
.A(n_9702),
.B(n_9048),
.Y(n_10600)
);

NOR2xp33_ASAP7_75t_L g10601 ( 
.A(n_9965),
.B(n_9990),
.Y(n_10601)
);

INVx2_ASAP7_75t_L g10602 ( 
.A(n_10325),
.Y(n_10602)
);

HB1xp67_ASAP7_75t_L g10603 ( 
.A(n_9728),
.Y(n_10603)
);

INVx3_ASAP7_75t_L g10604 ( 
.A(n_10274),
.Y(n_10604)
);

AND2x2_ASAP7_75t_L g10605 ( 
.A(n_9974),
.B(n_8117),
.Y(n_10605)
);

INVx1_ASAP7_75t_SL g10606 ( 
.A(n_10142),
.Y(n_10606)
);

BUFx2_ASAP7_75t_L g10607 ( 
.A(n_9758),
.Y(n_10607)
);

AND2x2_ASAP7_75t_L g10608 ( 
.A(n_9836),
.B(n_8162),
.Y(n_10608)
);

AND2x2_ASAP7_75t_L g10609 ( 
.A(n_9852),
.B(n_8162),
.Y(n_10609)
);

INVx1_ASAP7_75t_L g10610 ( 
.A(n_9940),
.Y(n_10610)
);

INVx1_ASAP7_75t_L g10611 ( 
.A(n_9942),
.Y(n_10611)
);

AND2x2_ASAP7_75t_L g10612 ( 
.A(n_9857),
.B(n_8162),
.Y(n_10612)
);

AND2x2_ASAP7_75t_L g10613 ( 
.A(n_9863),
.B(n_8162),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_9942),
.Y(n_10614)
);

INVx5_ASAP7_75t_L g10615 ( 
.A(n_9737),
.Y(n_10615)
);

AND2x2_ASAP7_75t_L g10616 ( 
.A(n_9865),
.B(n_8162),
.Y(n_10616)
);

INVx2_ASAP7_75t_L g10617 ( 
.A(n_10352),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_9995),
.Y(n_10618)
);

AND2x2_ASAP7_75t_L g10619 ( 
.A(n_9866),
.B(n_8173),
.Y(n_10619)
);

INVx1_ASAP7_75t_L g10620 ( 
.A(n_9995),
.Y(n_10620)
);

AND2x2_ASAP7_75t_L g10621 ( 
.A(n_9870),
.B(n_8173),
.Y(n_10621)
);

INVx2_ASAP7_75t_L g10622 ( 
.A(n_10274),
.Y(n_10622)
);

INVx4_ASAP7_75t_L g10623 ( 
.A(n_9822),
.Y(n_10623)
);

INVx1_ASAP7_75t_L g10624 ( 
.A(n_10004),
.Y(n_10624)
);

AND2x2_ASAP7_75t_L g10625 ( 
.A(n_9871),
.B(n_9874),
.Y(n_10625)
);

INVx2_ASAP7_75t_L g10626 ( 
.A(n_10319),
.Y(n_10626)
);

INVx2_ASAP7_75t_L g10627 ( 
.A(n_10319),
.Y(n_10627)
);

OR2x2_ASAP7_75t_L g10628 ( 
.A(n_9939),
.B(n_9301),
.Y(n_10628)
);

INVx1_ASAP7_75t_L g10629 ( 
.A(n_10004),
.Y(n_10629)
);

INVx1_ASAP7_75t_L g10630 ( 
.A(n_10019),
.Y(n_10630)
);

BUFx6f_ASAP7_75t_L g10631 ( 
.A(n_9770),
.Y(n_10631)
);

NAND2xp5_ASAP7_75t_L g10632 ( 
.A(n_9744),
.B(n_9054),
.Y(n_10632)
);

AND2x2_ASAP7_75t_L g10633 ( 
.A(n_9878),
.B(n_8173),
.Y(n_10633)
);

AND2x4_ASAP7_75t_L g10634 ( 
.A(n_10239),
.B(n_9097),
.Y(n_10634)
);

BUFx6f_ASAP7_75t_L g10635 ( 
.A(n_9798),
.Y(n_10635)
);

INVx2_ASAP7_75t_L g10636 ( 
.A(n_10320),
.Y(n_10636)
);

INVx2_ASAP7_75t_L g10637 ( 
.A(n_10320),
.Y(n_10637)
);

INVx2_ASAP7_75t_L g10638 ( 
.A(n_10322),
.Y(n_10638)
);

AND2x2_ASAP7_75t_L g10639 ( 
.A(n_9894),
.B(n_8173),
.Y(n_10639)
);

AND2x4_ASAP7_75t_L g10640 ( 
.A(n_10239),
.B(n_9183),
.Y(n_10640)
);

AND2x4_ASAP7_75t_L g10641 ( 
.A(n_9846),
.B(n_9183),
.Y(n_10641)
);

AND2x2_ASAP7_75t_L g10642 ( 
.A(n_9898),
.B(n_9986),
.Y(n_10642)
);

INVx1_ASAP7_75t_L g10643 ( 
.A(n_10019),
.Y(n_10643)
);

INVx2_ASAP7_75t_L g10644 ( 
.A(n_10322),
.Y(n_10644)
);

OAI33xp33_ASAP7_75t_L g10645 ( 
.A1(n_9808),
.A2(n_9060),
.A3(n_9054),
.B1(n_9063),
.B2(n_9062),
.B3(n_9055),
.Y(n_10645)
);

CKINVDCx8_ASAP7_75t_R g10646 ( 
.A(n_9846),
.Y(n_10646)
);

INVxp67_ASAP7_75t_SL g10647 ( 
.A(n_9922),
.Y(n_10647)
);

AND2x2_ASAP7_75t_L g10648 ( 
.A(n_9988),
.B(n_8173),
.Y(n_10648)
);

AND2x2_ASAP7_75t_L g10649 ( 
.A(n_9923),
.B(n_6927),
.Y(n_10649)
);

AND2x2_ASAP7_75t_L g10650 ( 
.A(n_9930),
.B(n_6927),
.Y(n_10650)
);

NAND2xp5_ASAP7_75t_L g10651 ( 
.A(n_9781),
.B(n_9055),
.Y(n_10651)
);

AND2x2_ASAP7_75t_L g10652 ( 
.A(n_9935),
.B(n_6927),
.Y(n_10652)
);

INVx1_ASAP7_75t_L g10653 ( 
.A(n_10038),
.Y(n_10653)
);

OAI21xp5_ASAP7_75t_L g10654 ( 
.A1(n_9712),
.A2(n_9502),
.B(n_9624),
.Y(n_10654)
);

AND2x2_ASAP7_75t_L g10655 ( 
.A(n_9905),
.B(n_6935),
.Y(n_10655)
);

HB1xp67_ASAP7_75t_L g10656 ( 
.A(n_9728),
.Y(n_10656)
);

INVx2_ASAP7_75t_SL g10657 ( 
.A(n_10116),
.Y(n_10657)
);

INVx2_ASAP7_75t_L g10658 ( 
.A(n_10326),
.Y(n_10658)
);

INVx1_ASAP7_75t_L g10659 ( 
.A(n_10038),
.Y(n_10659)
);

AND2x4_ASAP7_75t_L g10660 ( 
.A(n_9869),
.B(n_9768),
.Y(n_10660)
);

BUFx3_ASAP7_75t_L g10661 ( 
.A(n_10017),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_10059),
.Y(n_10662)
);

INVx1_ASAP7_75t_L g10663 ( 
.A(n_10059),
.Y(n_10663)
);

BUFx2_ASAP7_75t_L g10664 ( 
.A(n_9843),
.Y(n_10664)
);

AND2x2_ASAP7_75t_L g10665 ( 
.A(n_9977),
.B(n_6935),
.Y(n_10665)
);

OR2x2_ASAP7_75t_L g10666 ( 
.A(n_10422),
.B(n_9301),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_10067),
.Y(n_10667)
);

HB1xp67_ASAP7_75t_L g10668 ( 
.A(n_10011),
.Y(n_10668)
);

AND2x4_ASAP7_75t_L g10669 ( 
.A(n_9869),
.B(n_9183),
.Y(n_10669)
);

INVx1_ASAP7_75t_L g10670 ( 
.A(n_10067),
.Y(n_10670)
);

AOI22xp5_ASAP7_75t_SL g10671 ( 
.A1(n_9708),
.A2(n_6806),
.B1(n_6804),
.B2(n_6842),
.Y(n_10671)
);

INVx5_ASAP7_75t_L g10672 ( 
.A(n_9737),
.Y(n_10672)
);

BUFx3_ASAP7_75t_L g10673 ( 
.A(n_9737),
.Y(n_10673)
);

INVx2_ASAP7_75t_L g10674 ( 
.A(n_10326),
.Y(n_10674)
);

HB1xp67_ASAP7_75t_L g10675 ( 
.A(n_10366),
.Y(n_10675)
);

INVx1_ASAP7_75t_L g10676 ( 
.A(n_10068),
.Y(n_10676)
);

INVx1_ASAP7_75t_L g10677 ( 
.A(n_10068),
.Y(n_10677)
);

INVx2_ASAP7_75t_L g10678 ( 
.A(n_10117),
.Y(n_10678)
);

INVx2_ASAP7_75t_L g10679 ( 
.A(n_9962),
.Y(n_10679)
);

INVx2_ASAP7_75t_L g10680 ( 
.A(n_9962),
.Y(n_10680)
);

INVx1_ASAP7_75t_L g10681 ( 
.A(n_10087),
.Y(n_10681)
);

INVx1_ASAP7_75t_L g10682 ( 
.A(n_10087),
.Y(n_10682)
);

AND2x2_ASAP7_75t_L g10683 ( 
.A(n_9715),
.B(n_6935),
.Y(n_10683)
);

BUFx2_ASAP7_75t_L g10684 ( 
.A(n_10244),
.Y(n_10684)
);

AND2x2_ASAP7_75t_L g10685 ( 
.A(n_9920),
.B(n_8324),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_10088),
.Y(n_10686)
);

AO31x2_ASAP7_75t_L g10687 ( 
.A1(n_10106),
.A2(n_9062),
.A3(n_9063),
.B(n_9060),
.Y(n_10687)
);

AND2x4_ASAP7_75t_L g10688 ( 
.A(n_9907),
.B(n_9186),
.Y(n_10688)
);

INVx2_ASAP7_75t_SL g10689 ( 
.A(n_10116),
.Y(n_10689)
);

AND2x2_ASAP7_75t_L g10690 ( 
.A(n_9759),
.B(n_9767),
.Y(n_10690)
);

AND2x2_ASAP7_75t_L g10691 ( 
.A(n_9775),
.B(n_8324),
.Y(n_10691)
);

INVx1_ASAP7_75t_L g10692 ( 
.A(n_10088),
.Y(n_10692)
);

INVx1_ASAP7_75t_L g10693 ( 
.A(n_10112),
.Y(n_10693)
);

BUFx6f_ASAP7_75t_L g10694 ( 
.A(n_9798),
.Y(n_10694)
);

AND2x2_ASAP7_75t_L g10695 ( 
.A(n_10009),
.B(n_8324),
.Y(n_10695)
);

INVx1_ASAP7_75t_L g10696 ( 
.A(n_10112),
.Y(n_10696)
);

AND2x2_ASAP7_75t_L g10697 ( 
.A(n_10026),
.B(n_8421),
.Y(n_10697)
);

AND2x2_ASAP7_75t_L g10698 ( 
.A(n_10033),
.B(n_8421),
.Y(n_10698)
);

INVx2_ASAP7_75t_SL g10699 ( 
.A(n_9822),
.Y(n_10699)
);

NAND2xp5_ASAP7_75t_L g10700 ( 
.A(n_9837),
.B(n_9064),
.Y(n_10700)
);

INVx1_ASAP7_75t_L g10701 ( 
.A(n_10131),
.Y(n_10701)
);

INVx1_ASAP7_75t_L g10702 ( 
.A(n_10131),
.Y(n_10702)
);

AND2x2_ASAP7_75t_L g10703 ( 
.A(n_10035),
.B(n_8421),
.Y(n_10703)
);

NAND2xp5_ASAP7_75t_SL g10704 ( 
.A(n_10204),
.B(n_7826),
.Y(n_10704)
);

INVx2_ASAP7_75t_L g10705 ( 
.A(n_10368),
.Y(n_10705)
);

AO31x2_ASAP7_75t_L g10706 ( 
.A1(n_10106),
.A2(n_9922),
.A3(n_9913),
.B(n_10398),
.Y(n_10706)
);

INVx2_ASAP7_75t_L g10707 ( 
.A(n_10368),
.Y(n_10707)
);

AND2x4_ASAP7_75t_L g10708 ( 
.A(n_9907),
.B(n_9186),
.Y(n_10708)
);

AND2x2_ASAP7_75t_L g10709 ( 
.A(n_10040),
.B(n_8421),
.Y(n_10709)
);

INVx2_ASAP7_75t_L g10710 ( 
.A(n_10371),
.Y(n_10710)
);

INVx1_ASAP7_75t_L g10711 ( 
.A(n_10161),
.Y(n_10711)
);

INVx4_ASAP7_75t_L g10712 ( 
.A(n_9822),
.Y(n_10712)
);

INVx1_ASAP7_75t_L g10713 ( 
.A(n_10161),
.Y(n_10713)
);

AOI31xp33_ASAP7_75t_L g10714 ( 
.A1(n_10060),
.A2(n_6997),
.A3(n_6844),
.B(n_6889),
.Y(n_10714)
);

INVx2_ASAP7_75t_L g10715 ( 
.A(n_10371),
.Y(n_10715)
);

INVx2_ASAP7_75t_L g10716 ( 
.A(n_9883),
.Y(n_10716)
);

INVx1_ASAP7_75t_L g10717 ( 
.A(n_10181),
.Y(n_10717)
);

INVx2_ASAP7_75t_L g10718 ( 
.A(n_9883),
.Y(n_10718)
);

BUFx2_ASAP7_75t_L g10719 ( 
.A(n_10244),
.Y(n_10719)
);

AOI22xp33_ASAP7_75t_L g10720 ( 
.A1(n_9802),
.A2(n_8103),
.B1(n_9673),
.B2(n_9650),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_9985),
.B(n_8421),
.Y(n_10721)
);

AND2x2_ASAP7_75t_L g10722 ( 
.A(n_9985),
.B(n_8731),
.Y(n_10722)
);

INVx1_ASAP7_75t_L g10723 ( 
.A(n_10181),
.Y(n_10723)
);

AND2x2_ASAP7_75t_L g10724 ( 
.A(n_9997),
.B(n_8731),
.Y(n_10724)
);

INVxp67_ASAP7_75t_L g10725 ( 
.A(n_10210),
.Y(n_10725)
);

NAND2xp5_ASAP7_75t_L g10726 ( 
.A(n_9842),
.B(n_9064),
.Y(n_10726)
);

NAND2xp5_ASAP7_75t_L g10727 ( 
.A(n_9899),
.B(n_9072),
.Y(n_10727)
);

INVx1_ASAP7_75t_L g10728 ( 
.A(n_10190),
.Y(n_10728)
);

OR2x2_ASAP7_75t_L g10729 ( 
.A(n_9719),
.B(n_9312),
.Y(n_10729)
);

INVx2_ASAP7_75t_L g10730 ( 
.A(n_10352),
.Y(n_10730)
);

OR2x2_ASAP7_75t_L g10731 ( 
.A(n_9748),
.B(n_9312),
.Y(n_10731)
);

OR2x2_ASAP7_75t_L g10732 ( 
.A(n_9823),
.B(n_9164),
.Y(n_10732)
);

AO31x2_ASAP7_75t_L g10733 ( 
.A1(n_9913),
.A2(n_9076),
.A3(n_9077),
.B(n_9072),
.Y(n_10733)
);

INVxp67_ASAP7_75t_L g10734 ( 
.A(n_9701),
.Y(n_10734)
);

AND2x4_ASAP7_75t_L g10735 ( 
.A(n_9710),
.B(n_9186),
.Y(n_10735)
);

BUFx3_ASAP7_75t_L g10736 ( 
.A(n_10049),
.Y(n_10736)
);

INVx2_ASAP7_75t_L g10737 ( 
.A(n_10352),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_10190),
.Y(n_10738)
);

INVx2_ASAP7_75t_L g10739 ( 
.A(n_10185),
.Y(n_10739)
);

OR2x2_ASAP7_75t_L g10740 ( 
.A(n_9749),
.B(n_9164),
.Y(n_10740)
);

INVx1_ASAP7_75t_L g10741 ( 
.A(n_10247),
.Y(n_10741)
);

OR2x2_ASAP7_75t_L g10742 ( 
.A(n_9839),
.B(n_9622),
.Y(n_10742)
);

AND2x4_ASAP7_75t_L g10743 ( 
.A(n_9710),
.B(n_9219),
.Y(n_10743)
);

INVx2_ASAP7_75t_L g10744 ( 
.A(n_10185),
.Y(n_10744)
);

OAI21xp5_ASAP7_75t_L g10745 ( 
.A1(n_9845),
.A2(n_9833),
.B(n_9716),
.Y(n_10745)
);

INVx2_ASAP7_75t_L g10746 ( 
.A(n_10209),
.Y(n_10746)
);

CKINVDCx16_ASAP7_75t_R g10747 ( 
.A(n_9919),
.Y(n_10747)
);

INVx2_ASAP7_75t_L g10748 ( 
.A(n_10209),
.Y(n_10748)
);

AND2x4_ASAP7_75t_SL g10749 ( 
.A(n_9997),
.B(n_10072),
.Y(n_10749)
);

AND2x2_ASAP7_75t_L g10750 ( 
.A(n_10072),
.B(n_8731),
.Y(n_10750)
);

AO21x2_ASAP7_75t_L g10751 ( 
.A1(n_9814),
.A2(n_9077),
.B(n_9076),
.Y(n_10751)
);

BUFx2_ASAP7_75t_L g10752 ( 
.A(n_10244),
.Y(n_10752)
);

INVx2_ASAP7_75t_L g10753 ( 
.A(n_10302),
.Y(n_10753)
);

AOI22xp33_ASAP7_75t_L g10754 ( 
.A1(n_9795),
.A2(n_8103),
.B1(n_9673),
.B2(n_9650),
.Y(n_10754)
);

INVx1_ASAP7_75t_L g10755 ( 
.A(n_10247),
.Y(n_10755)
);

HB1xp67_ASAP7_75t_L g10756 ( 
.A(n_9926),
.Y(n_10756)
);

INVx2_ASAP7_75t_L g10757 ( 
.A(n_10302),
.Y(n_10757)
);

INVx1_ASAP7_75t_L g10758 ( 
.A(n_10278),
.Y(n_10758)
);

NAND2x1_ASAP7_75t_L g10759 ( 
.A(n_9697),
.B(n_10328),
.Y(n_10759)
);

AND2x2_ASAP7_75t_L g10760 ( 
.A(n_10101),
.B(n_10166),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_10168),
.Y(n_10761)
);

HB1xp67_ASAP7_75t_L g10762 ( 
.A(n_9936),
.Y(n_10762)
);

NAND2xp5_ASAP7_75t_L g10763 ( 
.A(n_9992),
.B(n_9082),
.Y(n_10763)
);

AND2x2_ASAP7_75t_L g10764 ( 
.A(n_10101),
.B(n_8731),
.Y(n_10764)
);

OAI22xp5_ASAP7_75t_L g10765 ( 
.A1(n_9713),
.A2(n_7796),
.B1(n_6745),
.B2(n_6747),
.Y(n_10765)
);

AND2x2_ASAP7_75t_L g10766 ( 
.A(n_10166),
.B(n_8731),
.Y(n_10766)
);

INVx2_ASAP7_75t_L g10767 ( 
.A(n_10168),
.Y(n_10767)
);

NOR2x1_ASAP7_75t_SL g10768 ( 
.A(n_10279),
.B(n_7406),
.Y(n_10768)
);

INVx1_ASAP7_75t_L g10769 ( 
.A(n_10278),
.Y(n_10769)
);

INVx3_ASAP7_75t_L g10770 ( 
.A(n_10061),
.Y(n_10770)
);

INVx2_ASAP7_75t_L g10771 ( 
.A(n_10184),
.Y(n_10771)
);

INVx2_ASAP7_75t_L g10772 ( 
.A(n_9765),
.Y(n_10772)
);

AND2x2_ASAP7_75t_L g10773 ( 
.A(n_9979),
.B(n_8806),
.Y(n_10773)
);

INVx1_ASAP7_75t_L g10774 ( 
.A(n_10341),
.Y(n_10774)
);

AND2x2_ASAP7_75t_L g10775 ( 
.A(n_10214),
.B(n_8806),
.Y(n_10775)
);

INVx2_ASAP7_75t_L g10776 ( 
.A(n_10184),
.Y(n_10776)
);

INVx2_ASAP7_75t_L g10777 ( 
.A(n_10199),
.Y(n_10777)
);

INVx1_ASAP7_75t_L g10778 ( 
.A(n_10341),
.Y(n_10778)
);

INVx1_ASAP7_75t_L g10779 ( 
.A(n_10363),
.Y(n_10779)
);

AND2x2_ASAP7_75t_L g10780 ( 
.A(n_10321),
.B(n_8806),
.Y(n_10780)
);

INVx2_ASAP7_75t_L g10781 ( 
.A(n_10199),
.Y(n_10781)
);

INVx2_ASAP7_75t_L g10782 ( 
.A(n_10224),
.Y(n_10782)
);

INVx2_ASAP7_75t_L g10783 ( 
.A(n_10224),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_L g10784 ( 
.A(n_10036),
.B(n_9082),
.Y(n_10784)
);

OR2x2_ASAP7_75t_L g10785 ( 
.A(n_9984),
.B(n_9622),
.Y(n_10785)
);

INVx5_ASAP7_75t_L g10786 ( 
.A(n_9798),
.Y(n_10786)
);

BUFx2_ASAP7_75t_L g10787 ( 
.A(n_10244),
.Y(n_10787)
);

INVx2_ASAP7_75t_L g10788 ( 
.A(n_10232),
.Y(n_10788)
);

AOI22xp33_ASAP7_75t_L g10789 ( 
.A1(n_9840),
.A2(n_8103),
.B1(n_9673),
.B2(n_9650),
.Y(n_10789)
);

INVx2_ASAP7_75t_L g10790 ( 
.A(n_10232),
.Y(n_10790)
);

AOI21xp5_ASAP7_75t_L g10791 ( 
.A1(n_9705),
.A2(n_9206),
.B(n_9502),
.Y(n_10791)
);

OR2x2_ASAP7_75t_L g10792 ( 
.A(n_9971),
.B(n_9692),
.Y(n_10792)
);

NOR2xp33_ASAP7_75t_L g10793 ( 
.A(n_10051),
.B(n_6986),
.Y(n_10793)
);

AND2x2_ASAP7_75t_L g10794 ( 
.A(n_10354),
.B(n_8806),
.Y(n_10794)
);

INVx1_ASAP7_75t_L g10795 ( 
.A(n_10363),
.Y(n_10795)
);

INVx2_ASAP7_75t_L g10796 ( 
.A(n_10249),
.Y(n_10796)
);

INVx4_ASAP7_75t_L g10797 ( 
.A(n_9924),
.Y(n_10797)
);

AOI22xp33_ASAP7_75t_SL g10798 ( 
.A1(n_9743),
.A2(n_9206),
.B1(n_7899),
.B2(n_8368),
.Y(n_10798)
);

AND2x2_ASAP7_75t_L g10799 ( 
.A(n_9735),
.B(n_8660),
.Y(n_10799)
);

BUFx3_ASAP7_75t_L g10800 ( 
.A(n_10049),
.Y(n_10800)
);

INVx2_ASAP7_75t_L g10801 ( 
.A(n_10249),
.Y(n_10801)
);

INVx2_ASAP7_75t_L g10802 ( 
.A(n_10255),
.Y(n_10802)
);

AND2x2_ASAP7_75t_L g10803 ( 
.A(n_9938),
.B(n_8678),
.Y(n_10803)
);

INVx1_ASAP7_75t_L g10804 ( 
.A(n_10412),
.Y(n_10804)
);

INVx5_ASAP7_75t_L g10805 ( 
.A(n_9924),
.Y(n_10805)
);

AND2x2_ASAP7_75t_L g10806 ( 
.A(n_9945),
.B(n_8678),
.Y(n_10806)
);

INVx4_ASAP7_75t_R g10807 ( 
.A(n_9750),
.Y(n_10807)
);

BUFx2_ASAP7_75t_SL g10808 ( 
.A(n_9889),
.Y(n_10808)
);

INVx2_ASAP7_75t_L g10809 ( 
.A(n_10255),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_10412),
.Y(n_10810)
);

INVx2_ASAP7_75t_L g10811 ( 
.A(n_10025),
.Y(n_10811)
);

INVx2_ASAP7_75t_L g10812 ( 
.A(n_10025),
.Y(n_10812)
);

INVxp67_ASAP7_75t_SL g10813 ( 
.A(n_10398),
.Y(n_10813)
);

INVx1_ASAP7_75t_SL g10814 ( 
.A(n_9717),
.Y(n_10814)
);

NAND2xp5_ASAP7_75t_L g10815 ( 
.A(n_10043),
.B(n_9093),
.Y(n_10815)
);

AND2x2_ASAP7_75t_L g10816 ( 
.A(n_10139),
.B(n_10140),
.Y(n_10816)
);

INVx1_ASAP7_75t_L g10817 ( 
.A(n_10437),
.Y(n_10817)
);

AND2x2_ASAP7_75t_L g10818 ( 
.A(n_10141),
.B(n_8678),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_10437),
.Y(n_10819)
);

HB1xp67_ASAP7_75t_L g10820 ( 
.A(n_10048),
.Y(n_10820)
);

INVx2_ASAP7_75t_L g10821 ( 
.A(n_10025),
.Y(n_10821)
);

INVx1_ASAP7_75t_L g10822 ( 
.A(n_10441),
.Y(n_10822)
);

BUFx3_ASAP7_75t_L g10823 ( 
.A(n_10049),
.Y(n_10823)
);

INVx1_ASAP7_75t_L g10824 ( 
.A(n_10441),
.Y(n_10824)
);

AO21x2_ASAP7_75t_L g10825 ( 
.A1(n_10357),
.A2(n_9094),
.B(n_9093),
.Y(n_10825)
);

INVx1_ASAP7_75t_L g10826 ( 
.A(n_10306),
.Y(n_10826)
);

AND2x2_ASAP7_75t_L g10827 ( 
.A(n_10154),
.B(n_8678),
.Y(n_10827)
);

CKINVDCx12_ASAP7_75t_R g10828 ( 
.A(n_10085),
.Y(n_10828)
);

INVx2_ASAP7_75t_L g10829 ( 
.A(n_10358),
.Y(n_10829)
);

NAND2xp5_ASAP7_75t_L g10830 ( 
.A(n_10079),
.B(n_9094),
.Y(n_10830)
);

AND2x2_ASAP7_75t_L g10831 ( 
.A(n_10156),
.B(n_8678),
.Y(n_10831)
);

INVx1_ASAP7_75t_L g10832 ( 
.A(n_10313),
.Y(n_10832)
);

INVx1_ASAP7_75t_L g10833 ( 
.A(n_10338),
.Y(n_10833)
);

BUFx3_ASAP7_75t_L g10834 ( 
.A(n_10049),
.Y(n_10834)
);

INVx4_ASAP7_75t_L g10835 ( 
.A(n_9924),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_10395),
.Y(n_10836)
);

INVx2_ASAP7_75t_L g10837 ( 
.A(n_9717),
.Y(n_10837)
);

INVx1_ASAP7_75t_L g10838 ( 
.A(n_10407),
.Y(n_10838)
);

INVx2_ASAP7_75t_L g10839 ( 
.A(n_10337),
.Y(n_10839)
);

AND2x2_ASAP7_75t_L g10840 ( 
.A(n_10158),
.B(n_10164),
.Y(n_10840)
);

INVx1_ASAP7_75t_L g10841 ( 
.A(n_10104),
.Y(n_10841)
);

AND2x4_ASAP7_75t_L g10842 ( 
.A(n_9736),
.B(n_9219),
.Y(n_10842)
);

INVx2_ASAP7_75t_L g10843 ( 
.A(n_10337),
.Y(n_10843)
);

INVx2_ASAP7_75t_SL g10844 ( 
.A(n_10086),
.Y(n_10844)
);

HB1xp67_ASAP7_75t_L g10845 ( 
.A(n_10157),
.Y(n_10845)
);

INVx2_ASAP7_75t_L g10846 ( 
.A(n_10122),
.Y(n_10846)
);

NAND2xp5_ASAP7_75t_L g10847 ( 
.A(n_10348),
.B(n_9096),
.Y(n_10847)
);

INVx1_ASAP7_75t_L g10848 ( 
.A(n_9848),
.Y(n_10848)
);

BUFx2_ASAP7_75t_L g10849 ( 
.A(n_9697),
.Y(n_10849)
);

INVx1_ASAP7_75t_L g10850 ( 
.A(n_9872),
.Y(n_10850)
);

NAND2xp5_ASAP7_75t_L g10851 ( 
.A(n_9730),
.B(n_9096),
.Y(n_10851)
);

AND2x2_ASAP7_75t_L g10852 ( 
.A(n_10170),
.B(n_8754),
.Y(n_10852)
);

BUFx2_ASAP7_75t_L g10853 ( 
.A(n_10149),
.Y(n_10853)
);

AND2x2_ASAP7_75t_L g10854 ( 
.A(n_9747),
.B(n_8754),
.Y(n_10854)
);

NAND2xp5_ASAP7_75t_L g10855 ( 
.A(n_9917),
.B(n_9098),
.Y(n_10855)
);

INVx1_ASAP7_75t_L g10856 ( 
.A(n_9895),
.Y(n_10856)
);

INVx1_ASAP7_75t_SL g10857 ( 
.A(n_10109),
.Y(n_10857)
);

BUFx2_ASAP7_75t_L g10858 ( 
.A(n_10240),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_9696),
.Y(n_10859)
);

INVx1_ASAP7_75t_L g10860 ( 
.A(n_9706),
.Y(n_10860)
);

INVx2_ASAP7_75t_L g10861 ( 
.A(n_10122),
.Y(n_10861)
);

AND2x4_ASAP7_75t_SL g10862 ( 
.A(n_9727),
.B(n_6677),
.Y(n_10862)
);

INVx2_ASAP7_75t_L g10863 ( 
.A(n_10125),
.Y(n_10863)
);

INVx2_ASAP7_75t_L g10864 ( 
.A(n_10125),
.Y(n_10864)
);

AND2x4_ASAP7_75t_L g10865 ( 
.A(n_9736),
.B(n_9219),
.Y(n_10865)
);

AND2x2_ASAP7_75t_L g10866 ( 
.A(n_10042),
.B(n_8754),
.Y(n_10866)
);

INVx2_ASAP7_75t_L g10867 ( 
.A(n_10251),
.Y(n_10867)
);

INVx2_ASAP7_75t_L g10868 ( 
.A(n_10057),
.Y(n_10868)
);

NOR2xp33_ASAP7_75t_L g10869 ( 
.A(n_10051),
.B(n_6822),
.Y(n_10869)
);

NAND2xp5_ASAP7_75t_L g10870 ( 
.A(n_9954),
.B(n_9098),
.Y(n_10870)
);

AND2x2_ASAP7_75t_L g10871 ( 
.A(n_9779),
.B(n_8754),
.Y(n_10871)
);

BUFx6f_ASAP7_75t_L g10872 ( 
.A(n_9873),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_9772),
.Y(n_10873)
);

AND2x2_ASAP7_75t_L g10874 ( 
.A(n_10047),
.B(n_8754),
.Y(n_10874)
);

HB1xp67_ASAP7_75t_L g10875 ( 
.A(n_10282),
.Y(n_10875)
);

NAND2xp5_ASAP7_75t_L g10876 ( 
.A(n_10350),
.B(n_9948),
.Y(n_10876)
);

AND2x4_ASAP7_75t_L g10877 ( 
.A(n_9755),
.B(n_9290),
.Y(n_10877)
);

AND2x2_ASAP7_75t_L g10878 ( 
.A(n_10058),
.B(n_6677),
.Y(n_10878)
);

AND2x2_ASAP7_75t_L g10879 ( 
.A(n_9788),
.B(n_6736),
.Y(n_10879)
);

OAI22xp5_ASAP7_75t_L g10880 ( 
.A1(n_9793),
.A2(n_7796),
.B1(n_6928),
.B2(n_7623),
.Y(n_10880)
);

AND2x2_ASAP7_75t_L g10881 ( 
.A(n_9797),
.B(n_6736),
.Y(n_10881)
);

AND2x2_ASAP7_75t_L g10882 ( 
.A(n_10126),
.B(n_6736),
.Y(n_10882)
);

INVx2_ASAP7_75t_L g10883 ( 
.A(n_10057),
.Y(n_10883)
);

NOR2x1_ASAP7_75t_SL g10884 ( 
.A(n_10159),
.B(n_7406),
.Y(n_10884)
);

INVx2_ASAP7_75t_L g10885 ( 
.A(n_9953),
.Y(n_10885)
);

INVx1_ASAP7_75t_L g10886 ( 
.A(n_9799),
.Y(n_10886)
);

OAI22xp5_ASAP7_75t_L g10887 ( 
.A1(n_9762),
.A2(n_9850),
.B1(n_10350),
.B2(n_9902),
.Y(n_10887)
);

OR2x2_ASAP7_75t_L g10888 ( 
.A(n_9811),
.B(n_9692),
.Y(n_10888)
);

INVx1_ASAP7_75t_L g10889 ( 
.A(n_9807),
.Y(n_10889)
);

AND2x2_ASAP7_75t_L g10890 ( 
.A(n_10128),
.B(n_6736),
.Y(n_10890)
);

INVx1_ASAP7_75t_L g10891 ( 
.A(n_9834),
.Y(n_10891)
);

INVx1_ASAP7_75t_L g10892 ( 
.A(n_9885),
.Y(n_10892)
);

OR2x2_ASAP7_75t_L g10893 ( 
.A(n_9956),
.B(n_8823),
.Y(n_10893)
);

INVx1_ASAP7_75t_L g10894 ( 
.A(n_9893),
.Y(n_10894)
);

OR2x2_ASAP7_75t_L g10895 ( 
.A(n_9994),
.B(n_8823),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_10130),
.B(n_6969),
.Y(n_10896)
);

INVx1_ASAP7_75t_L g10897 ( 
.A(n_9906),
.Y(n_10897)
);

OR2x2_ASAP7_75t_L g10898 ( 
.A(n_10195),
.B(n_8826),
.Y(n_10898)
);

INVx1_ASAP7_75t_L g10899 ( 
.A(n_9921),
.Y(n_10899)
);

BUFx3_ASAP7_75t_L g10900 ( 
.A(n_9933),
.Y(n_10900)
);

INVx1_ASAP7_75t_L g10901 ( 
.A(n_9929),
.Y(n_10901)
);

BUFx3_ASAP7_75t_L g10902 ( 
.A(n_9937),
.Y(n_10902)
);

NAND4xp25_ASAP7_75t_L g10903 ( 
.A(n_9841),
.B(n_6689),
.C(n_7130),
.D(n_7051),
.Y(n_10903)
);

INVx1_ASAP7_75t_L g10904 ( 
.A(n_9947),
.Y(n_10904)
);

CKINVDCx5p33_ASAP7_75t_R g10905 ( 
.A(n_10186),
.Y(n_10905)
);

NAND2xp5_ASAP7_75t_L g10906 ( 
.A(n_10052),
.B(n_9100),
.Y(n_10906)
);

NAND2xp5_ASAP7_75t_L g10907 ( 
.A(n_10083),
.B(n_9100),
.Y(n_10907)
);

NOR2xp33_ASAP7_75t_L g10908 ( 
.A(n_9873),
.B(n_6822),
.Y(n_10908)
);

AOI22xp33_ASAP7_75t_SL g10909 ( 
.A1(n_9741),
.A2(n_7899),
.B1(n_8368),
.B2(n_9624),
.Y(n_10909)
);

INVx1_ASAP7_75t_L g10910 ( 
.A(n_9958),
.Y(n_10910)
);

AND2x2_ASAP7_75t_L g10911 ( 
.A(n_9745),
.B(n_10066),
.Y(n_10911)
);

AND2x4_ASAP7_75t_L g10912 ( 
.A(n_9755),
.B(n_9290),
.Y(n_10912)
);

AND2x2_ASAP7_75t_L g10913 ( 
.A(n_10069),
.B(n_6969),
.Y(n_10913)
);

NAND2xp5_ASAP7_75t_L g10914 ( 
.A(n_10173),
.B(n_9103),
.Y(n_10914)
);

HB1xp67_ASAP7_75t_L g10915 ( 
.A(n_10291),
.Y(n_10915)
);

INVx1_ASAP7_75t_L g10916 ( 
.A(n_9963),
.Y(n_10916)
);

INVx1_ASAP7_75t_L g10917 ( 
.A(n_9968),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_9998),
.Y(n_10918)
);

HB1xp67_ASAP7_75t_L g10919 ( 
.A(n_10292),
.Y(n_10919)
);

INVx1_ASAP7_75t_L g10920 ( 
.A(n_10001),
.Y(n_10920)
);

BUFx6f_ASAP7_75t_L g10921 ( 
.A(n_9816),
.Y(n_10921)
);

INVxp67_ASAP7_75t_SL g10922 ( 
.A(n_9944),
.Y(n_10922)
);

AND2x4_ASAP7_75t_SL g10923 ( 
.A(n_9727),
.B(n_6969),
.Y(n_10923)
);

INVxp67_ASAP7_75t_L g10924 ( 
.A(n_10024),
.Y(n_10924)
);

INVx2_ASAP7_75t_L g10925 ( 
.A(n_9953),
.Y(n_10925)
);

OAI222xp33_ASAP7_75t_L g10926 ( 
.A1(n_9875),
.A2(n_9646),
.B1(n_8819),
.B2(n_6928),
.C1(n_7629),
.C2(n_7680),
.Y(n_10926)
);

AOI22xp33_ASAP7_75t_L g10927 ( 
.A1(n_9800),
.A2(n_7814),
.B1(n_7838),
.B2(n_7899),
.Y(n_10927)
);

AND2x2_ASAP7_75t_L g10928 ( 
.A(n_10078),
.B(n_6969),
.Y(n_10928)
);

NAND2xp5_ASAP7_75t_L g10929 ( 
.A(n_10056),
.B(n_9103),
.Y(n_10929)
);

INVx1_ASAP7_75t_L g10930 ( 
.A(n_10094),
.Y(n_10930)
);

BUFx3_ASAP7_75t_L g10931 ( 
.A(n_9964),
.Y(n_10931)
);

INVx1_ASAP7_75t_L g10932 ( 
.A(n_10096),
.Y(n_10932)
);

BUFx3_ASAP7_75t_L g10933 ( 
.A(n_9783),
.Y(n_10933)
);

OR2x2_ASAP7_75t_L g10934 ( 
.A(n_9761),
.B(n_8826),
.Y(n_10934)
);

AND2x2_ASAP7_75t_L g10935 ( 
.A(n_10080),
.B(n_8828),
.Y(n_10935)
);

INVx1_ASAP7_75t_L g10936 ( 
.A(n_10107),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_10137),
.Y(n_10937)
);

INVx2_ASAP7_75t_SL g10938 ( 
.A(n_9757),
.Y(n_10938)
);

AND2x2_ASAP7_75t_L g10939 ( 
.A(n_10081),
.B(n_8828),
.Y(n_10939)
);

INVx1_ASAP7_75t_L g10940 ( 
.A(n_10138),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_10177),
.Y(n_10941)
);

AND2x2_ASAP7_75t_L g10942 ( 
.A(n_10084),
.B(n_10089),
.Y(n_10942)
);

OR2x2_ASAP7_75t_L g10943 ( 
.A(n_9782),
.B(n_8834),
.Y(n_10943)
);

AND2x2_ASAP7_75t_L g10944 ( 
.A(n_10110),
.B(n_8834),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_10201),
.Y(n_10945)
);

BUFx3_ASAP7_75t_L g10946 ( 
.A(n_9757),
.Y(n_10946)
);

INVx2_ASAP7_75t_L g10947 ( 
.A(n_9765),
.Y(n_10947)
);

INVx2_ASAP7_75t_L g10948 ( 
.A(n_9927),
.Y(n_10948)
);

AOI22xp33_ASAP7_75t_L g10949 ( 
.A1(n_9738),
.A2(n_7814),
.B1(n_7838),
.B2(n_7126),
.Y(n_10949)
);

AND2x2_ASAP7_75t_L g10950 ( 
.A(n_10120),
.B(n_8835),
.Y(n_10950)
);

AND2x2_ASAP7_75t_L g10951 ( 
.A(n_10111),
.B(n_8835),
.Y(n_10951)
);

NAND2xp5_ASAP7_75t_L g10952 ( 
.A(n_10211),
.B(n_9107),
.Y(n_10952)
);

INVx2_ASAP7_75t_L g10953 ( 
.A(n_9927),
.Y(n_10953)
);

AND2x2_ASAP7_75t_L g10954 ( 
.A(n_9951),
.B(n_8840),
.Y(n_10954)
);

INVx2_ASAP7_75t_L g10955 ( 
.A(n_9959),
.Y(n_10955)
);

INVx1_ASAP7_75t_L g10956 ( 
.A(n_10231),
.Y(n_10956)
);

INVx1_ASAP7_75t_L g10957 ( 
.A(n_10238),
.Y(n_10957)
);

INVx1_ASAP7_75t_L g10958 ( 
.A(n_10243),
.Y(n_10958)
);

INVx2_ASAP7_75t_L g10959 ( 
.A(n_9959),
.Y(n_10959)
);

INVx2_ASAP7_75t_L g10960 ( 
.A(n_10133),
.Y(n_10960)
);

AND2x2_ASAP7_75t_L g10961 ( 
.A(n_10276),
.B(n_8840),
.Y(n_10961)
);

AND2x2_ASAP7_75t_L g10962 ( 
.A(n_10276),
.B(n_8845),
.Y(n_10962)
);

AND2x4_ASAP7_75t_SL g10963 ( 
.A(n_10207),
.B(n_7032),
.Y(n_10963)
);

AND2x2_ASAP7_75t_L g10964 ( 
.A(n_10176),
.B(n_8845),
.Y(n_10964)
);

NAND2xp5_ASAP7_75t_L g10965 ( 
.A(n_10277),
.B(n_9107),
.Y(n_10965)
);

INVx2_ASAP7_75t_L g10966 ( 
.A(n_9953),
.Y(n_10966)
);

AND2x2_ASAP7_75t_L g10967 ( 
.A(n_10187),
.B(n_8848),
.Y(n_10967)
);

INVx2_ASAP7_75t_L g10968 ( 
.A(n_10005),
.Y(n_10968)
);

NAND3xp33_ASAP7_75t_L g10969 ( 
.A(n_10039),
.B(n_8312),
.C(n_9624),
.Y(n_10969)
);

INVx2_ASAP7_75t_L g10970 ( 
.A(n_10005),
.Y(n_10970)
);

AND2x2_ASAP7_75t_L g10971 ( 
.A(n_10188),
.B(n_8848),
.Y(n_10971)
);

AND2x2_ASAP7_75t_L g10972 ( 
.A(n_10219),
.B(n_8849),
.Y(n_10972)
);

INVx1_ASAP7_75t_L g10973 ( 
.A(n_10196),
.Y(n_10973)
);

INVxp67_ASAP7_75t_SL g10974 ( 
.A(n_10357),
.Y(n_10974)
);

AND2x2_ASAP7_75t_L g10975 ( 
.A(n_10222),
.B(n_8849),
.Y(n_10975)
);

OAI21xp33_ASAP7_75t_L g10976 ( 
.A1(n_9975),
.A2(n_9646),
.B(n_6686),
.Y(n_10976)
);

INVx2_ASAP7_75t_L g10977 ( 
.A(n_10005),
.Y(n_10977)
);

INVx1_ASAP7_75t_L g10978 ( 
.A(n_10202),
.Y(n_10978)
);

INVx1_ASAP7_75t_L g10979 ( 
.A(n_10206),
.Y(n_10979)
);

INVx1_ASAP7_75t_L g10980 ( 
.A(n_10233),
.Y(n_10980)
);

INVx2_ASAP7_75t_L g10981 ( 
.A(n_10369),
.Y(n_10981)
);

INVx1_ASAP7_75t_L g10982 ( 
.A(n_10248),
.Y(n_10982)
);

AND2x2_ASAP7_75t_L g10983 ( 
.A(n_10225),
.B(n_8868),
.Y(n_10983)
);

NAND2xp5_ASAP7_75t_L g10984 ( 
.A(n_10182),
.B(n_9108),
.Y(n_10984)
);

INVx1_ASAP7_75t_SL g10985 ( 
.A(n_9763),
.Y(n_10985)
);

AND2x2_ASAP7_75t_L g10986 ( 
.A(n_10227),
.B(n_8868),
.Y(n_10986)
);

HB1xp67_ASAP7_75t_L g10987 ( 
.A(n_10312),
.Y(n_10987)
);

AND2x2_ASAP7_75t_L g10988 ( 
.A(n_10229),
.B(n_8869),
.Y(n_10988)
);

AND2x2_ASAP7_75t_L g10989 ( 
.A(n_10241),
.B(n_8869),
.Y(n_10989)
);

INVx2_ASAP7_75t_L g10990 ( 
.A(n_10298),
.Y(n_10990)
);

BUFx6f_ASAP7_75t_L g10991 ( 
.A(n_9821),
.Y(n_10991)
);

BUFx6f_ASAP7_75t_L g10992 ( 
.A(n_9832),
.Y(n_10992)
);

AND2x2_ASAP7_75t_L g10993 ( 
.A(n_10246),
.B(n_10268),
.Y(n_10993)
);

INVx2_ASAP7_75t_L g10994 ( 
.A(n_10360),
.Y(n_10994)
);

INVx2_ASAP7_75t_L g10995 ( 
.A(n_10361),
.Y(n_10995)
);

AND2x2_ASAP7_75t_L g10996 ( 
.A(n_10272),
.B(n_8870),
.Y(n_10996)
);

INVx2_ASAP7_75t_L g10997 ( 
.A(n_10365),
.Y(n_10997)
);

OAI221xp5_ASAP7_75t_L g10998 ( 
.A1(n_10108),
.A2(n_7130),
.B1(n_7143),
.B2(n_7051),
.C(n_7155),
.Y(n_10998)
);

INVx1_ASAP7_75t_L g10999 ( 
.A(n_10253),
.Y(n_10999)
);

INVx2_ASAP7_75t_L g11000 ( 
.A(n_10384),
.Y(n_11000)
);

INVx2_ASAP7_75t_L g11001 ( 
.A(n_10386),
.Y(n_11001)
);

INVx2_ASAP7_75t_L g11002 ( 
.A(n_10392),
.Y(n_11002)
);

INVx2_ASAP7_75t_L g11003 ( 
.A(n_10399),
.Y(n_11003)
);

AND2x2_ASAP7_75t_L g11004 ( 
.A(n_10281),
.B(n_8870),
.Y(n_11004)
);

INVx1_ASAP7_75t_L g11005 ( 
.A(n_9763),
.Y(n_11005)
);

AND2x2_ASAP7_75t_L g11006 ( 
.A(n_10290),
.B(n_8871),
.Y(n_11006)
);

NAND2xp5_ASAP7_75t_L g11007 ( 
.A(n_10031),
.B(n_9108),
.Y(n_11007)
);

INVx1_ASAP7_75t_L g11008 ( 
.A(n_9778),
.Y(n_11008)
);

BUFx2_ASAP7_75t_L g11009 ( 
.A(n_9778),
.Y(n_11009)
);

INVx1_ASAP7_75t_L g11010 ( 
.A(n_9787),
.Y(n_11010)
);

INVx1_ASAP7_75t_L g11011 ( 
.A(n_9787),
.Y(n_11011)
);

HB1xp67_ASAP7_75t_L g11012 ( 
.A(n_9849),
.Y(n_11012)
);

INVx1_ASAP7_75t_L g11013 ( 
.A(n_9844),
.Y(n_11013)
);

INVx1_ASAP7_75t_L g11014 ( 
.A(n_9844),
.Y(n_11014)
);

AND2x2_ASAP7_75t_L g11015 ( 
.A(n_10295),
.B(n_8871),
.Y(n_11015)
);

AND2x2_ASAP7_75t_L g11016 ( 
.A(n_10301),
.B(n_8872),
.Y(n_11016)
);

NOR2xp67_ASAP7_75t_L g11017 ( 
.A(n_9742),
.B(n_9290),
.Y(n_11017)
);

INVx2_ASAP7_75t_SL g11018 ( 
.A(n_9854),
.Y(n_11018)
);

INVx2_ASAP7_75t_L g11019 ( 
.A(n_10405),
.Y(n_11019)
);

AND2x2_ASAP7_75t_L g11020 ( 
.A(n_10308),
.B(n_8872),
.Y(n_11020)
);

BUFx2_ASAP7_75t_L g11021 ( 
.A(n_9854),
.Y(n_11021)
);

OR2x2_ASAP7_75t_L g11022 ( 
.A(n_9794),
.B(n_8874),
.Y(n_11022)
);

BUFx6f_ASAP7_75t_L g11023 ( 
.A(n_9901),
.Y(n_11023)
);

AND2x2_ASAP7_75t_L g11024 ( 
.A(n_10310),
.B(n_8874),
.Y(n_11024)
);

NOR2x1_ASAP7_75t_SL g11025 ( 
.A(n_9756),
.B(n_9914),
.Y(n_11025)
);

AND2x2_ASAP7_75t_L g11026 ( 
.A(n_10311),
.B(n_7051),
.Y(n_11026)
);

INVx2_ASAP7_75t_SL g11027 ( 
.A(n_9879),
.Y(n_11027)
);

BUFx3_ASAP7_75t_L g11028 ( 
.A(n_9879),
.Y(n_11028)
);

AO21x2_ASAP7_75t_L g11029 ( 
.A1(n_10250),
.A2(n_9113),
.B(n_9109),
.Y(n_11029)
);

HB1xp67_ASAP7_75t_L g11030 ( 
.A(n_10335),
.Y(n_11030)
);

AND2x2_ASAP7_75t_L g11031 ( 
.A(n_10314),
.B(n_7051),
.Y(n_11031)
);

HB1xp67_ASAP7_75t_L g11032 ( 
.A(n_10344),
.Y(n_11032)
);

INVx1_ASAP7_75t_L g11033 ( 
.A(n_10376),
.Y(n_11033)
);

AO31x2_ASAP7_75t_L g11034 ( 
.A1(n_10250),
.A2(n_9113),
.A3(n_9114),
.B(n_9109),
.Y(n_11034)
);

AND2x2_ASAP7_75t_L g11035 ( 
.A(n_10316),
.B(n_7130),
.Y(n_11035)
);

AND2x2_ASAP7_75t_L g11036 ( 
.A(n_10334),
.B(n_7130),
.Y(n_11036)
);

NAND2xp5_ASAP7_75t_L g11037 ( 
.A(n_10213),
.B(n_9114),
.Y(n_11037)
);

NAND2xp5_ASAP7_75t_L g11038 ( 
.A(n_10006),
.B(n_9118),
.Y(n_11038)
);

INVxp67_ASAP7_75t_SL g11039 ( 
.A(n_10351),
.Y(n_11039)
);

HB1xp67_ASAP7_75t_L g11040 ( 
.A(n_10377),
.Y(n_11040)
);

INVxp67_ASAP7_75t_L g11041 ( 
.A(n_10150),
.Y(n_11041)
);

HB1xp67_ASAP7_75t_L g11042 ( 
.A(n_10381),
.Y(n_11042)
);

OR2x2_ASAP7_75t_L g11043 ( 
.A(n_10178),
.B(n_9021),
.Y(n_11043)
);

INVx1_ASAP7_75t_L g11044 ( 
.A(n_10383),
.Y(n_11044)
);

OR2x2_ASAP7_75t_L g11045 ( 
.A(n_10374),
.B(n_9021),
.Y(n_11045)
);

INVx1_ASAP7_75t_L g11046 ( 
.A(n_10396),
.Y(n_11046)
);

OR2x2_ASAP7_75t_L g11047 ( 
.A(n_10375),
.B(n_8875),
.Y(n_11047)
);

OR2x2_ASAP7_75t_L g11048 ( 
.A(n_10385),
.B(n_8875),
.Y(n_11048)
);

NAND2xp5_ASAP7_75t_L g11049 ( 
.A(n_10427),
.B(n_9118),
.Y(n_11049)
);

BUFx2_ASAP7_75t_L g11050 ( 
.A(n_9909),
.Y(n_11050)
);

INVx1_ASAP7_75t_L g11051 ( 
.A(n_10343),
.Y(n_11051)
);

INVx1_ASAP7_75t_L g11052 ( 
.A(n_10364),
.Y(n_11052)
);

INVx2_ASAP7_75t_L g11053 ( 
.A(n_10409),
.Y(n_11053)
);

INVx1_ASAP7_75t_L g11054 ( 
.A(n_10014),
.Y(n_11054)
);

AND2x2_ASAP7_75t_L g11055 ( 
.A(n_10339),
.B(n_7143),
.Y(n_11055)
);

NOR2x1_ASAP7_75t_SL g11056 ( 
.A(n_10064),
.B(n_6989),
.Y(n_11056)
);

INVx2_ASAP7_75t_L g11057 ( 
.A(n_10411),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10014),
.Y(n_11058)
);

NOR4xp25_ASAP7_75t_SL g11059 ( 
.A(n_10329),
.B(n_6864),
.C(n_7129),
.D(n_8627),
.Y(n_11059)
);

AND2x2_ASAP7_75t_L g11060 ( 
.A(n_10346),
.B(n_7143),
.Y(n_11060)
);

OR2x2_ASAP7_75t_L g11061 ( 
.A(n_10075),
.B(n_8876),
.Y(n_11061)
);

AND2x2_ASAP7_75t_L g11062 ( 
.A(n_10355),
.B(n_7143),
.Y(n_11062)
);

INVx1_ASAP7_75t_L g11063 ( 
.A(n_10014),
.Y(n_11063)
);

AND2x2_ASAP7_75t_L g11064 ( 
.A(n_10356),
.B(n_10134),
.Y(n_11064)
);

INVx1_ASAP7_75t_L g11065 ( 
.A(n_10074),
.Y(n_11065)
);

INVx2_ASAP7_75t_SL g11066 ( 
.A(n_9909),
.Y(n_11066)
);

NAND2xp5_ASAP7_75t_SL g11067 ( 
.A(n_9916),
.B(n_7826),
.Y(n_11067)
);

AOI22xp33_ASAP7_75t_L g11068 ( 
.A1(n_9876),
.A2(n_7814),
.B1(n_7838),
.B2(n_7126),
.Y(n_11068)
);

INVx1_ASAP7_75t_L g11069 ( 
.A(n_10284),
.Y(n_11069)
);

AND2x2_ASAP7_75t_L g11070 ( 
.A(n_10194),
.B(n_8876),
.Y(n_11070)
);

INVx1_ASAP7_75t_L g11071 ( 
.A(n_10285),
.Y(n_11071)
);

AND2x2_ASAP7_75t_L g11072 ( 
.A(n_10102),
.B(n_8877),
.Y(n_11072)
);

AND2x2_ASAP7_75t_L g11073 ( 
.A(n_10309),
.B(n_8877),
.Y(n_11073)
);

OR2x2_ASAP7_75t_L g11074 ( 
.A(n_10082),
.B(n_8887),
.Y(n_11074)
);

INVx1_ASAP7_75t_L g11075 ( 
.A(n_10397),
.Y(n_11075)
);

INVx2_ASAP7_75t_L g11076 ( 
.A(n_10413),
.Y(n_11076)
);

AND2x2_ASAP7_75t_L g11077 ( 
.A(n_9818),
.B(n_8887),
.Y(n_11077)
);

INVx2_ASAP7_75t_L g11078 ( 
.A(n_10414),
.Y(n_11078)
);

AND2x4_ASAP7_75t_L g11079 ( 
.A(n_9903),
.B(n_8433),
.Y(n_11079)
);

AND2x2_ASAP7_75t_L g11080 ( 
.A(n_9853),
.B(n_8889),
.Y(n_11080)
);

AND2x2_ASAP7_75t_L g11081 ( 
.A(n_10286),
.B(n_10256),
.Y(n_11081)
);

NAND2xp5_ASAP7_75t_L g11082 ( 
.A(n_10442),
.B(n_9121),
.Y(n_11082)
);

AOI22xp33_ASAP7_75t_L g11083 ( 
.A1(n_10260),
.A2(n_7838),
.B1(n_7814),
.B2(n_9652),
.Y(n_11083)
);

INVx2_ASAP7_75t_SL g11084 ( 
.A(n_10015),
.Y(n_11084)
);

INVx1_ASAP7_75t_L g11085 ( 
.A(n_10404),
.Y(n_11085)
);

AND2x2_ASAP7_75t_L g11086 ( 
.A(n_10258),
.B(n_8889),
.Y(n_11086)
);

AND2x4_ASAP7_75t_L g11087 ( 
.A(n_9966),
.B(n_8450),
.Y(n_11087)
);

INVxp67_ASAP7_75t_L g11088 ( 
.A(n_10163),
.Y(n_11088)
);

INVx1_ASAP7_75t_L g11089 ( 
.A(n_10347),
.Y(n_11089)
);

BUFx2_ASAP7_75t_L g11090 ( 
.A(n_10015),
.Y(n_11090)
);

NOR2x1_ASAP7_75t_SL g11091 ( 
.A(n_9820),
.B(n_9949),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10347),
.Y(n_11092)
);

HB1xp67_ASAP7_75t_L g11093 ( 
.A(n_10237),
.Y(n_11093)
);

AND2x2_ASAP7_75t_L g11094 ( 
.A(n_9969),
.B(n_8896),
.Y(n_11094)
);

INVx2_ASAP7_75t_L g11095 ( 
.A(n_10418),
.Y(n_11095)
);

INVx2_ASAP7_75t_L g11096 ( 
.A(n_10431),
.Y(n_11096)
);

INVx1_ASAP7_75t_L g11097 ( 
.A(n_10347),
.Y(n_11097)
);

INVx1_ASAP7_75t_L g11098 ( 
.A(n_10193),
.Y(n_11098)
);

OR2x2_ASAP7_75t_L g11099 ( 
.A(n_10444),
.B(n_10197),
.Y(n_11099)
);

AND2x2_ASAP7_75t_L g11100 ( 
.A(n_9973),
.B(n_8896),
.Y(n_11100)
);

INVx1_ASAP7_75t_L g11101 ( 
.A(n_10421),
.Y(n_11101)
);

INVx1_ASAP7_75t_L g11102 ( 
.A(n_10421),
.Y(n_11102)
);

BUFx3_ASAP7_75t_L g11103 ( 
.A(n_10076),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_10421),
.Y(n_11104)
);

INVx2_ASAP7_75t_L g11105 ( 
.A(n_10434),
.Y(n_11105)
);

AND2x2_ASAP7_75t_L g11106 ( 
.A(n_10002),
.B(n_8904),
.Y(n_11106)
);

HB1xp67_ASAP7_75t_L g11107 ( 
.A(n_10378),
.Y(n_11107)
);

NOR2xp33_ASAP7_75t_L g11108 ( 
.A(n_10217),
.B(n_6890),
.Y(n_11108)
);

INVx1_ASAP7_75t_L g11109 ( 
.A(n_10054),
.Y(n_11109)
);

BUFx2_ASAP7_75t_L g11110 ( 
.A(n_10034),
.Y(n_11110)
);

BUFx2_ASAP7_75t_L g11111 ( 
.A(n_10034),
.Y(n_11111)
);

INVx1_ASAP7_75t_L g11112 ( 
.A(n_10054),
.Y(n_11112)
);

AND2x4_ASAP7_75t_L g11113 ( 
.A(n_10003),
.B(n_8450),
.Y(n_11113)
);

NAND2xp5_ASAP7_75t_L g11114 ( 
.A(n_10423),
.B(n_9121),
.Y(n_11114)
);

AND2x2_ASAP7_75t_L g11115 ( 
.A(n_10324),
.B(n_8904),
.Y(n_11115)
);

INVx1_ASAP7_75t_L g11116 ( 
.A(n_10054),
.Y(n_11116)
);

INVx2_ASAP7_75t_L g11117 ( 
.A(n_9721),
.Y(n_11117)
);

NAND2xp5_ASAP7_75t_L g11118 ( 
.A(n_10010),
.B(n_9124),
.Y(n_11118)
);

INVx1_ASAP7_75t_L g11119 ( 
.A(n_10212),
.Y(n_11119)
);

INVx2_ASAP7_75t_L g11120 ( 
.A(n_9721),
.Y(n_11120)
);

NAND2xp5_ASAP7_75t_L g11121 ( 
.A(n_10297),
.B(n_9124),
.Y(n_11121)
);

INVx2_ASAP7_75t_L g11122 ( 
.A(n_9829),
.Y(n_11122)
);

AND2x2_ASAP7_75t_L g11123 ( 
.A(n_10283),
.B(n_8906),
.Y(n_11123)
);

INVx2_ASAP7_75t_L g11124 ( 
.A(n_9829),
.Y(n_11124)
);

OR2x2_ASAP7_75t_L g11125 ( 
.A(n_10223),
.B(n_8906),
.Y(n_11125)
);

INVxp67_ASAP7_75t_L g11126 ( 
.A(n_10077),
.Y(n_11126)
);

OA21x2_ASAP7_75t_L g11127 ( 
.A1(n_10340),
.A2(n_9209),
.B(n_9144),
.Y(n_11127)
);

AND2x2_ASAP7_75t_L g11128 ( 
.A(n_10236),
.B(n_8908),
.Y(n_11128)
);

AND2x2_ASAP7_75t_L g11129 ( 
.A(n_10296),
.B(n_8908),
.Y(n_11129)
);

AND2x2_ASAP7_75t_L g11130 ( 
.A(n_10439),
.B(n_8914),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_L g11131 ( 
.A(n_10391),
.B(n_9126),
.Y(n_11131)
);

INVx1_ASAP7_75t_L g11132 ( 
.A(n_10257),
.Y(n_11132)
);

AND2x2_ASAP7_75t_L g11133 ( 
.A(n_10529),
.B(n_10151),
.Y(n_11133)
);

AND2x2_ASAP7_75t_L g11134 ( 
.A(n_10593),
.B(n_9809),
.Y(n_11134)
);

NAND2xp5_ASAP7_75t_L g11135 ( 
.A(n_10585),
.B(n_10315),
.Y(n_11135)
);

AND2x2_ASAP7_75t_L g11136 ( 
.A(n_10573),
.B(n_10200),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_L g11137 ( 
.A(n_10585),
.B(n_10606),
.Y(n_11137)
);

NOR2xp33_ASAP7_75t_L g11138 ( 
.A(n_10536),
.B(n_9766),
.Y(n_11138)
);

OAI22xp5_ASAP7_75t_L g11139 ( 
.A1(n_10515),
.A2(n_9851),
.B1(n_9803),
.B2(n_10175),
.Y(n_11139)
);

OAI221xp5_ASAP7_75t_SL g11140 ( 
.A1(n_10515),
.A2(n_10440),
.B1(n_10266),
.B2(n_10153),
.C(n_9897),
.Y(n_11140)
);

AND2x2_ASAP7_75t_L g11141 ( 
.A(n_10573),
.B(n_10165),
.Y(n_11141)
);

NAND3xp33_ASAP7_75t_L g11142 ( 
.A(n_10603),
.B(n_10146),
.C(n_9911),
.Y(n_11142)
);

OAI21xp5_ASAP7_75t_SL g11143 ( 
.A1(n_10745),
.A2(n_9817),
.B(n_9858),
.Y(n_11143)
);

NAND2xp5_ASAP7_75t_L g11144 ( 
.A(n_10606),
.B(n_10267),
.Y(n_11144)
);

NAND2xp5_ASAP7_75t_L g11145 ( 
.A(n_10668),
.B(n_10029),
.Y(n_11145)
);

AOI22xp33_ASAP7_75t_SL g11146 ( 
.A1(n_10887),
.A2(n_10162),
.B1(n_10121),
.B2(n_10362),
.Y(n_11146)
);

NOR2xp67_ASAP7_75t_L g11147 ( 
.A(n_10463),
.B(n_9835),
.Y(n_11147)
);

NAND4xp25_ASAP7_75t_L g11148 ( 
.A(n_10745),
.B(n_10021),
.C(n_10288),
.D(n_9867),
.Y(n_11148)
);

NAND2xp5_ASAP7_75t_L g11149 ( 
.A(n_10668),
.B(n_10095),
.Y(n_11149)
);

AND2x2_ASAP7_75t_L g11150 ( 
.A(n_10661),
.B(n_10191),
.Y(n_11150)
);

AOI21xp5_ASAP7_75t_L g11151 ( 
.A1(n_10599),
.A2(n_9890),
.B(n_10030),
.Y(n_11151)
);

NAND3xp33_ASAP7_75t_L g11152 ( 
.A(n_10603),
.B(n_10216),
.C(n_10379),
.Y(n_11152)
);

AND2x2_ASAP7_75t_L g11153 ( 
.A(n_10661),
.B(n_10092),
.Y(n_11153)
);

AND2x2_ASAP7_75t_L g11154 ( 
.A(n_10524),
.B(n_10132),
.Y(n_11154)
);

NAND2xp5_ASAP7_75t_L g11155 ( 
.A(n_10448),
.B(n_9884),
.Y(n_11155)
);

NAND3xp33_ASAP7_75t_L g11156 ( 
.A(n_10656),
.B(n_10198),
.C(n_10123),
.Y(n_11156)
);

AND2x2_ASAP7_75t_SL g11157 ( 
.A(n_10551),
.B(n_10660),
.Y(n_11157)
);

AND2x2_ASAP7_75t_L g11158 ( 
.A(n_10857),
.B(n_9943),
.Y(n_11158)
);

NAND3xp33_ASAP7_75t_L g11159 ( 
.A(n_10656),
.B(n_9978),
.C(n_9864),
.Y(n_11159)
);

NAND2xp5_ASAP7_75t_L g11160 ( 
.A(n_10454),
.B(n_10380),
.Y(n_11160)
);

NAND2xp5_ASAP7_75t_L g11161 ( 
.A(n_10462),
.B(n_9855),
.Y(n_11161)
);

NOR3xp33_ASAP7_75t_L g11162 ( 
.A(n_10887),
.B(n_10294),
.C(n_9934),
.Y(n_11162)
);

AND2x2_ASAP7_75t_L g11163 ( 
.A(n_10857),
.B(n_9886),
.Y(n_11163)
);

NAND2xp5_ASAP7_75t_L g11164 ( 
.A(n_10473),
.B(n_9928),
.Y(n_11164)
);

AND2x2_ASAP7_75t_L g11165 ( 
.A(n_10625),
.B(n_9776),
.Y(n_11165)
);

NAND2xp5_ASAP7_75t_L g11166 ( 
.A(n_10734),
.B(n_8819),
.Y(n_11166)
);

AOI22xp33_ASAP7_75t_SL g11167 ( 
.A1(n_11025),
.A2(n_10599),
.B1(n_11091),
.B2(n_10765),
.Y(n_11167)
);

AOI22xp33_ASAP7_75t_L g11168 ( 
.A1(n_10765),
.A2(n_9931),
.B1(n_10016),
.B2(n_9925),
.Y(n_11168)
);

AND2x2_ASAP7_75t_SL g11169 ( 
.A(n_10551),
.B(n_10023),
.Y(n_11169)
);

NAND2xp5_ASAP7_75t_SL g11170 ( 
.A(n_10467),
.B(n_10234),
.Y(n_11170)
);

NAND3xp33_ASAP7_75t_L g11171 ( 
.A(n_10467),
.B(n_9896),
.C(n_9877),
.Y(n_11171)
);

OAI221xp5_ASAP7_75t_SL g11172 ( 
.A1(n_10520),
.A2(n_10228),
.B1(n_10416),
.B2(n_9862),
.C(n_10046),
.Y(n_11172)
);

NAND2xp5_ASAP7_75t_L g11173 ( 
.A(n_10734),
.B(n_8819),
.Y(n_11173)
);

NAND2xp5_ASAP7_75t_L g11174 ( 
.A(n_10814),
.B(n_8819),
.Y(n_11174)
);

NAND2xp5_ASAP7_75t_L g11175 ( 
.A(n_10814),
.B(n_10564),
.Y(n_11175)
);

NAND2xp5_ASAP7_75t_L g11176 ( 
.A(n_10564),
.B(n_8819),
.Y(n_11176)
);

OAI221xp5_ASAP7_75t_L g11177 ( 
.A1(n_10571),
.A2(n_9868),
.B1(n_10044),
.B2(n_10037),
.C(n_10091),
.Y(n_11177)
);

AOI22xp5_ASAP7_75t_L g11178 ( 
.A1(n_10571),
.A2(n_9932),
.B1(n_9996),
.B2(n_10018),
.Y(n_11178)
);

AND2x2_ASAP7_75t_L g11179 ( 
.A(n_10536),
.B(n_9776),
.Y(n_11179)
);

NAND2xp5_ASAP7_75t_L g11180 ( 
.A(n_10583),
.B(n_10443),
.Y(n_11180)
);

OAI221xp5_ASAP7_75t_SL g11181 ( 
.A1(n_10520),
.A2(n_9967),
.B1(n_10400),
.B2(n_10433),
.C(n_10073),
.Y(n_11181)
);

AOI22xp33_ASAP7_75t_SL g11182 ( 
.A1(n_10671),
.A2(n_10121),
.B1(n_10162),
.B2(n_10362),
.Y(n_11182)
);

AOI22xp33_ASAP7_75t_L g11183 ( 
.A1(n_10880),
.A2(n_10008),
.B1(n_10167),
.B2(n_10147),
.Y(n_11183)
);

NAND3xp33_ASAP7_75t_L g11184 ( 
.A(n_10720),
.B(n_9993),
.C(n_10370),
.Y(n_11184)
);

NAND2xp5_ASAP7_75t_L g11185 ( 
.A(n_10583),
.B(n_10013),
.Y(n_11185)
);

AOI22xp5_ASAP7_75t_L g11186 ( 
.A1(n_10880),
.A2(n_9991),
.B1(n_9960),
.B2(n_10245),
.Y(n_11186)
);

OA21x2_ASAP7_75t_L g11187 ( 
.A1(n_10791),
.A2(n_10432),
.B(n_10353),
.Y(n_11187)
);

OAI22xp5_ASAP7_75t_L g11188 ( 
.A1(n_10720),
.A2(n_10789),
.B1(n_10754),
.B2(n_10476),
.Y(n_11188)
);

NAND2xp5_ASAP7_75t_L g11189 ( 
.A(n_10447),
.B(n_10408),
.Y(n_11189)
);

NAND3xp33_ASAP7_75t_L g11190 ( 
.A(n_10789),
.B(n_10235),
.C(n_10280),
.Y(n_11190)
);

OA21x2_ASAP7_75t_L g11191 ( 
.A1(n_10791),
.A2(n_10429),
.B(n_9847),
.Y(n_11191)
);

NAND2xp5_ASAP7_75t_L g11192 ( 
.A(n_10447),
.B(n_10382),
.Y(n_11192)
);

NAND2xp5_ASAP7_75t_SL g11193 ( 
.A(n_10536),
.B(n_10262),
.Y(n_11193)
);

NAND2xp5_ASAP7_75t_L g11194 ( 
.A(n_10452),
.B(n_10388),
.Y(n_11194)
);

NAND2xp5_ASAP7_75t_L g11195 ( 
.A(n_10452),
.B(n_10545),
.Y(n_11195)
);

NAND2xp5_ASAP7_75t_L g11196 ( 
.A(n_10545),
.B(n_10390),
.Y(n_11196)
);

NAND4xp25_ASAP7_75t_L g11197 ( 
.A(n_10851),
.B(n_10359),
.C(n_10041),
.D(n_10269),
.Y(n_11197)
);

NAND2xp5_ASAP7_75t_L g11198 ( 
.A(n_10558),
.B(n_10858),
.Y(n_11198)
);

AND2x2_ASAP7_75t_L g11199 ( 
.A(n_10642),
.B(n_9776),
.Y(n_11199)
);

AND2x2_ASAP7_75t_L g11200 ( 
.A(n_10660),
.B(n_9805),
.Y(n_11200)
);

NAND2xp5_ASAP7_75t_SL g11201 ( 
.A(n_10798),
.B(n_9957),
.Y(n_11201)
);

OAI221xp5_ASAP7_75t_L g11202 ( 
.A1(n_10903),
.A2(n_10203),
.B1(n_10022),
.B2(n_10007),
.C(n_10055),
.Y(n_11202)
);

NOR2xp33_ASAP7_75t_R g11203 ( 
.A(n_10580),
.B(n_6989),
.Y(n_11203)
);

NOR2xp33_ASAP7_75t_L g11204 ( 
.A(n_10457),
.B(n_6890),
.Y(n_11204)
);

INVx2_ASAP7_75t_L g11205 ( 
.A(n_10451),
.Y(n_11205)
);

AOI22xp33_ASAP7_75t_SL g11206 ( 
.A1(n_10671),
.A2(n_9805),
.B1(n_10119),
.B2(n_10372),
.Y(n_11206)
);

AND2x2_ASAP7_75t_L g11207 ( 
.A(n_10579),
.B(n_9805),
.Y(n_11207)
);

NAND2xp5_ASAP7_75t_L g11208 ( 
.A(n_10558),
.B(n_10402),
.Y(n_11208)
);

NAND2xp5_ASAP7_75t_L g11209 ( 
.A(n_10479),
.B(n_10417),
.Y(n_11209)
);

INVx1_ASAP7_75t_L g11210 ( 
.A(n_10587),
.Y(n_11210)
);

NAND3xp33_ASAP7_75t_L g11211 ( 
.A(n_10922),
.B(n_10430),
.C(n_9982),
.Y(n_11211)
);

INVx1_ASAP7_75t_L g11212 ( 
.A(n_10587),
.Y(n_11212)
);

AOI22xp33_ASAP7_75t_SL g11213 ( 
.A1(n_10751),
.A2(n_10144),
.B1(n_10172),
.B2(n_10424),
.Y(n_11213)
);

NAND2xp5_ASAP7_75t_L g11214 ( 
.A(n_10482),
.B(n_10287),
.Y(n_11214)
);

NOR3xp33_ASAP7_75t_L g11215 ( 
.A(n_10747),
.B(n_10259),
.C(n_10438),
.Y(n_11215)
);

AOI22xp33_ASAP7_75t_SL g11216 ( 
.A1(n_10751),
.A2(n_10420),
.B1(n_10299),
.B2(n_10171),
.Y(n_11216)
);

NAND3xp33_ASAP7_75t_L g11217 ( 
.A(n_10922),
.B(n_11012),
.C(n_10458),
.Y(n_11217)
);

NAND3xp33_ASAP7_75t_L g11218 ( 
.A(n_11012),
.B(n_10304),
.C(n_10275),
.Y(n_11218)
);

OAI22xp5_ASAP7_75t_L g11219 ( 
.A1(n_10754),
.A2(n_7623),
.B1(n_7629),
.B2(n_7597),
.Y(n_11219)
);

AND2x2_ASAP7_75t_L g11220 ( 
.A(n_10808),
.B(n_9835),
.Y(n_11220)
);

NAND2xp5_ASAP7_75t_L g11221 ( 
.A(n_10484),
.B(n_10328),
.Y(n_11221)
);

OAI221xp5_ASAP7_75t_L g11222 ( 
.A1(n_10903),
.A2(n_10263),
.B1(n_10090),
.B2(n_10065),
.C(n_10105),
.Y(n_11222)
);

NAND3xp33_ASAP7_75t_L g11223 ( 
.A(n_10458),
.B(n_10271),
.C(n_10336),
.Y(n_11223)
);

NAND2xp5_ASAP7_75t_L g11224 ( 
.A(n_10487),
.B(n_10328),
.Y(n_11224)
);

NAND4xp25_ASAP7_75t_L g11225 ( 
.A(n_10851),
.B(n_10428),
.C(n_10289),
.D(n_10100),
.Y(n_11225)
);

NAND2xp5_ASAP7_75t_L g11226 ( 
.A(n_10494),
.B(n_10500),
.Y(n_11226)
);

NAND3xp33_ASAP7_75t_L g11227 ( 
.A(n_10847),
.B(n_10476),
.C(n_10566),
.Y(n_11227)
);

AND2x2_ASAP7_75t_L g11228 ( 
.A(n_10690),
.B(n_7032),
.Y(n_11228)
);

NAND2xp5_ASAP7_75t_L g11229 ( 
.A(n_10489),
.B(n_10328),
.Y(n_11229)
);

AND2x2_ASAP7_75t_L g11230 ( 
.A(n_10595),
.B(n_10816),
.Y(n_11230)
);

NAND3xp33_ASAP7_75t_L g11231 ( 
.A(n_10798),
.B(n_10342),
.C(n_10221),
.Y(n_11231)
);

NAND2xp5_ASAP7_75t_L g11232 ( 
.A(n_10489),
.B(n_10032),
.Y(n_11232)
);

OAI22xp5_ASAP7_75t_L g11233 ( 
.A1(n_10568),
.A2(n_7697),
.B1(n_7721),
.B2(n_7680),
.Y(n_11233)
);

NAND2xp5_ASAP7_75t_L g11234 ( 
.A(n_10506),
.B(n_10160),
.Y(n_11234)
);

AOI221xp5_ASAP7_75t_L g11235 ( 
.A1(n_10645),
.A2(n_10566),
.B1(n_10926),
.B2(n_10468),
.C(n_10654),
.Y(n_11235)
);

OAI221xp5_ASAP7_75t_SL g11236 ( 
.A1(n_11068),
.A2(n_10332),
.B1(n_10230),
.B2(n_10393),
.C(n_10387),
.Y(n_11236)
);

AND2x2_ASAP7_75t_L g11237 ( 
.A(n_10840),
.B(n_10525),
.Y(n_11237)
);

NAND2xp5_ASAP7_75t_L g11238 ( 
.A(n_10506),
.B(n_10406),
.Y(n_11238)
);

NOR2xp33_ASAP7_75t_L g11239 ( 
.A(n_10457),
.B(n_10580),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_10522),
.B(n_10318),
.Y(n_11240)
);

NAND2xp5_ASAP7_75t_L g11241 ( 
.A(n_10522),
.B(n_10327),
.Y(n_11241)
);

OA211x2_ASAP7_75t_L g11242 ( 
.A1(n_10759),
.A2(n_11108),
.B(n_10976),
.C(n_10704),
.Y(n_11242)
);

AND2x2_ASAP7_75t_L g11243 ( 
.A(n_10853),
.B(n_7032),
.Y(n_11243)
);

OAI21xp5_ASAP7_75t_SL g11244 ( 
.A1(n_10714),
.A2(n_10415),
.B(n_6841),
.Y(n_11244)
);

OAI21xp5_ASAP7_75t_SL g11245 ( 
.A1(n_10714),
.A2(n_6841),
.B(n_10205),
.Y(n_11245)
);

NOR2xp33_ASAP7_75t_L g11246 ( 
.A(n_10457),
.B(n_6890),
.Y(n_11246)
);

AND2x2_ASAP7_75t_L g11247 ( 
.A(n_10466),
.B(n_11064),
.Y(n_11247)
);

NAND2xp5_ASAP7_75t_L g11248 ( 
.A(n_10530),
.B(n_9037),
.Y(n_11248)
);

NAND3xp33_ASAP7_75t_L g11249 ( 
.A(n_10568),
.B(n_10654),
.C(n_10909),
.Y(n_11249)
);

AND2x2_ASAP7_75t_L g11250 ( 
.A(n_10449),
.B(n_7032),
.Y(n_11250)
);

INVx1_ASAP7_75t_L g11251 ( 
.A(n_10530),
.Y(n_11251)
);

INVx2_ASAP7_75t_L g11252 ( 
.A(n_10451),
.Y(n_11252)
);

AND2x2_ASAP7_75t_L g11253 ( 
.A(n_10508),
.B(n_9037),
.Y(n_11253)
);

OAI221xp5_ASAP7_75t_SL g11254 ( 
.A1(n_11068),
.A2(n_10394),
.B1(n_10426),
.B2(n_10425),
.C(n_10401),
.Y(n_11254)
);

AND2x2_ASAP7_75t_L g11255 ( 
.A(n_10509),
.B(n_9041),
.Y(n_11255)
);

OAI221xp5_ASAP7_75t_SL g11256 ( 
.A1(n_10949),
.A2(n_10436),
.B1(n_6729),
.B2(n_7161),
.C(n_6782),
.Y(n_11256)
);

NAND2xp5_ASAP7_75t_L g11257 ( 
.A(n_10477),
.B(n_9041),
.Y(n_11257)
);

OAI21xp5_ASAP7_75t_SL g11258 ( 
.A1(n_10926),
.A2(n_10215),
.B(n_10208),
.Y(n_11258)
);

INVx1_ASAP7_75t_L g11259 ( 
.A(n_10756),
.Y(n_11259)
);

NAND2xp5_ASAP7_75t_L g11260 ( 
.A(n_10478),
.B(n_9044),
.Y(n_11260)
);

NAND2xp5_ASAP7_75t_L g11261 ( 
.A(n_10985),
.B(n_9044),
.Y(n_11261)
);

NAND2xp5_ASAP7_75t_L g11262 ( 
.A(n_10985),
.B(n_9049),
.Y(n_11262)
);

NAND2xp5_ASAP7_75t_L g11263 ( 
.A(n_10675),
.B(n_10455),
.Y(n_11263)
);

AND2x2_ASAP7_75t_L g11264 ( 
.A(n_10517),
.B(n_9049),
.Y(n_11264)
);

NAND3xp33_ASAP7_75t_L g11265 ( 
.A(n_10909),
.B(n_10317),
.C(n_10305),
.Y(n_11265)
);

OAI21xp5_ASAP7_75t_L g11266 ( 
.A1(n_10976),
.A2(n_9796),
.B(n_10226),
.Y(n_11266)
);

NAND3xp33_ASAP7_75t_L g11267 ( 
.A(n_10468),
.B(n_10345),
.C(n_9674),
.Y(n_11267)
);

NAND2xp5_ASAP7_75t_SL g11268 ( 
.A(n_10556),
.B(n_10463),
.Y(n_11268)
);

NAND2xp5_ASAP7_75t_L g11269 ( 
.A(n_10675),
.B(n_9058),
.Y(n_11269)
);

NAND2xp5_ASAP7_75t_L g11270 ( 
.A(n_10456),
.B(n_9058),
.Y(n_11270)
);

AND2x2_ASAP7_75t_L g11271 ( 
.A(n_10481),
.B(n_9073),
.Y(n_11271)
);

NAND2xp5_ASAP7_75t_SL g11272 ( 
.A(n_10463),
.B(n_10115),
.Y(n_11272)
);

AND2x2_ASAP7_75t_L g11273 ( 
.A(n_10488),
.B(n_10749),
.Y(n_11273)
);

NAND2xp5_ASAP7_75t_L g11274 ( 
.A(n_10459),
.B(n_9073),
.Y(n_11274)
);

AND2x2_ASAP7_75t_L g11275 ( 
.A(n_10749),
.B(n_8914),
.Y(n_11275)
);

AND2x2_ASAP7_75t_L g11276 ( 
.A(n_10854),
.B(n_8927),
.Y(n_11276)
);

NAND2xp5_ASAP7_75t_L g11277 ( 
.A(n_10464),
.B(n_10367),
.Y(n_11277)
);

AND2x2_ASAP7_75t_L g11278 ( 
.A(n_10446),
.B(n_8927),
.Y(n_11278)
);

AND2x2_ASAP7_75t_L g11279 ( 
.A(n_10445),
.B(n_8935),
.Y(n_11279)
);

OAI21xp5_ASAP7_75t_SL g11280 ( 
.A1(n_11108),
.A2(n_7118),
.B(n_7520),
.Y(n_11280)
);

NAND2xp5_ASAP7_75t_L g11281 ( 
.A(n_10739),
.B(n_10331),
.Y(n_11281)
);

AND2x2_ASAP7_75t_L g11282 ( 
.A(n_10483),
.B(n_8935),
.Y(n_11282)
);

NAND2xp5_ASAP7_75t_L g11283 ( 
.A(n_10744),
.B(n_10678),
.Y(n_11283)
);

NOR3xp33_ASAP7_75t_L g11284 ( 
.A(n_10505),
.B(n_9338),
.C(n_9324),
.Y(n_11284)
);

NAND2xp5_ASAP7_75t_L g11285 ( 
.A(n_11039),
.B(n_8938),
.Y(n_11285)
);

NAND2xp5_ASAP7_75t_L g11286 ( 
.A(n_11039),
.B(n_8938),
.Y(n_11286)
);

AND2x2_ASAP7_75t_L g11287 ( 
.A(n_10485),
.B(n_8942),
.Y(n_11287)
);

AND2x2_ASAP7_75t_L g11288 ( 
.A(n_10760),
.B(n_8942),
.Y(n_11288)
);

OAI22xp5_ASAP7_75t_L g11289 ( 
.A1(n_11059),
.A2(n_7721),
.B1(n_7738),
.B2(n_7697),
.Y(n_11289)
);

OAI221xp5_ASAP7_75t_SL g11290 ( 
.A1(n_10949),
.A2(n_6796),
.B1(n_6685),
.B2(n_7162),
.C(n_7756),
.Y(n_11290)
);

AND2x2_ASAP7_75t_L g11291 ( 
.A(n_10844),
.B(n_8950),
.Y(n_11291)
);

OAI22xp5_ASAP7_75t_L g11292 ( 
.A1(n_11059),
.A2(n_7764),
.B1(n_7778),
.B2(n_7738),
.Y(n_11292)
);

NAND3xp33_ASAP7_75t_L g11293 ( 
.A(n_10453),
.B(n_9674),
.C(n_9652),
.Y(n_11293)
);

OAI22xp5_ASAP7_75t_L g11294 ( 
.A1(n_10974),
.A2(n_7778),
.B1(n_7786),
.B2(n_7764),
.Y(n_11294)
);

NAND2xp5_ASAP7_75t_SL g11295 ( 
.A(n_10463),
.B(n_10183),
.Y(n_11295)
);

NAND2xp5_ASAP7_75t_L g11296 ( 
.A(n_11126),
.B(n_8950),
.Y(n_11296)
);

OAI22xp5_ASAP7_75t_L g11297 ( 
.A1(n_10974),
.A2(n_7786),
.B1(n_7594),
.B2(n_7624),
.Y(n_11297)
);

NAND2xp5_ASAP7_75t_SL g11298 ( 
.A(n_10615),
.B(n_7109),
.Y(n_11298)
);

AND2x2_ASAP7_75t_L g11299 ( 
.A(n_11103),
.B(n_8951),
.Y(n_11299)
);

NAND4xp25_ASAP7_75t_L g11300 ( 
.A(n_10453),
.B(n_10330),
.C(n_7546),
.D(n_7551),
.Y(n_11300)
);

NAND3xp33_ASAP7_75t_L g11301 ( 
.A(n_10927),
.B(n_9674),
.C(n_9652),
.Y(n_11301)
);

AND2x2_ASAP7_75t_L g11302 ( 
.A(n_11103),
.B(n_8951),
.Y(n_11302)
);

NAND2xp5_ASAP7_75t_L g11303 ( 
.A(n_11126),
.B(n_8958),
.Y(n_11303)
);

AND2x2_ASAP7_75t_L g11304 ( 
.A(n_10523),
.B(n_8958),
.Y(n_11304)
);

INVx2_ASAP7_75t_L g11305 ( 
.A(n_10604),
.Y(n_11305)
);

NAND2xp5_ASAP7_75t_L g11306 ( 
.A(n_10849),
.B(n_8960),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_10879),
.B(n_8960),
.Y(n_11307)
);

NOR2xp33_ASAP7_75t_R g11308 ( 
.A(n_10646),
.B(n_7040),
.Y(n_11308)
);

NAND2xp5_ASAP7_75t_L g11309 ( 
.A(n_10491),
.B(n_8961),
.Y(n_11309)
);

NAND2xp5_ASAP7_75t_L g11310 ( 
.A(n_10491),
.B(n_8961),
.Y(n_11310)
);

NAND3xp33_ASAP7_75t_L g11311 ( 
.A(n_10927),
.B(n_9680),
.C(n_9674),
.Y(n_11311)
);

NAND2xp5_ASAP7_75t_L g11312 ( 
.A(n_11009),
.B(n_8963),
.Y(n_11312)
);

OAI21xp5_ASAP7_75t_SL g11313 ( 
.A1(n_10497),
.A2(n_7282),
.B(n_7153),
.Y(n_11313)
);

NAND2x1p5_ASAP7_75t_L g11314 ( 
.A(n_10615),
.B(n_7083),
.Y(n_11314)
);

OAI221xp5_ASAP7_75t_SL g11315 ( 
.A1(n_10984),
.A2(n_9477),
.B1(n_9507),
.B2(n_9492),
.C(n_9446),
.Y(n_11315)
);

NAND2xp5_ASAP7_75t_L g11316 ( 
.A(n_11021),
.B(n_8963),
.Y(n_11316)
);

OAI21xp5_ASAP7_75t_L g11317 ( 
.A1(n_10969),
.A2(n_10179),
.B(n_8537),
.Y(n_11317)
);

NAND2xp5_ASAP7_75t_L g11318 ( 
.A(n_10867),
.B(n_8969),
.Y(n_11318)
);

AND2x2_ASAP7_75t_L g11319 ( 
.A(n_10881),
.B(n_8969),
.Y(n_11319)
);

OAI21xp5_ASAP7_75t_SL g11320 ( 
.A1(n_10497),
.A2(n_7138),
.B(n_7306),
.Y(n_11320)
);

NAND2xp5_ASAP7_75t_L g11321 ( 
.A(n_10924),
.B(n_8985),
.Y(n_11321)
);

AOI22xp33_ASAP7_75t_L g11322 ( 
.A1(n_10645),
.A2(n_7838),
.B1(n_7814),
.B2(n_7951),
.Y(n_11322)
);

AND2x2_ASAP7_75t_L g11323 ( 
.A(n_10803),
.B(n_8985),
.Y(n_11323)
);

OAI21xp33_ASAP7_75t_L g11324 ( 
.A1(n_10537),
.A2(n_10145),
.B(n_10124),
.Y(n_11324)
);

NAND2xp5_ASAP7_75t_L g11325 ( 
.A(n_10924),
.B(n_8986),
.Y(n_11325)
);

INVx1_ASAP7_75t_L g11326 ( 
.A(n_10756),
.Y(n_11326)
);

AND2x2_ASAP7_75t_L g11327 ( 
.A(n_10806),
.B(n_8986),
.Y(n_11327)
);

AOI221xp5_ASAP7_75t_L g11328 ( 
.A1(n_10847),
.A2(n_9131),
.B1(n_9135),
.B2(n_9130),
.C(n_9126),
.Y(n_11328)
);

AND2x2_ASAP7_75t_L g11329 ( 
.A(n_10799),
.B(n_8987),
.Y(n_11329)
);

NAND2xp5_ASAP7_75t_L g11330 ( 
.A(n_10725),
.B(n_8987),
.Y(n_11330)
);

NAND2xp5_ASAP7_75t_L g11331 ( 
.A(n_10725),
.B(n_8999),
.Y(n_11331)
);

OAI21xp5_ASAP7_75t_SL g11332 ( 
.A1(n_10998),
.A2(n_7307),
.B(n_9477),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_L g11333 ( 
.A(n_10859),
.B(n_8999),
.Y(n_11333)
);

AND2x2_ASAP7_75t_L g11334 ( 
.A(n_10528),
.B(n_9001),
.Y(n_11334)
);

NAND2xp5_ASAP7_75t_L g11335 ( 
.A(n_10860),
.B(n_10873),
.Y(n_11335)
);

NAND2xp5_ASAP7_75t_L g11336 ( 
.A(n_10886),
.B(n_9001),
.Y(n_11336)
);

AOI22xp33_ASAP7_75t_L g11337 ( 
.A1(n_10933),
.A2(n_10902),
.B1(n_10931),
.B2(n_10900),
.Y(n_11337)
);

OAI21xp5_ASAP7_75t_L g11338 ( 
.A1(n_10969),
.A2(n_8537),
.B(n_8516),
.Y(n_11338)
);

AOI221xp5_ASAP7_75t_L g11339 ( 
.A1(n_10984),
.A2(n_9135),
.B1(n_9140),
.B2(n_9131),
.C(n_9130),
.Y(n_11339)
);

AOI221xp5_ASAP7_75t_L g11340 ( 
.A1(n_10537),
.A2(n_9150),
.B1(n_9159),
.B2(n_9149),
.C(n_9140),
.Y(n_11340)
);

OAI221xp5_ASAP7_75t_SL g11341 ( 
.A1(n_11083),
.A2(n_9492),
.B1(n_9523),
.B2(n_9507),
.C(n_9477),
.Y(n_11341)
);

NAND2xp5_ASAP7_75t_L g11342 ( 
.A(n_10889),
.B(n_9008),
.Y(n_11342)
);

AND2x2_ASAP7_75t_L g11343 ( 
.A(n_10539),
.B(n_10933),
.Y(n_11343)
);

NAND2xp5_ASAP7_75t_L g11344 ( 
.A(n_10891),
.B(n_9008),
.Y(n_11344)
);

AOI22xp33_ASAP7_75t_L g11345 ( 
.A1(n_10900),
.A2(n_7951),
.B1(n_8312),
.B2(n_8356),
.Y(n_11345)
);

OAI221xp5_ASAP7_75t_L g11346 ( 
.A1(n_10998),
.A2(n_9523),
.B1(n_9533),
.B2(n_9507),
.C(n_9492),
.Y(n_11346)
);

AND2x2_ASAP7_75t_L g11347 ( 
.A(n_10878),
.B(n_9010),
.Y(n_11347)
);

OAI22xp5_ASAP7_75t_L g11348 ( 
.A1(n_10647),
.A2(n_11065),
.B1(n_10586),
.B2(n_10813),
.Y(n_11348)
);

OAI22xp5_ASAP7_75t_L g11349 ( 
.A1(n_10647),
.A2(n_10586),
.B1(n_10813),
.B2(n_11093),
.Y(n_11349)
);

NAND2xp5_ASAP7_75t_L g11350 ( 
.A(n_10892),
.B(n_9010),
.Y(n_11350)
);

AND2x2_ASAP7_75t_L g11351 ( 
.A(n_10691),
.B(n_9011),
.Y(n_11351)
);

NAND2xp5_ASAP7_75t_L g11352 ( 
.A(n_10894),
.B(n_9011),
.Y(n_11352)
);

OAI221xp5_ASAP7_75t_L g11353 ( 
.A1(n_11083),
.A2(n_9569),
.B1(n_9587),
.B2(n_9533),
.C(n_9523),
.Y(n_11353)
);

OAI21xp33_ASAP7_75t_L g11354 ( 
.A1(n_10829),
.A2(n_7563),
.B(n_10293),
.Y(n_11354)
);

NAND2xp5_ASAP7_75t_L g11355 ( 
.A(n_10897),
.B(n_9013),
.Y(n_11355)
);

NOR3xp33_ASAP7_75t_SL g11356 ( 
.A(n_10601),
.B(n_7504),
.C(n_7413),
.Y(n_11356)
);

NAND2xp5_ASAP7_75t_SL g11357 ( 
.A(n_10615),
.B(n_7109),
.Y(n_11357)
);

NAND3xp33_ASAP7_75t_L g11358 ( 
.A(n_10704),
.B(n_9680),
.C(n_7951),
.Y(n_11358)
);

AND2x2_ASAP7_75t_L g11359 ( 
.A(n_10911),
.B(n_9013),
.Y(n_11359)
);

NAND2xp5_ASAP7_75t_L g11360 ( 
.A(n_10899),
.B(n_9680),
.Y(n_11360)
);

NAND2xp5_ASAP7_75t_L g11361 ( 
.A(n_10901),
.B(n_9680),
.Y(n_11361)
);

NAND2xp5_ASAP7_75t_L g11362 ( 
.A(n_10904),
.B(n_8628),
.Y(n_11362)
);

AND2x2_ASAP7_75t_L g11363 ( 
.A(n_10695),
.B(n_8629),
.Y(n_11363)
);

NAND3xp33_ASAP7_75t_L g11364 ( 
.A(n_11107),
.B(n_11093),
.C(n_11067),
.Y(n_11364)
);

NOR3xp33_ASAP7_75t_SL g11365 ( 
.A(n_10601),
.B(n_7787),
.C(n_7669),
.Y(n_11365)
);

NAND2xp5_ASAP7_75t_L g11366 ( 
.A(n_10910),
.B(n_8629),
.Y(n_11366)
);

NOR2xp33_ASAP7_75t_SL g11367 ( 
.A(n_10505),
.B(n_7040),
.Y(n_11367)
);

AND2x2_ASAP7_75t_L g11368 ( 
.A(n_10697),
.B(n_8629),
.Y(n_11368)
);

OAI22xp5_ASAP7_75t_L g11369 ( 
.A1(n_10493),
.A2(n_7617),
.B1(n_7624),
.B2(n_7594),
.Y(n_11369)
);

AOI221xp5_ASAP7_75t_L g11370 ( 
.A1(n_11067),
.A2(n_9159),
.B1(n_9160),
.B2(n_9150),
.C(n_9149),
.Y(n_11370)
);

NAND2xp5_ASAP7_75t_L g11371 ( 
.A(n_10916),
.B(n_8650),
.Y(n_11371)
);

OAI21xp5_ASAP7_75t_SL g11372 ( 
.A1(n_10908),
.A2(n_9569),
.B(n_9533),
.Y(n_11372)
);

OAI221xp5_ASAP7_75t_L g11373 ( 
.A1(n_10607),
.A2(n_9640),
.B1(n_9665),
.B2(n_9587),
.C(n_9569),
.Y(n_11373)
);

OAI22xp5_ASAP7_75t_L g11374 ( 
.A1(n_10493),
.A2(n_7617),
.B1(n_7624),
.B2(n_7594),
.Y(n_11374)
);

NAND2xp5_ASAP7_75t_SL g11375 ( 
.A(n_10615),
.B(n_7109),
.Y(n_11375)
);

AND2x2_ASAP7_75t_L g11376 ( 
.A(n_10698),
.B(n_8650),
.Y(n_11376)
);

NAND2xp5_ASAP7_75t_L g11377 ( 
.A(n_10917),
.B(n_8650),
.Y(n_11377)
);

NAND2xp5_ASAP7_75t_L g11378 ( 
.A(n_10918),
.B(n_8651),
.Y(n_11378)
);

AND2x2_ASAP7_75t_L g11379 ( 
.A(n_10703),
.B(n_8651),
.Y(n_11379)
);

AND2x2_ASAP7_75t_L g11380 ( 
.A(n_10709),
.B(n_8651),
.Y(n_11380)
);

NAND2xp5_ASAP7_75t_L g11381 ( 
.A(n_10920),
.B(n_10930),
.Y(n_11381)
);

NAND2xp5_ASAP7_75t_SL g11382 ( 
.A(n_10672),
.B(n_7109),
.Y(n_11382)
);

NAND2xp5_ASAP7_75t_L g11383 ( 
.A(n_10932),
.B(n_8669),
.Y(n_11383)
);

AND2x2_ASAP7_75t_L g11384 ( 
.A(n_10902),
.B(n_8669),
.Y(n_11384)
);

AND2x2_ASAP7_75t_SL g11385 ( 
.A(n_10963),
.B(n_6648),
.Y(n_11385)
);

NAND2xp5_ASAP7_75t_L g11386 ( 
.A(n_10936),
.B(n_8669),
.Y(n_11386)
);

NAND2xp5_ASAP7_75t_L g11387 ( 
.A(n_10937),
.B(n_10940),
.Y(n_11387)
);

OAI22xp5_ASAP7_75t_L g11388 ( 
.A1(n_11107),
.A2(n_7617),
.B1(n_7624),
.B2(n_7594),
.Y(n_11388)
);

NOR3xp33_ASAP7_75t_L g11389 ( 
.A(n_10664),
.B(n_9338),
.C(n_9324),
.Y(n_11389)
);

AOI221xp5_ASAP7_75t_L g11390 ( 
.A1(n_10762),
.A2(n_10845),
.B1(n_10820),
.B2(n_11102),
.C(n_11101),
.Y(n_11390)
);

NAND3xp33_ASAP7_75t_L g11391 ( 
.A(n_11104),
.B(n_7951),
.C(n_9567),
.Y(n_11391)
);

NAND3xp33_ASAP7_75t_L g11392 ( 
.A(n_10672),
.B(n_9621),
.C(n_9567),
.Y(n_11392)
);

AND2x2_ASAP7_75t_L g11393 ( 
.A(n_10931),
.B(n_10655),
.Y(n_11393)
);

AND2x2_ASAP7_75t_L g11394 ( 
.A(n_10942),
.B(n_8782),
.Y(n_11394)
);

OAI221xp5_ASAP7_75t_L g11395 ( 
.A1(n_11017),
.A2(n_9665),
.B1(n_9640),
.B2(n_9587),
.C(n_9357),
.Y(n_11395)
);

OAI22xp5_ASAP7_75t_L g11396 ( 
.A1(n_10533),
.A2(n_7624),
.B1(n_7641),
.B2(n_7617),
.Y(n_11396)
);

NAND3xp33_ASAP7_75t_L g11397 ( 
.A(n_10672),
.B(n_11118),
.C(n_10947),
.Y(n_11397)
);

NAND2xp5_ASAP7_75t_L g11398 ( 
.A(n_10941),
.B(n_8782),
.Y(n_11398)
);

NOR2xp33_ASAP7_75t_L g11399 ( 
.A(n_10498),
.B(n_7040),
.Y(n_11399)
);

AND2x2_ASAP7_75t_L g11400 ( 
.A(n_10963),
.B(n_10913),
.Y(n_11400)
);

OAI21xp5_ASAP7_75t_SL g11401 ( 
.A1(n_10908),
.A2(n_9665),
.B(n_9640),
.Y(n_11401)
);

AND2x2_ASAP7_75t_L g11402 ( 
.A(n_10928),
.B(n_8782),
.Y(n_11402)
);

AND2x2_ASAP7_75t_L g11403 ( 
.A(n_10882),
.B(n_8791),
.Y(n_11403)
);

AOI221xp5_ASAP7_75t_L g11404 ( 
.A1(n_10762),
.A2(n_9167),
.B1(n_9172),
.B2(n_9165),
.C(n_9160),
.Y(n_11404)
);

NAND2xp5_ASAP7_75t_L g11405 ( 
.A(n_10945),
.B(n_8791),
.Y(n_11405)
);

NAND3xp33_ASAP7_75t_L g11406 ( 
.A(n_10672),
.B(n_11118),
.C(n_10947),
.Y(n_11406)
);

AOI22xp33_ASAP7_75t_SL g11407 ( 
.A1(n_11115),
.A2(n_8312),
.B1(n_6711),
.B2(n_6840),
.Y(n_11407)
);

NAND3xp33_ASAP7_75t_L g11408 ( 
.A(n_10772),
.B(n_9621),
.C(n_9567),
.Y(n_11408)
);

AND2x2_ASAP7_75t_L g11409 ( 
.A(n_10890),
.B(n_8791),
.Y(n_11409)
);

NAND3xp33_ASAP7_75t_L g11410 ( 
.A(n_10772),
.B(n_9621),
.C(n_9567),
.Y(n_11410)
);

NAND2xp5_ASAP7_75t_L g11411 ( 
.A(n_10956),
.B(n_9165),
.Y(n_11411)
);

AND2x2_ASAP7_75t_L g11412 ( 
.A(n_10896),
.B(n_9280),
.Y(n_11412)
);

HB1xp67_ASAP7_75t_L g11413 ( 
.A(n_11029),
.Y(n_11413)
);

AND2x2_ASAP7_75t_L g11414 ( 
.A(n_10685),
.B(n_9280),
.Y(n_11414)
);

OAI21xp5_ASAP7_75t_SL g11415 ( 
.A1(n_10869),
.A2(n_9338),
.B(n_9324),
.Y(n_11415)
);

NAND4xp25_ASAP7_75t_L g11416 ( 
.A(n_11077),
.B(n_7614),
.C(n_7540),
.D(n_7167),
.Y(n_11416)
);

AND2x2_ASAP7_75t_SL g11417 ( 
.A(n_10532),
.B(n_7230),
.Y(n_11417)
);

NAND2xp5_ASAP7_75t_L g11418 ( 
.A(n_10957),
.B(n_9167),
.Y(n_11418)
);

AOI22xp33_ASAP7_75t_L g11419 ( 
.A1(n_11073),
.A2(n_8312),
.B1(n_8356),
.B2(n_8207),
.Y(n_11419)
);

OAI21xp5_ASAP7_75t_SL g11420 ( 
.A1(n_10869),
.A2(n_9380),
.B(n_9357),
.Y(n_11420)
);

NOR3xp33_ASAP7_75t_L g11421 ( 
.A(n_10797),
.B(n_9380),
.C(n_9357),
.Y(n_11421)
);

AOI22xp5_ASAP7_75t_L g11422 ( 
.A1(n_10472),
.A2(n_6704),
.B1(n_6840),
.B2(n_6711),
.Y(n_11422)
);

OAI21xp33_ASAP7_75t_L g11423 ( 
.A1(n_10954),
.A2(n_7563),
.B(n_6950),
.Y(n_11423)
);

AND2x2_ASAP7_75t_L g11424 ( 
.A(n_10649),
.B(n_9292),
.Y(n_11424)
);

AND2x2_ASAP7_75t_L g11425 ( 
.A(n_10650),
.B(n_9292),
.Y(n_11425)
);

AND2x2_ASAP7_75t_L g11426 ( 
.A(n_10652),
.B(n_10546),
.Y(n_11426)
);

AND2x2_ASAP7_75t_L g11427 ( 
.A(n_10553),
.B(n_9298),
.Y(n_11427)
);

NAND3xp33_ASAP7_75t_L g11428 ( 
.A(n_10820),
.B(n_9621),
.C(n_9028),
.Y(n_11428)
);

NAND2xp5_ASAP7_75t_L g11429 ( 
.A(n_10958),
.B(n_10845),
.Y(n_11429)
);

NAND3xp33_ASAP7_75t_L g11430 ( 
.A(n_10960),
.B(n_9028),
.C(n_9173),
.Y(n_11430)
);

NOR3xp33_ASAP7_75t_L g11431 ( 
.A(n_10797),
.B(n_9389),
.C(n_9380),
.Y(n_11431)
);

NAND2xp5_ASAP7_75t_L g11432 ( 
.A(n_10839),
.B(n_9172),
.Y(n_11432)
);

NAND2xp5_ASAP7_75t_L g11433 ( 
.A(n_10843),
.B(n_9174),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_10716),
.B(n_9174),
.Y(n_11434)
);

NOR3xp33_ASAP7_75t_L g11435 ( 
.A(n_10835),
.B(n_9398),
.C(n_9389),
.Y(n_11435)
);

NAND2xp5_ASAP7_75t_L g11436 ( 
.A(n_10718),
.B(n_9178),
.Y(n_11436)
);

AND2x2_ASAP7_75t_L g11437 ( 
.A(n_10555),
.B(n_9298),
.Y(n_11437)
);

AOI221xp5_ASAP7_75t_L g11438 ( 
.A1(n_10841),
.A2(n_10559),
.B1(n_11092),
.B2(n_11097),
.C(n_11089),
.Y(n_11438)
);

NAND3xp33_ASAP7_75t_L g11439 ( 
.A(n_10960),
.B(n_9028),
.C(n_9173),
.Y(n_11439)
);

AND2x2_ASAP7_75t_L g11440 ( 
.A(n_10561),
.B(n_9299),
.Y(n_11440)
);

NAND3xp33_ASAP7_75t_L g11441 ( 
.A(n_10876),
.B(n_11058),
.C(n_11054),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_L g11442 ( 
.A(n_10837),
.B(n_10679),
.Y(n_11442)
);

NAND3xp33_ASAP7_75t_L g11443 ( 
.A(n_10876),
.B(n_9028),
.C(n_9173),
.Y(n_11443)
);

AND2x2_ASAP7_75t_L g11444 ( 
.A(n_10569),
.B(n_9299),
.Y(n_11444)
);

NAND2xp5_ASAP7_75t_L g11445 ( 
.A(n_10680),
.B(n_9178),
.Y(n_11445)
);

NOR2xp33_ASAP7_75t_L g11446 ( 
.A(n_10498),
.B(n_7056),
.Y(n_11446)
);

AND2x2_ASAP7_75t_SL g11447 ( 
.A(n_10532),
.B(n_7230),
.Y(n_11447)
);

NAND2xp5_ASAP7_75t_L g11448 ( 
.A(n_11005),
.B(n_9179),
.Y(n_11448)
);

NOR3xp33_ASAP7_75t_L g11449 ( 
.A(n_10835),
.B(n_9398),
.C(n_9389),
.Y(n_11449)
);

NAND2xp5_ASAP7_75t_L g11450 ( 
.A(n_11008),
.B(n_9179),
.Y(n_11450)
);

INVx1_ASAP7_75t_L g11451 ( 
.A(n_10470),
.Y(n_11451)
);

OR2x2_ASAP7_75t_L g11452 ( 
.A(n_10588),
.B(n_9181),
.Y(n_11452)
);

NAND2xp5_ASAP7_75t_L g11453 ( 
.A(n_11010),
.B(n_11011),
.Y(n_11453)
);

NAND2xp5_ASAP7_75t_L g11454 ( 
.A(n_11013),
.B(n_9181),
.Y(n_11454)
);

NAND2xp5_ASAP7_75t_L g11455 ( 
.A(n_11014),
.B(n_9184),
.Y(n_11455)
);

NAND2xp5_ASAP7_75t_L g11456 ( 
.A(n_11050),
.B(n_9184),
.Y(n_11456)
);

NAND2xp5_ASAP7_75t_L g11457 ( 
.A(n_11090),
.B(n_9188),
.Y(n_11457)
);

NAND3xp33_ASAP7_75t_L g11458 ( 
.A(n_11063),
.B(n_11112),
.C(n_11109),
.Y(n_11458)
);

AND2x2_ASAP7_75t_L g11459 ( 
.A(n_10574),
.B(n_9316),
.Y(n_11459)
);

NAND2xp5_ASAP7_75t_L g11460 ( 
.A(n_11110),
.B(n_11111),
.Y(n_11460)
);

NAND4xp25_ASAP7_75t_L g11461 ( 
.A(n_11080),
.B(n_9422),
.C(n_9398),
.D(n_7147),
.Y(n_11461)
);

NAND2xp5_ASAP7_75t_L g11462 ( 
.A(n_10938),
.B(n_9188),
.Y(n_11462)
);

NAND2xp5_ASAP7_75t_L g11463 ( 
.A(n_11018),
.B(n_9191),
.Y(n_11463)
);

NAND3xp33_ASAP7_75t_L g11464 ( 
.A(n_11116),
.B(n_9173),
.C(n_9191),
.Y(n_11464)
);

NAND2xp5_ASAP7_75t_L g11465 ( 
.A(n_11027),
.B(n_9192),
.Y(n_11465)
);

INVx1_ASAP7_75t_L g11466 ( 
.A(n_10471),
.Y(n_11466)
);

NAND2xp5_ASAP7_75t_L g11467 ( 
.A(n_11119),
.B(n_9192),
.Y(n_11467)
);

OAI22xp5_ASAP7_75t_L g11468 ( 
.A1(n_10450),
.A2(n_7641),
.B1(n_7644),
.B2(n_7617),
.Y(n_11468)
);

NAND3xp33_ASAP7_75t_L g11469 ( 
.A(n_10623),
.B(n_9201),
.C(n_9195),
.Y(n_11469)
);

NAND2xp5_ASAP7_75t_L g11470 ( 
.A(n_11132),
.B(n_9195),
.Y(n_11470)
);

NAND2xp5_ASAP7_75t_SL g11471 ( 
.A(n_10641),
.B(n_7826),
.Y(n_11471)
);

OAI21xp5_ASAP7_75t_L g11472 ( 
.A1(n_10461),
.A2(n_8537),
.B(n_8516),
.Y(n_11472)
);

OAI22xp33_ASAP7_75t_L g11473 ( 
.A1(n_10591),
.A2(n_7149),
.B1(n_7284),
.B2(n_7083),
.Y(n_11473)
);

NAND2xp5_ASAP7_75t_L g11474 ( 
.A(n_11069),
.B(n_9201),
.Y(n_11474)
);

AOI21xp5_ASAP7_75t_SL g11475 ( 
.A1(n_10496),
.A2(n_8596),
.B(n_8516),
.Y(n_11475)
);

NAND2xp5_ASAP7_75t_L g11476 ( 
.A(n_11071),
.B(n_9208),
.Y(n_11476)
);

NAND2xp5_ASAP7_75t_L g11477 ( 
.A(n_11041),
.B(n_9208),
.Y(n_11477)
);

INVx2_ASAP7_75t_L g11478 ( 
.A(n_10604),
.Y(n_11478)
);

AOI22xp33_ASAP7_75t_L g11479 ( 
.A1(n_11070),
.A2(n_8356),
.B1(n_8207),
.B2(n_8241),
.Y(n_11479)
);

AND2x2_ASAP7_75t_L g11480 ( 
.A(n_10575),
.B(n_9316),
.Y(n_11480)
);

OAI22xp5_ASAP7_75t_L g11481 ( 
.A1(n_10469),
.A2(n_7644),
.B1(n_7664),
.B2(n_7641),
.Y(n_11481)
);

NAND2xp5_ASAP7_75t_L g11482 ( 
.A(n_11041),
.B(n_11088),
.Y(n_11482)
);

OAI221xp5_ASAP7_75t_L g11483 ( 
.A1(n_10472),
.A2(n_9422),
.B1(n_8698),
.B2(n_8596),
.C(n_7895),
.Y(n_11483)
);

NAND2xp5_ASAP7_75t_L g11484 ( 
.A(n_11088),
.B(n_9212),
.Y(n_11484)
);

NAND2x1_ASAP7_75t_L g11485 ( 
.A(n_10465),
.B(n_10435),
.Y(n_11485)
);

NAND3xp33_ASAP7_75t_L g11486 ( 
.A(n_10623),
.B(n_9217),
.C(n_9212),
.Y(n_11486)
);

AOI21xp5_ASAP7_75t_SL g11487 ( 
.A1(n_10596),
.A2(n_8698),
.B(n_8596),
.Y(n_11487)
);

AND2x2_ASAP7_75t_L g11488 ( 
.A(n_10584),
.B(n_9322),
.Y(n_11488)
);

NAND3xp33_ASAP7_75t_L g11489 ( 
.A(n_10712),
.B(n_9220),
.C(n_9217),
.Y(n_11489)
);

NOR3xp33_ASAP7_75t_L g11490 ( 
.A(n_11081),
.B(n_10712),
.C(n_10699),
.Y(n_11490)
);

NAND3xp33_ASAP7_75t_L g11491 ( 
.A(n_11007),
.B(n_9234),
.C(n_9220),
.Y(n_11491)
);

OAI21xp33_ASAP7_75t_L g11492 ( 
.A1(n_11094),
.A2(n_6945),
.B(n_7110),
.Y(n_11492)
);

NOR2xp33_ASAP7_75t_L g11493 ( 
.A(n_10598),
.B(n_10905),
.Y(n_11493)
);

AND2x2_ASAP7_75t_L g11494 ( 
.A(n_10773),
.B(n_9322),
.Y(n_11494)
);

AND2x2_ASAP7_75t_L g11495 ( 
.A(n_10594),
.B(n_10605),
.Y(n_11495)
);

NAND2xp5_ASAP7_75t_L g11496 ( 
.A(n_10557),
.B(n_9234),
.Y(n_11496)
);

OAI22xp33_ASAP7_75t_L g11497 ( 
.A1(n_10591),
.A2(n_7284),
.B1(n_7438),
.B2(n_7149),
.Y(n_11497)
);

OAI21xp5_ASAP7_75t_SL g11498 ( 
.A1(n_10793),
.A2(n_9422),
.B(n_6902),
.Y(n_11498)
);

AND2x2_ASAP7_75t_L g11499 ( 
.A(n_10665),
.B(n_9327),
.Y(n_11499)
);

AOI221xp5_ASAP7_75t_L g11500 ( 
.A1(n_10559),
.A2(n_9248),
.B1(n_9252),
.B2(n_9241),
.C(n_9237),
.Y(n_11500)
);

INVx1_ASAP7_75t_L g11501 ( 
.A(n_10475),
.Y(n_11501)
);

NAND2xp5_ASAP7_75t_L g11502 ( 
.A(n_11033),
.B(n_9237),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_10608),
.B(n_9327),
.Y(n_11503)
);

NAND2xp5_ASAP7_75t_L g11504 ( 
.A(n_11044),
.B(n_9241),
.Y(n_11504)
);

NAND3xp33_ASAP7_75t_L g11505 ( 
.A(n_11007),
.B(n_9252),
.C(n_9248),
.Y(n_11505)
);

AND2x2_ASAP7_75t_L g11506 ( 
.A(n_10609),
.B(n_9336),
.Y(n_11506)
);

AOI22xp33_ASAP7_75t_SL g11507 ( 
.A1(n_10884),
.A2(n_10499),
.B1(n_11087),
.B2(n_11079),
.Y(n_11507)
);

OR2x6_ASAP7_75t_SL g11508 ( 
.A(n_10905),
.B(n_6995),
.Y(n_11508)
);

NAND3xp33_ASAP7_75t_L g11509 ( 
.A(n_11114),
.B(n_9257),
.C(n_9256),
.Y(n_11509)
);

AND2x2_ASAP7_75t_L g11510 ( 
.A(n_10612),
.B(n_10613),
.Y(n_11510)
);

OAI22xp5_ASAP7_75t_L g11511 ( 
.A1(n_10465),
.A2(n_7644),
.B1(n_7664),
.B2(n_7641),
.Y(n_11511)
);

NAND2xp5_ASAP7_75t_L g11512 ( 
.A(n_11046),
.B(n_9256),
.Y(n_11512)
);

AND2x2_ASAP7_75t_L g11513 ( 
.A(n_10616),
.B(n_9336),
.Y(n_11513)
);

AOI221xp5_ASAP7_75t_L g11514 ( 
.A1(n_10848),
.A2(n_10856),
.B1(n_10850),
.B2(n_10503),
.C(n_10531),
.Y(n_11514)
);

NAND2xp5_ASAP7_75t_SL g11515 ( 
.A(n_10641),
.B(n_7826),
.Y(n_11515)
);

NAND2xp5_ASAP7_75t_L g11516 ( 
.A(n_11098),
.B(n_9257),
.Y(n_11516)
);

OAI21xp5_ASAP7_75t_SL g11517 ( 
.A1(n_10793),
.A2(n_7176),
.B(n_7526),
.Y(n_11517)
);

NOR3xp33_ASAP7_75t_L g11518 ( 
.A(n_10495),
.B(n_10261),
.C(n_10012),
.Y(n_11518)
);

AOI21xp33_ASAP7_75t_L g11519 ( 
.A1(n_10499),
.A2(n_8698),
.B(n_9258),
.Y(n_11519)
);

NAND2xp5_ASAP7_75t_L g11520 ( 
.A(n_11066),
.B(n_9258),
.Y(n_11520)
);

NAND2xp5_ASAP7_75t_SL g11521 ( 
.A(n_10669),
.B(n_7826),
.Y(n_11521)
);

AOI21xp5_ASAP7_75t_SL g11522 ( 
.A1(n_11056),
.A2(n_10192),
.B(n_10435),
.Y(n_11522)
);

OAI22xp5_ASAP7_75t_L g11523 ( 
.A1(n_10705),
.A2(n_7644),
.B1(n_7664),
.B2(n_7641),
.Y(n_11523)
);

AND2x2_ASAP7_75t_L g11524 ( 
.A(n_10619),
.B(n_9342),
.Y(n_11524)
);

AND2x2_ASAP7_75t_L g11525 ( 
.A(n_10621),
.B(n_9342),
.Y(n_11525)
);

NAND2xp5_ASAP7_75t_L g11526 ( 
.A(n_11084),
.B(n_9261),
.Y(n_11526)
);

NAND2xp5_ASAP7_75t_L g11527 ( 
.A(n_10868),
.B(n_9261),
.Y(n_11527)
);

NOR2xp33_ASAP7_75t_R g11528 ( 
.A(n_10598),
.B(n_7056),
.Y(n_11528)
);

NAND2xp5_ASAP7_75t_L g11529 ( 
.A(n_10883),
.B(n_9262),
.Y(n_11529)
);

NAND2xp5_ASAP7_75t_L g11530 ( 
.A(n_10761),
.B(n_9262),
.Y(n_11530)
);

AOI22xp5_ASAP7_75t_L g11531 ( 
.A1(n_10548),
.A2(n_6704),
.B1(n_6954),
.B2(n_6878),
.Y(n_11531)
);

NOR3xp33_ASAP7_75t_L g11532 ( 
.A(n_10657),
.B(n_9987),
.C(n_10071),
.Y(n_11532)
);

AND2x2_ASAP7_75t_L g11533 ( 
.A(n_10633),
.B(n_9353),
.Y(n_11533)
);

OAI22xp5_ASAP7_75t_L g11534 ( 
.A1(n_10707),
.A2(n_10710),
.B1(n_10715),
.B2(n_10628),
.Y(n_11534)
);

AND2x2_ASAP7_75t_L g11535 ( 
.A(n_10639),
.B(n_9353),
.Y(n_11535)
);

NAND3xp33_ASAP7_75t_L g11536 ( 
.A(n_11114),
.B(n_10915),
.C(n_10875),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_10767),
.B(n_10771),
.Y(n_11537)
);

NAND2xp5_ASAP7_75t_SL g11538 ( 
.A(n_10669),
.B(n_7826),
.Y(n_11538)
);

NOR2xp33_ASAP7_75t_SL g11539 ( 
.A(n_10689),
.B(n_7071),
.Y(n_11539)
);

NAND2xp5_ASAP7_75t_L g11540 ( 
.A(n_10776),
.B(n_9263),
.Y(n_11540)
);

NAND2xp5_ASAP7_75t_L g11541 ( 
.A(n_10777),
.B(n_9263),
.Y(n_11541)
);

NAND2xp5_ASAP7_75t_L g11542 ( 
.A(n_10781),
.B(n_9264),
.Y(n_11542)
);

NAND2xp5_ASAP7_75t_L g11543 ( 
.A(n_10782),
.B(n_9264),
.Y(n_11543)
);

OA211x2_ASAP7_75t_L g11544 ( 
.A1(n_11037),
.A2(n_6995),
.B(n_7062),
.C(n_9915),
.Y(n_11544)
);

NAND3xp33_ASAP7_75t_L g11545 ( 
.A(n_10875),
.B(n_9266),
.C(n_9265),
.Y(n_11545)
);

NAND2xp5_ASAP7_75t_L g11546 ( 
.A(n_10783),
.B(n_9265),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_L g11547 ( 
.A(n_10788),
.B(n_9266),
.Y(n_11547)
);

NAND2xp5_ASAP7_75t_L g11548 ( 
.A(n_10790),
.B(n_9267),
.Y(n_11548)
);

AND2x2_ASAP7_75t_L g11549 ( 
.A(n_10871),
.B(n_9363),
.Y(n_11549)
);

OA21x2_ASAP7_75t_L g11550 ( 
.A1(n_10948),
.A2(n_10129),
.B(n_9275),
.Y(n_11550)
);

NAND3xp33_ASAP7_75t_L g11551 ( 
.A(n_10915),
.B(n_9275),
.C(n_9267),
.Y(n_11551)
);

NAND2xp5_ASAP7_75t_L g11552 ( 
.A(n_10796),
.B(n_9281),
.Y(n_11552)
);

INVx2_ASAP7_75t_SL g11553 ( 
.A(n_10807),
.Y(n_11553)
);

AND2x2_ASAP7_75t_L g11554 ( 
.A(n_10874),
.B(n_9363),
.Y(n_11554)
);

NAND2xp5_ASAP7_75t_L g11555 ( 
.A(n_10801),
.B(n_9281),
.Y(n_11555)
);

AND2x2_ASAP7_75t_L g11556 ( 
.A(n_10648),
.B(n_10501),
.Y(n_11556)
);

OAI21xp33_ASAP7_75t_L g11557 ( 
.A1(n_11100),
.A2(n_7293),
.B(n_7260),
.Y(n_11557)
);

AND2x2_ASAP7_75t_SL g11558 ( 
.A(n_10862),
.B(n_7230),
.Y(n_11558)
);

AND2x2_ASAP7_75t_L g11559 ( 
.A(n_10511),
.B(n_9377),
.Y(n_11559)
);

NOR2xp33_ASAP7_75t_SL g11560 ( 
.A(n_10683),
.B(n_7071),
.Y(n_11560)
);

NAND4xp25_ASAP7_75t_L g11561 ( 
.A(n_11106),
.B(n_11072),
.C(n_11086),
.D(n_10673),
.Y(n_11561)
);

NAND3xp33_ASAP7_75t_L g11562 ( 
.A(n_10919),
.B(n_7928),
.C(n_9980),
.Y(n_11562)
);

NAND3xp33_ASAP7_75t_L g11563 ( 
.A(n_10919),
.B(n_7928),
.C(n_9980),
.Y(n_11563)
);

OAI22xp5_ASAP7_75t_L g11564 ( 
.A1(n_11079),
.A2(n_7664),
.B1(n_7674),
.B2(n_7644),
.Y(n_11564)
);

NAND3xp33_ASAP7_75t_L g11565 ( 
.A(n_10987),
.B(n_7928),
.C(n_9989),
.Y(n_11565)
);

NAND2xp5_ASAP7_75t_L g11566 ( 
.A(n_10802),
.B(n_8885),
.Y(n_11566)
);

AOI22xp5_ASAP7_75t_L g11567 ( 
.A1(n_11087),
.A2(n_11113),
.B1(n_11123),
.B2(n_10722),
.Y(n_11567)
);

OAI21xp5_ASAP7_75t_SL g11568 ( 
.A1(n_11113),
.A2(n_10923),
.B(n_10862),
.Y(n_11568)
);

AOI22xp5_ASAP7_75t_L g11569 ( 
.A1(n_10721),
.A2(n_6878),
.B1(n_6954),
.B2(n_7664),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_L g11570 ( 
.A(n_10809),
.B(n_8892),
.Y(n_11570)
);

NAND2xp5_ASAP7_75t_L g11571 ( 
.A(n_11030),
.B(n_8892),
.Y(n_11571)
);

NAND2xp5_ASAP7_75t_SL g11572 ( 
.A(n_10872),
.B(n_7826),
.Y(n_11572)
);

AND2x2_ASAP7_75t_SL g11573 ( 
.A(n_10923),
.B(n_7230),
.Y(n_11573)
);

OAI21xp33_ASAP7_75t_L g11574 ( 
.A1(n_10951),
.A2(n_11128),
.B(n_11130),
.Y(n_11574)
);

NOR3xp33_ASAP7_75t_L g11575 ( 
.A(n_10684),
.B(n_7250),
.C(n_7237),
.Y(n_11575)
);

AOI221xp5_ASAP7_75t_L g11576 ( 
.A1(n_10502),
.A2(n_7099),
.B1(n_7075),
.B2(n_7189),
.C(n_7065),
.Y(n_11576)
);

OA211x2_ASAP7_75t_L g11577 ( 
.A1(n_11037),
.A2(n_11131),
.B(n_11121),
.C(n_10552),
.Y(n_11577)
);

NAND2xp5_ASAP7_75t_L g11578 ( 
.A(n_11030),
.B(n_11032),
.Y(n_11578)
);

AND2x2_ASAP7_75t_L g11579 ( 
.A(n_10512),
.B(n_9377),
.Y(n_11579)
);

OAI221xp5_ASAP7_75t_L g11580 ( 
.A1(n_10673),
.A2(n_7895),
.B1(n_8681),
.B2(n_8702),
.C(n_8663),
.Y(n_11580)
);

AND2x2_ASAP7_75t_SL g11581 ( 
.A(n_10719),
.B(n_7240),
.Y(n_11581)
);

NAND2x1_ASAP7_75t_L g11582 ( 
.A(n_10770),
.B(n_10192),
.Y(n_11582)
);

AND2x2_ASAP7_75t_L g11583 ( 
.A(n_10514),
.B(n_9383),
.Y(n_11583)
);

NAND2xp5_ASAP7_75t_L g11584 ( 
.A(n_11032),
.B(n_8895),
.Y(n_11584)
);

AND2x2_ASAP7_75t_L g11585 ( 
.A(n_10866),
.B(n_9383),
.Y(n_11585)
);

INVx2_ASAP7_75t_L g11586 ( 
.A(n_10534),
.Y(n_11586)
);

OA21x2_ASAP7_75t_L g11587 ( 
.A1(n_10948),
.A2(n_9078),
.B(n_9075),
.Y(n_11587)
);

OAI21xp33_ASAP7_75t_L g11588 ( 
.A1(n_11129),
.A2(n_7293),
.B(n_7260),
.Y(n_11588)
);

NAND2xp5_ASAP7_75t_L g11589 ( 
.A(n_11040),
.B(n_8895),
.Y(n_11589)
);

NAND2xp5_ASAP7_75t_L g11590 ( 
.A(n_11040),
.B(n_8897),
.Y(n_11590)
);

HB1xp67_ASAP7_75t_L g11591 ( 
.A(n_11029),
.Y(n_11591)
);

OAI21xp5_ASAP7_75t_L g11592 ( 
.A1(n_11121),
.A2(n_7915),
.B(n_7896),
.Y(n_11592)
);

OAI22xp5_ASAP7_75t_L g11593 ( 
.A1(n_10562),
.A2(n_7683),
.B1(n_7725),
.B2(n_7674),
.Y(n_11593)
);

OAI21xp5_ASAP7_75t_SL g11594 ( 
.A1(n_10724),
.A2(n_7176),
.B(n_7010),
.Y(n_11594)
);

AND2x2_ASAP7_75t_L g11595 ( 
.A(n_10993),
.B(n_9416),
.Y(n_11595)
);

NAND2xp5_ASAP7_75t_L g11596 ( 
.A(n_11042),
.B(n_8897),
.Y(n_11596)
);

OAI22xp5_ASAP7_75t_L g11597 ( 
.A1(n_11099),
.A2(n_7683),
.B1(n_7725),
.B2(n_7674),
.Y(n_11597)
);

NAND2xp5_ASAP7_75t_L g11598 ( 
.A(n_11042),
.B(n_8898),
.Y(n_11598)
);

NAND2xp5_ASAP7_75t_L g11599 ( 
.A(n_10973),
.B(n_8898),
.Y(n_11599)
);

NAND2xp5_ASAP7_75t_L g11600 ( 
.A(n_10978),
.B(n_8899),
.Y(n_11600)
);

NAND3xp33_ASAP7_75t_L g11601 ( 
.A(n_10987),
.B(n_7928),
.C(n_9989),
.Y(n_11601)
);

OAI22xp5_ASAP7_75t_L g11602 ( 
.A1(n_10597),
.A2(n_7683),
.B1(n_7725),
.B2(n_7674),
.Y(n_11602)
);

AND2x2_ASAP7_75t_L g11603 ( 
.A(n_10750),
.B(n_9416),
.Y(n_11603)
);

OA21x2_ASAP7_75t_L g11604 ( 
.A1(n_10953),
.A2(n_9078),
.B(n_9075),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_L g11605 ( 
.A(n_10979),
.B(n_8899),
.Y(n_11605)
);

AND2x2_ASAP7_75t_L g11606 ( 
.A(n_10764),
.B(n_9418),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_10480),
.Y(n_11607)
);

OAI22xp5_ASAP7_75t_L g11608 ( 
.A1(n_10597),
.A2(n_7683),
.B1(n_7725),
.B2(n_7674),
.Y(n_11608)
);

NAND2xp5_ASAP7_75t_L g11609 ( 
.A(n_10980),
.B(n_10982),
.Y(n_11609)
);

NAND2xp5_ASAP7_75t_L g11610 ( 
.A(n_10999),
.B(n_8902),
.Y(n_11610)
);

AND2x2_ASAP7_75t_L g11611 ( 
.A(n_10766),
.B(n_9418),
.Y(n_11611)
);

AND2x2_ASAP7_75t_L g11612 ( 
.A(n_10570),
.B(n_9434),
.Y(n_11612)
);

NAND4xp25_ASAP7_75t_L g11613 ( 
.A(n_10946),
.B(n_7147),
.C(n_7535),
.D(n_7528),
.Y(n_11613)
);

OAI21xp5_ASAP7_75t_SL g11614 ( 
.A1(n_11026),
.A2(n_7010),
.B(n_6998),
.Y(n_11614)
);

OAI22xp33_ASAP7_75t_L g11615 ( 
.A1(n_10602),
.A2(n_7284),
.B1(n_7438),
.B2(n_7149),
.Y(n_11615)
);

OAI221xp5_ASAP7_75t_SL g11616 ( 
.A1(n_11131),
.A2(n_9941),
.B1(n_9915),
.B2(n_7067),
.C(n_7068),
.Y(n_11616)
);

NAND3xp33_ASAP7_75t_L g11617 ( 
.A(n_10786),
.B(n_10805),
.C(n_10872),
.Y(n_11617)
);

OAI21xp5_ASAP7_75t_SL g11618 ( 
.A1(n_11031),
.A2(n_6998),
.B(n_7389),
.Y(n_11618)
);

NAND2xp5_ASAP7_75t_L g11619 ( 
.A(n_10946),
.B(n_8902),
.Y(n_11619)
);

NAND2xp5_ASAP7_75t_L g11620 ( 
.A(n_11028),
.B(n_8905),
.Y(n_11620)
);

AND2x2_ASAP7_75t_L g11621 ( 
.A(n_10576),
.B(n_9434),
.Y(n_11621)
);

AOI22xp33_ASAP7_75t_SL g11622 ( 
.A1(n_10825),
.A2(n_8356),
.B1(n_7099),
.B2(n_7075),
.Y(n_11622)
);

AND2x2_ASAP7_75t_L g11623 ( 
.A(n_10622),
.B(n_9436),
.Y(n_11623)
);

AND2x2_ASAP7_75t_L g11624 ( 
.A(n_10626),
.B(n_9436),
.Y(n_11624)
);

OAI22xp5_ASAP7_75t_L g11625 ( 
.A1(n_10602),
.A2(n_7725),
.B1(n_7732),
.B2(n_7683),
.Y(n_11625)
);

NAND2xp5_ASAP7_75t_L g11626 ( 
.A(n_11028),
.B(n_8905),
.Y(n_11626)
);

OAI22xp5_ASAP7_75t_L g11627 ( 
.A1(n_10617),
.A2(n_10666),
.B1(n_10538),
.B2(n_10504),
.Y(n_11627)
);

OAI22xp5_ASAP7_75t_L g11628 ( 
.A1(n_10617),
.A2(n_7750),
.B1(n_7757),
.B2(n_7732),
.Y(n_11628)
);

INVx2_ASAP7_75t_L g11629 ( 
.A(n_10534),
.Y(n_11629)
);

NAND2xp5_ASAP7_75t_L g11630 ( 
.A(n_10921),
.B(n_8912),
.Y(n_11630)
);

NAND2xp5_ASAP7_75t_L g11631 ( 
.A(n_10921),
.B(n_8912),
.Y(n_11631)
);

OAI21xp5_ASAP7_75t_SL g11632 ( 
.A1(n_11035),
.A2(n_7389),
.B(n_7511),
.Y(n_11632)
);

NAND2xp5_ASAP7_75t_L g11633 ( 
.A(n_10921),
.B(n_8922),
.Y(n_11633)
);

OR2x2_ASAP7_75t_L g11634 ( 
.A(n_10729),
.B(n_8922),
.Y(n_11634)
);

AND2x2_ASAP7_75t_L g11635 ( 
.A(n_10627),
.B(n_9438),
.Y(n_11635)
);

NAND2xp5_ASAP7_75t_L g11636 ( 
.A(n_10991),
.B(n_8930),
.Y(n_11636)
);

NAND2xp5_ASAP7_75t_L g11637 ( 
.A(n_10991),
.B(n_8930),
.Y(n_11637)
);

NOR2xp33_ASAP7_75t_SL g11638 ( 
.A(n_10752),
.B(n_7071),
.Y(n_11638)
);

NAND2xp5_ASAP7_75t_L g11639 ( 
.A(n_10991),
.B(n_8931),
.Y(n_11639)
);

NAND2xp5_ASAP7_75t_L g11640 ( 
.A(n_10992),
.B(n_8931),
.Y(n_11640)
);

AND2x2_ASAP7_75t_L g11641 ( 
.A(n_10636),
.B(n_9438),
.Y(n_11641)
);

OAI21xp5_ASAP7_75t_SL g11642 ( 
.A1(n_11036),
.A2(n_11060),
.B(n_11055),
.Y(n_11642)
);

AND2x2_ASAP7_75t_L g11643 ( 
.A(n_10637),
.B(n_9439),
.Y(n_11643)
);

NOR2xp33_ASAP7_75t_L g11644 ( 
.A(n_10828),
.B(n_7134),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_10638),
.B(n_9439),
.Y(n_11645)
);

NAND2xp5_ASAP7_75t_L g11646 ( 
.A(n_10992),
.B(n_8936),
.Y(n_11646)
);

NAND3xp33_ASAP7_75t_L g11647 ( 
.A(n_10786),
.B(n_8356),
.C(n_7928),
.Y(n_11647)
);

AOI221xp5_ASAP7_75t_L g11648 ( 
.A1(n_10502),
.A2(n_7453),
.B1(n_7462),
.B2(n_7392),
.C(n_7321),
.Y(n_11648)
);

NAND3xp33_ASAP7_75t_L g11649 ( 
.A(n_10786),
.B(n_8038),
.C(n_7840),
.Y(n_11649)
);

AND2x2_ASAP7_75t_L g11650 ( 
.A(n_10644),
.B(n_9453),
.Y(n_11650)
);

AND2x2_ASAP7_75t_L g11651 ( 
.A(n_10658),
.B(n_9453),
.Y(n_11651)
);

NAND3xp33_ASAP7_75t_L g11652 ( 
.A(n_10786),
.B(n_8038),
.C(n_7840),
.Y(n_11652)
);

NAND2xp5_ASAP7_75t_L g11653 ( 
.A(n_10992),
.B(n_8936),
.Y(n_11653)
);

NAND2xp5_ASAP7_75t_L g11654 ( 
.A(n_11023),
.B(n_8937),
.Y(n_11654)
);

AOI22xp33_ASAP7_75t_L g11655 ( 
.A1(n_11062),
.A2(n_8207),
.B1(n_8241),
.B2(n_8191),
.Y(n_11655)
);

OAI21xp5_ASAP7_75t_SL g11656 ( 
.A1(n_10787),
.A2(n_7515),
.B(n_7429),
.Y(n_11656)
);

NAND2xp5_ASAP7_75t_L g11657 ( 
.A(n_11023),
.B(n_8937),
.Y(n_11657)
);

NAND2xp5_ASAP7_75t_L g11658 ( 
.A(n_11023),
.B(n_8944),
.Y(n_11658)
);

OAI22xp5_ASAP7_75t_L g11659 ( 
.A1(n_10507),
.A2(n_7750),
.B1(n_7757),
.B2(n_7732),
.Y(n_11659)
);

NAND4xp25_ASAP7_75t_L g11660 ( 
.A(n_10567),
.B(n_7147),
.C(n_7430),
.D(n_7114),
.Y(n_11660)
);

AND2x4_ASAP7_75t_L g11661 ( 
.A(n_10805),
.B(n_9465),
.Y(n_11661)
);

NAND2xp5_ASAP7_75t_L g11662 ( 
.A(n_10846),
.B(n_8944),
.Y(n_11662)
);

AOI22xp33_ASAP7_75t_L g11663 ( 
.A1(n_11051),
.A2(n_8207),
.B1(n_8241),
.B2(n_8191),
.Y(n_11663)
);

OA21x2_ASAP7_75t_L g11664 ( 
.A1(n_10953),
.A2(n_9081),
.B(n_9079),
.Y(n_11664)
);

NAND3xp33_ASAP7_75t_L g11665 ( 
.A(n_10805),
.B(n_8038),
.C(n_7840),
.Y(n_11665)
);

NAND3xp33_ASAP7_75t_L g11666 ( 
.A(n_10805),
.B(n_8038),
.C(n_7840),
.Y(n_11666)
);

AND2x2_ASAP7_75t_L g11667 ( 
.A(n_10674),
.B(n_9465),
.Y(n_11667)
);

NAND3xp33_ASAP7_75t_L g11668 ( 
.A(n_10872),
.B(n_8038),
.C(n_7840),
.Y(n_11668)
);

NAND2xp5_ASAP7_75t_L g11669 ( 
.A(n_10861),
.B(n_8946),
.Y(n_11669)
);

NAND2xp5_ASAP7_75t_SL g11670 ( 
.A(n_10474),
.B(n_7840),
.Y(n_11670)
);

AND2x2_ASAP7_75t_L g11671 ( 
.A(n_10818),
.B(n_9466),
.Y(n_11671)
);

NAND2xp5_ASAP7_75t_L g11672 ( 
.A(n_10863),
.B(n_8946),
.Y(n_11672)
);

OAI221xp5_ASAP7_75t_L g11673 ( 
.A1(n_11052),
.A2(n_7895),
.B1(n_8702),
.B2(n_8681),
.C(n_8038),
.Y(n_11673)
);

NAND2xp5_ASAP7_75t_L g11674 ( 
.A(n_10864),
.B(n_8956),
.Y(n_11674)
);

NAND3xp33_ASAP7_75t_SL g11675 ( 
.A(n_10513),
.B(n_8658),
.C(n_8646),
.Y(n_11675)
);

OAI22xp33_ASAP7_75t_SL g11676 ( 
.A1(n_10526),
.A2(n_8203),
.B1(n_8219),
.B2(n_8177),
.Y(n_11676)
);

NAND2xp5_ASAP7_75t_SL g11677 ( 
.A(n_10474),
.B(n_7840),
.Y(n_11677)
);

NAND2xp5_ASAP7_75t_SL g11678 ( 
.A(n_10735),
.B(n_8038),
.Y(n_11678)
);

OAI21xp33_ASAP7_75t_L g11679 ( 
.A1(n_10961),
.A2(n_7052),
.B(n_7392),
.Y(n_11679)
);

NAND2xp33_ASAP7_75t_R g11680 ( 
.A(n_10565),
.B(n_9827),
.Y(n_11680)
);

AND2x2_ASAP7_75t_L g11681 ( 
.A(n_10827),
.B(n_9466),
.Y(n_11681)
);

AOI22xp33_ASAP7_75t_L g11682 ( 
.A1(n_11075),
.A2(n_8207),
.B1(n_8241),
.B2(n_8191),
.Y(n_11682)
);

NAND2xp5_ASAP7_75t_L g11683 ( 
.A(n_10581),
.B(n_8956),
.Y(n_11683)
);

OAI21xp33_ASAP7_75t_L g11684 ( 
.A1(n_10962),
.A2(n_7462),
.B(n_7453),
.Y(n_11684)
);

OAI21xp33_ASAP7_75t_SL g11685 ( 
.A1(n_10544),
.A2(n_9486),
.B(n_9470),
.Y(n_11685)
);

NAND2xp5_ASAP7_75t_L g11686 ( 
.A(n_10581),
.B(n_8959),
.Y(n_11686)
);

AND2x2_ASAP7_75t_L g11687 ( 
.A(n_10831),
.B(n_9470),
.Y(n_11687)
);

NAND2xp5_ASAP7_75t_L g11688 ( 
.A(n_10581),
.B(n_8959),
.Y(n_11688)
);

AND2x2_ASAP7_75t_L g11689 ( 
.A(n_10852),
.B(n_10590),
.Y(n_11689)
);

NAND2xp5_ASAP7_75t_L g11690 ( 
.A(n_10589),
.B(n_8966),
.Y(n_11690)
);

OAI21xp33_ASAP7_75t_L g11691 ( 
.A1(n_10731),
.A2(n_7179),
.B(n_7191),
.Y(n_11691)
);

OAI22xp5_ASAP7_75t_L g11692 ( 
.A1(n_10554),
.A2(n_7750),
.B1(n_7757),
.B2(n_7732),
.Y(n_11692)
);

OAI22xp5_ASAP7_75t_L g11693 ( 
.A1(n_10994),
.A2(n_7750),
.B1(n_7757),
.B2(n_7732),
.Y(n_11693)
);

NAND2xp5_ASAP7_75t_SL g11694 ( 
.A(n_10735),
.B(n_8060),
.Y(n_11694)
);

NAND2xp5_ASAP7_75t_L g11695 ( 
.A(n_10589),
.B(n_8966),
.Y(n_11695)
);

NAND4xp25_ASAP7_75t_L g11696 ( 
.A(n_10567),
.B(n_7116),
.C(n_7500),
.D(n_7371),
.Y(n_11696)
);

NAND2xp5_ASAP7_75t_L g11697 ( 
.A(n_10589),
.B(n_8968),
.Y(n_11697)
);

AND2x2_ASAP7_75t_L g11698 ( 
.A(n_10775),
.B(n_9486),
.Y(n_11698)
);

AOI221xp5_ASAP7_75t_L g11699 ( 
.A1(n_10503),
.A2(n_7321),
.B1(n_7123),
.B2(n_7502),
.C(n_8968),
.Y(n_11699)
);

OAI22xp5_ASAP7_75t_L g11700 ( 
.A1(n_10995),
.A2(n_7757),
.B1(n_7777),
.B2(n_7750),
.Y(n_11700)
);

OAI21xp33_ASAP7_75t_L g11701 ( 
.A1(n_10935),
.A2(n_7363),
.B(n_7537),
.Y(n_11701)
);

NAND2xp5_ASAP7_75t_L g11702 ( 
.A(n_10631),
.B(n_8970),
.Y(n_11702)
);

AND2x2_ASAP7_75t_L g11703 ( 
.A(n_10780),
.B(n_10794),
.Y(n_11703)
);

HB1xp67_ASAP7_75t_L g11704 ( 
.A(n_10825),
.Y(n_11704)
);

AND2x2_ASAP7_75t_L g11705 ( 
.A(n_10542),
.B(n_9490),
.Y(n_11705)
);

AOI21xp5_ASAP7_75t_SL g11706 ( 
.A1(n_10736),
.A2(n_9912),
.B(n_9827),
.Y(n_11706)
);

NAND2xp5_ASAP7_75t_SL g11707 ( 
.A(n_10743),
.B(n_8060),
.Y(n_11707)
);

AOI22xp33_ASAP7_75t_SL g11708 ( 
.A1(n_10768),
.A2(n_6939),
.B1(n_6974),
.B2(n_6932),
.Y(n_11708)
);

NAND4xp25_ASAP7_75t_L g11709 ( 
.A(n_10600),
.B(n_10651),
.C(n_10700),
.D(n_10632),
.Y(n_11709)
);

AND2x2_ASAP7_75t_L g11710 ( 
.A(n_10542),
.B(n_9490),
.Y(n_11710)
);

NOR3xp33_ASAP7_75t_L g11711 ( 
.A(n_10486),
.B(n_7345),
.C(n_7341),
.Y(n_11711)
);

AOI22xp33_ASAP7_75t_SL g11712 ( 
.A1(n_10736),
.A2(n_6939),
.B1(n_6974),
.B2(n_6932),
.Y(n_11712)
);

AOI221xp5_ASAP7_75t_L g11713 ( 
.A1(n_10510),
.A2(n_7123),
.B1(n_8973),
.B2(n_8971),
.C(n_8970),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_10939),
.B(n_9500),
.Y(n_11714)
);

AND2x2_ASAP7_75t_L g11715 ( 
.A(n_10944),
.B(n_9500),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_10950),
.B(n_8681),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_10631),
.B(n_8971),
.Y(n_11717)
);

AND2x2_ASAP7_75t_L g11718 ( 
.A(n_11053),
.B(n_8702),
.Y(n_11718)
);

AND2x2_ASAP7_75t_L g11719 ( 
.A(n_11057),
.B(n_11076),
.Y(n_11719)
);

NAND3xp33_ASAP7_75t_L g11720 ( 
.A(n_11117),
.B(n_8119),
.C(n_8060),
.Y(n_11720)
);

AND2x4_ASAP7_75t_L g11721 ( 
.A(n_11553),
.B(n_10565),
.Y(n_11721)
);

INVx1_ASAP7_75t_SL g11722 ( 
.A(n_11179),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_11259),
.Y(n_11723)
);

OAI221xp5_ASAP7_75t_L g11724 ( 
.A1(n_11167),
.A2(n_10800),
.B1(n_10834),
.B2(n_10823),
.C(n_11085),
.Y(n_11724)
);

AND2x2_ASAP7_75t_L g11725 ( 
.A(n_11239),
.B(n_10631),
.Y(n_11725)
);

AOI22xp33_ASAP7_75t_L g11726 ( 
.A1(n_11206),
.A2(n_11000),
.B1(n_11001),
.B2(n_10997),
.Y(n_11726)
);

OR2x2_ASAP7_75t_L g11727 ( 
.A(n_11137),
.B(n_11198),
.Y(n_11727)
);

INVx1_ASAP7_75t_L g11728 ( 
.A(n_11326),
.Y(n_11728)
);

INVx2_ASAP7_75t_L g11729 ( 
.A(n_11661),
.Y(n_11729)
);

INVxp67_ASAP7_75t_SL g11730 ( 
.A(n_11195),
.Y(n_11730)
);

INVx1_ASAP7_75t_L g11731 ( 
.A(n_11413),
.Y(n_11731)
);

AND2x4_ASAP7_75t_L g11732 ( 
.A(n_11617),
.B(n_10800),
.Y(n_11732)
);

INVx4_ASAP7_75t_L g11733 ( 
.A(n_11150),
.Y(n_11733)
);

INVx2_ASAP7_75t_L g11734 ( 
.A(n_11661),
.Y(n_11734)
);

AND2x2_ASAP7_75t_L g11735 ( 
.A(n_11230),
.B(n_10635),
.Y(n_11735)
);

AND2x2_ASAP7_75t_L g11736 ( 
.A(n_11158),
.B(n_10635),
.Y(n_11736)
);

NAND2xp5_ASAP7_75t_L g11737 ( 
.A(n_11207),
.B(n_10635),
.Y(n_11737)
);

NAND3xp33_ASAP7_75t_L g11738 ( 
.A(n_11235),
.B(n_10694),
.C(n_10552),
.Y(n_11738)
);

INVx1_ASAP7_75t_L g11739 ( 
.A(n_11591),
.Y(n_11739)
);

OAI33xp33_ASAP7_75t_L g11740 ( 
.A1(n_11188),
.A2(n_10486),
.A3(n_10510),
.B1(n_10531),
.B2(n_10907),
.B3(n_10906),
.Y(n_11740)
);

BUFx3_ASAP7_75t_L g11741 ( 
.A(n_11273),
.Y(n_11741)
);

INVx2_ASAP7_75t_L g11742 ( 
.A(n_11314),
.Y(n_11742)
);

NAND2xp5_ASAP7_75t_L g11743 ( 
.A(n_11200),
.B(n_11165),
.Y(n_11743)
);

NOR2xp33_ASAP7_75t_L g11744 ( 
.A(n_11138),
.B(n_10694),
.Y(n_11744)
);

INVxp67_ASAP7_75t_L g11745 ( 
.A(n_11199),
.Y(n_11745)
);

INVx2_ASAP7_75t_L g11746 ( 
.A(n_11582),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_11704),
.Y(n_11747)
);

BUFx2_ASAP7_75t_L g11748 ( 
.A(n_11203),
.Y(n_11748)
);

NOR2xp33_ASAP7_75t_L g11749 ( 
.A(n_11367),
.B(n_10694),
.Y(n_11749)
);

INVx2_ASAP7_75t_L g11750 ( 
.A(n_11205),
.Y(n_11750)
);

AND2x2_ASAP7_75t_L g11751 ( 
.A(n_11153),
.B(n_11078),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_11578),
.Y(n_11752)
);

INVx2_ASAP7_75t_L g11753 ( 
.A(n_11252),
.Y(n_11753)
);

AOI33xp33_ASAP7_75t_L g11754 ( 
.A1(n_11213),
.A2(n_11096),
.A3(n_11105),
.B1(n_11095),
.B2(n_11019),
.B3(n_11002),
.Y(n_11754)
);

AOI21xp5_ASAP7_75t_L g11755 ( 
.A1(n_11170),
.A2(n_10737),
.B(n_10730),
.Y(n_11755)
);

INVx1_ASAP7_75t_L g11756 ( 
.A(n_11251),
.Y(n_11756)
);

INVx1_ASAP7_75t_L g11757 ( 
.A(n_11175),
.Y(n_11757)
);

INVx1_ASAP7_75t_L g11758 ( 
.A(n_11210),
.Y(n_11758)
);

INVx1_ASAP7_75t_L g11759 ( 
.A(n_11212),
.Y(n_11759)
);

AND2x2_ASAP7_75t_L g11760 ( 
.A(n_11247),
.B(n_11003),
.Y(n_11760)
);

INVx1_ASAP7_75t_L g11761 ( 
.A(n_11263),
.Y(n_11761)
);

AND2x4_ASAP7_75t_L g11762 ( 
.A(n_11305),
.B(n_10823),
.Y(n_11762)
);

OR2x2_ASAP7_75t_L g11763 ( 
.A(n_11627),
.B(n_10560),
.Y(n_11763)
);

INVxp67_ASAP7_75t_L g11764 ( 
.A(n_11193),
.Y(n_11764)
);

HB1xp67_ASAP7_75t_L g11765 ( 
.A(n_11187),
.Y(n_11765)
);

INVx1_ASAP7_75t_L g11766 ( 
.A(n_11429),
.Y(n_11766)
);

INVx1_ASAP7_75t_L g11767 ( 
.A(n_11269),
.Y(n_11767)
);

NAND2xp5_ASAP7_75t_L g11768 ( 
.A(n_11586),
.B(n_10746),
.Y(n_11768)
);

NAND2xp33_ASAP7_75t_L g11769 ( 
.A(n_11337),
.B(n_10740),
.Y(n_11769)
);

HB1xp67_ASAP7_75t_L g11770 ( 
.A(n_11187),
.Y(n_11770)
);

HB1xp67_ASAP7_75t_L g11771 ( 
.A(n_11460),
.Y(n_11771)
);

NAND3xp33_ASAP7_75t_L g11772 ( 
.A(n_11249),
.B(n_10907),
.C(n_10906),
.Y(n_11772)
);

HB1xp67_ASAP7_75t_L g11773 ( 
.A(n_11680),
.Y(n_11773)
);

INVx1_ASAP7_75t_L g11774 ( 
.A(n_11248),
.Y(n_11774)
);

INVx4_ASAP7_75t_L g11775 ( 
.A(n_11393),
.Y(n_11775)
);

AOI22xp33_ASAP7_75t_L g11776 ( 
.A1(n_11139),
.A2(n_10834),
.B1(n_10888),
.B2(n_10964),
.Y(n_11776)
);

AND2x4_ASAP7_75t_L g11777 ( 
.A(n_11478),
.B(n_10743),
.Y(n_11777)
);

INVx2_ASAP7_75t_L g11778 ( 
.A(n_11705),
.Y(n_11778)
);

AND2x2_ASAP7_75t_L g11779 ( 
.A(n_11220),
.B(n_10688),
.Y(n_11779)
);

HB1xp67_ASAP7_75t_L g11780 ( 
.A(n_11629),
.Y(n_11780)
);

NOR2x1_ASAP7_75t_SL g11781 ( 
.A(n_11268),
.B(n_7134),
.Y(n_11781)
);

HB1xp67_ASAP7_75t_L g11782 ( 
.A(n_11384),
.Y(n_11782)
);

INVx1_ASAP7_75t_L g11783 ( 
.A(n_11452),
.Y(n_11783)
);

INVx1_ASAP7_75t_L g11784 ( 
.A(n_11232),
.Y(n_11784)
);

BUFx2_ASAP7_75t_L g11785 ( 
.A(n_11308),
.Y(n_11785)
);

AND2x2_ASAP7_75t_L g11786 ( 
.A(n_11204),
.B(n_10688),
.Y(n_11786)
);

INVx1_ASAP7_75t_L g11787 ( 
.A(n_11234),
.Y(n_11787)
);

INVx2_ASAP7_75t_L g11788 ( 
.A(n_11710),
.Y(n_11788)
);

OR2x2_ASAP7_75t_L g11789 ( 
.A(n_11145),
.B(n_11049),
.Y(n_11789)
);

AND2x2_ASAP7_75t_L g11790 ( 
.A(n_11246),
.B(n_10708),
.Y(n_11790)
);

INVx1_ASAP7_75t_L g11791 ( 
.A(n_11456),
.Y(n_11791)
);

INVxp67_ASAP7_75t_L g11792 ( 
.A(n_11638),
.Y(n_11792)
);

AND2x2_ASAP7_75t_L g11793 ( 
.A(n_11237),
.B(n_10708),
.Y(n_11793)
);

INVxp67_ASAP7_75t_SL g11794 ( 
.A(n_11217),
.Y(n_11794)
);

AND2x2_ASAP7_75t_L g11795 ( 
.A(n_11343),
.B(n_11154),
.Y(n_11795)
);

INVx2_ASAP7_75t_L g11796 ( 
.A(n_11157),
.Y(n_11796)
);

HB1xp67_ASAP7_75t_L g11797 ( 
.A(n_11147),
.Y(n_11797)
);

NAND4xp25_ASAP7_75t_L g11798 ( 
.A(n_11227),
.B(n_10632),
.C(n_10651),
.D(n_10600),
.Y(n_11798)
);

AND2x2_ASAP7_75t_L g11799 ( 
.A(n_11133),
.B(n_10634),
.Y(n_11799)
);

INVx1_ASAP7_75t_L g11800 ( 
.A(n_11457),
.Y(n_11800)
);

AO21x2_ASAP7_75t_L g11801 ( 
.A1(n_11217),
.A2(n_10460),
.B(n_10955),
.Y(n_11801)
);

INVx2_ASAP7_75t_L g11802 ( 
.A(n_11243),
.Y(n_11802)
);

OR2x2_ASAP7_75t_L g11803 ( 
.A(n_11185),
.B(n_11049),
.Y(n_11803)
);

NAND4xp25_ASAP7_75t_L g11804 ( 
.A(n_11227),
.B(n_10726),
.C(n_10727),
.D(n_10700),
.Y(n_11804)
);

INVx1_ASAP7_75t_L g11805 ( 
.A(n_11571),
.Y(n_11805)
);

AND2x2_ASAP7_75t_L g11806 ( 
.A(n_11136),
.B(n_10634),
.Y(n_11806)
);

AND2x2_ASAP7_75t_L g11807 ( 
.A(n_11134),
.B(n_10640),
.Y(n_11807)
);

NAND2xp5_ASAP7_75t_L g11808 ( 
.A(n_11163),
.B(n_10748),
.Y(n_11808)
);

OAI22xp5_ASAP7_75t_L g11809 ( 
.A1(n_11168),
.A2(n_10732),
.B1(n_10785),
.B2(n_10792),
.Y(n_11809)
);

OAI21xp5_ASAP7_75t_SL g11810 ( 
.A1(n_11143),
.A2(n_10727),
.B(n_10726),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_11584),
.Y(n_11811)
);

OAI221xp5_ASAP7_75t_L g11812 ( 
.A1(n_11216),
.A2(n_11082),
.B1(n_11038),
.B2(n_10784),
.C(n_10830),
.Y(n_11812)
);

HB1xp67_ASAP7_75t_L g11813 ( 
.A(n_11485),
.Y(n_11813)
);

AND2x2_ASAP7_75t_L g11814 ( 
.A(n_11141),
.B(n_10640),
.Y(n_11814)
);

AND2x2_ASAP7_75t_L g11815 ( 
.A(n_11644),
.B(n_10842),
.Y(n_11815)
);

INVx1_ASAP7_75t_L g11816 ( 
.A(n_11589),
.Y(n_11816)
);

AND2x4_ASAP7_75t_L g11817 ( 
.A(n_11490),
.B(n_10578),
.Y(n_11817)
);

AND2x2_ASAP7_75t_L g11818 ( 
.A(n_11228),
.B(n_10842),
.Y(n_11818)
);

AND2x2_ASAP7_75t_L g11819 ( 
.A(n_11556),
.B(n_10865),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11250),
.B(n_10865),
.Y(n_11820)
);

OAI22xp5_ASAP7_75t_L g11821 ( 
.A1(n_11183),
.A2(n_10742),
.B1(n_11122),
.B2(n_11120),
.Y(n_11821)
);

OR2x2_ASAP7_75t_L g11822 ( 
.A(n_11240),
.B(n_11082),
.Y(n_11822)
);

HB1xp67_ASAP7_75t_L g11823 ( 
.A(n_11149),
.Y(n_11823)
);

INVx2_ASAP7_75t_L g11824 ( 
.A(n_11587),
.Y(n_11824)
);

NAND3xp33_ASAP7_75t_L g11825 ( 
.A(n_11152),
.B(n_10914),
.C(n_11124),
.Y(n_11825)
);

OAI321xp33_ASAP7_75t_L g11826 ( 
.A1(n_11181),
.A2(n_10965),
.A3(n_10784),
.B1(n_10815),
.B2(n_10830),
.C(n_10763),
.Y(n_11826)
);

NAND2x1p5_ASAP7_75t_L g11827 ( 
.A(n_11298),
.B(n_10578),
.Y(n_11827)
);

AND2x2_ASAP7_75t_L g11828 ( 
.A(n_11703),
.B(n_10877),
.Y(n_11828)
);

INVx2_ASAP7_75t_L g11829 ( 
.A(n_11587),
.Y(n_11829)
);

INVx1_ASAP7_75t_L g11830 ( 
.A(n_11590),
.Y(n_11830)
);

INVx2_ASAP7_75t_L g11831 ( 
.A(n_11604),
.Y(n_11831)
);

AND2x2_ASAP7_75t_L g11832 ( 
.A(n_11426),
.B(n_10877),
.Y(n_11832)
);

AOI31xp33_ASAP7_75t_L g11833 ( 
.A1(n_11146),
.A2(n_10527),
.A3(n_10914),
.B(n_10815),
.Y(n_11833)
);

INVx2_ASAP7_75t_L g11834 ( 
.A(n_11604),
.Y(n_11834)
);

INVx1_ASAP7_75t_L g11835 ( 
.A(n_11596),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_11598),
.Y(n_11836)
);

INVx4_ASAP7_75t_L g11837 ( 
.A(n_11400),
.Y(n_11837)
);

HB1xp67_ASAP7_75t_L g11838 ( 
.A(n_11349),
.Y(n_11838)
);

INVx2_ASAP7_75t_L g11839 ( 
.A(n_11664),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_11261),
.Y(n_11840)
);

HB1xp67_ASAP7_75t_L g11841 ( 
.A(n_11189),
.Y(n_11841)
);

INVx3_ASAP7_75t_L g11842 ( 
.A(n_11558),
.Y(n_11842)
);

BUFx2_ASAP7_75t_L g11843 ( 
.A(n_11528),
.Y(n_11843)
);

INVx4_ASAP7_75t_L g11844 ( 
.A(n_11581),
.Y(n_11844)
);

AOI211xp5_ASAP7_75t_L g11845 ( 
.A1(n_11140),
.A2(n_10763),
.B(n_10952),
.C(n_10929),
.Y(n_11845)
);

INVx1_ASAP7_75t_L g11846 ( 
.A(n_11262),
.Y(n_11846)
);

INVx2_ASAP7_75t_L g11847 ( 
.A(n_11664),
.Y(n_11847)
);

INVx1_ASAP7_75t_L g11848 ( 
.A(n_11634),
.Y(n_11848)
);

BUFx2_ASAP7_75t_L g11849 ( 
.A(n_11508),
.Y(n_11849)
);

AO221x2_ASAP7_75t_L g11850 ( 
.A1(n_11152),
.A2(n_10757),
.B1(n_10753),
.B2(n_10990),
.C(n_10812),
.Y(n_11850)
);

OR2x2_ASAP7_75t_L g11851 ( 
.A(n_11241),
.B(n_11038),
.Y(n_11851)
);

INVx1_ASAP7_75t_L g11852 ( 
.A(n_11180),
.Y(n_11852)
);

OAI221xp5_ASAP7_75t_L g11853 ( 
.A1(n_11148),
.A2(n_10855),
.B1(n_10870),
.B2(n_10893),
.C(n_10895),
.Y(n_11853)
);

INVx2_ASAP7_75t_L g11854 ( 
.A(n_11554),
.Y(n_11854)
);

INVx1_ASAP7_75t_L g11855 ( 
.A(n_11448),
.Y(n_11855)
);

INVx1_ASAP7_75t_L g11856 ( 
.A(n_11450),
.Y(n_11856)
);

INVx2_ASAP7_75t_L g11857 ( 
.A(n_11689),
.Y(n_11857)
);

NAND4xp25_ASAP7_75t_SL g11858 ( 
.A(n_11151),
.B(n_10870),
.C(n_10855),
.D(n_10821),
.Y(n_11858)
);

OR2x2_ASAP7_75t_L g11859 ( 
.A(n_11453),
.B(n_10898),
.Y(n_11859)
);

AND2x2_ASAP7_75t_L g11860 ( 
.A(n_11271),
.B(n_10912),
.Y(n_11860)
);

INVx2_ASAP7_75t_L g11861 ( 
.A(n_11585),
.Y(n_11861)
);

INVx1_ASAP7_75t_L g11862 ( 
.A(n_11454),
.Y(n_11862)
);

AND2x2_ASAP7_75t_L g11863 ( 
.A(n_11493),
.B(n_10912),
.Y(n_11863)
);

NOR2x1_ASAP7_75t_SL g11864 ( 
.A(n_11357),
.B(n_7134),
.Y(n_11864)
);

INVx3_ASAP7_75t_L g11865 ( 
.A(n_11573),
.Y(n_11865)
);

INVx2_ASAP7_75t_SL g11866 ( 
.A(n_11385),
.Y(n_11866)
);

INVx2_ASAP7_75t_L g11867 ( 
.A(n_11671),
.Y(n_11867)
);

AND2x2_ASAP7_75t_L g11868 ( 
.A(n_11299),
.B(n_10582),
.Y(n_11868)
);

OAI211xp5_ASAP7_75t_L g11869 ( 
.A1(n_11201),
.A2(n_10929),
.B(n_10952),
.C(n_10811),
.Y(n_11869)
);

OAI211xp5_ASAP7_75t_SL g11870 ( 
.A1(n_11178),
.A2(n_10965),
.B(n_10925),
.C(n_10885),
.Y(n_11870)
);

AND2x2_ASAP7_75t_L g11871 ( 
.A(n_11302),
.B(n_10582),
.Y(n_11871)
);

INVx1_ASAP7_75t_SL g11872 ( 
.A(n_11417),
.Y(n_11872)
);

NAND2xp5_ASAP7_75t_L g11873 ( 
.A(n_11291),
.B(n_10826),
.Y(n_11873)
);

INVx1_ASAP7_75t_L g11874 ( 
.A(n_11455),
.Y(n_11874)
);

NOR2xp33_ASAP7_75t_SL g11875 ( 
.A(n_11169),
.B(n_7062),
.Y(n_11875)
);

INVx2_ASAP7_75t_L g11876 ( 
.A(n_11681),
.Y(n_11876)
);

AND2x2_ASAP7_75t_L g11877 ( 
.A(n_11495),
.B(n_10967),
.Y(n_11877)
);

NAND2xp5_ASAP7_75t_L g11878 ( 
.A(n_11574),
.B(n_10832),
.Y(n_11878)
);

BUFx6f_ASAP7_75t_L g11879 ( 
.A(n_11375),
.Y(n_11879)
);

NAND2xp5_ASAP7_75t_L g11880 ( 
.A(n_11340),
.B(n_10833),
.Y(n_11880)
);

AO21x2_ASAP7_75t_L g11881 ( 
.A1(n_11364),
.A2(n_10959),
.B(n_10955),
.Y(n_11881)
);

OAI33xp33_ASAP7_75t_L g11882 ( 
.A1(n_11348),
.A2(n_10838),
.A3(n_10836),
.B1(n_10518),
.B2(n_10492),
.B3(n_10519),
.Y(n_11882)
);

AND2x2_ASAP7_75t_L g11883 ( 
.A(n_11575),
.B(n_10971),
.Y(n_11883)
);

OR2x2_ASAP7_75t_L g11884 ( 
.A(n_11238),
.B(n_10934),
.Y(n_11884)
);

AOI322xp5_ASAP7_75t_L g11885 ( 
.A1(n_11675),
.A2(n_10970),
.A3(n_10966),
.B1(n_10977),
.B2(n_10968),
.C1(n_10959),
.C2(n_10540),
.Y(n_11885)
);

INVx1_ASAP7_75t_SL g11886 ( 
.A(n_11447),
.Y(n_11886)
);

AO31x2_ASAP7_75t_L g11887 ( 
.A1(n_11144),
.A2(n_10516),
.A3(n_10521),
.B(n_10490),
.Y(n_11887)
);

OAI221xp5_ASAP7_75t_L g11888 ( 
.A1(n_11172),
.A2(n_11258),
.B1(n_11177),
.B2(n_11244),
.C(n_11236),
.Y(n_11888)
);

HB1xp67_ASAP7_75t_L g11889 ( 
.A(n_11469),
.Y(n_11889)
);

INVx2_ASAP7_75t_L g11890 ( 
.A(n_11687),
.Y(n_11890)
);

INVx1_ASAP7_75t_L g11891 ( 
.A(n_11491),
.Y(n_11891)
);

INVx1_ASAP7_75t_L g11892 ( 
.A(n_11491),
.Y(n_11892)
);

AND2x2_ASAP7_75t_L g11893 ( 
.A(n_11510),
.B(n_10972),
.Y(n_11893)
);

AND2x2_ASAP7_75t_L g11894 ( 
.A(n_11275),
.B(n_10975),
.Y(n_11894)
);

INVx3_ASAP7_75t_L g11895 ( 
.A(n_11716),
.Y(n_11895)
);

AOI22xp33_ASAP7_75t_L g11896 ( 
.A1(n_11162),
.A2(n_10986),
.B1(n_10988),
.B2(n_10983),
.Y(n_11896)
);

NAND2xp5_ASAP7_75t_SL g11897 ( 
.A(n_11182),
.B(n_10770),
.Y(n_11897)
);

NAND2xp5_ASAP7_75t_L g11898 ( 
.A(n_11534),
.B(n_10989),
.Y(n_11898)
);

AND2x2_ASAP7_75t_L g11899 ( 
.A(n_11215),
.B(n_11288),
.Y(n_11899)
);

INVx2_ASAP7_75t_L g11900 ( 
.A(n_11559),
.Y(n_11900)
);

INVx2_ASAP7_75t_L g11901 ( 
.A(n_11579),
.Y(n_11901)
);

AND2x2_ASAP7_75t_L g11902 ( 
.A(n_11359),
.B(n_10996),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_11467),
.Y(n_11903)
);

INVx2_ASAP7_75t_L g11904 ( 
.A(n_11583),
.Y(n_11904)
);

INVx1_ASAP7_75t_L g11905 ( 
.A(n_11470),
.Y(n_11905)
);

HB1xp67_ASAP7_75t_L g11906 ( 
.A(n_11469),
.Y(n_11906)
);

INVx1_ASAP7_75t_L g11907 ( 
.A(n_11474),
.Y(n_11907)
);

OAI33xp33_ASAP7_75t_L g11908 ( 
.A1(n_11142),
.A2(n_10547),
.A3(n_10541),
.B1(n_10549),
.B2(n_10543),
.B3(n_10535),
.Y(n_11908)
);

NAND2xp5_ASAP7_75t_L g11909 ( 
.A(n_11438),
.B(n_11004),
.Y(n_11909)
);

INVx1_ASAP7_75t_L g11910 ( 
.A(n_11476),
.Y(n_11910)
);

AND2x2_ASAP7_75t_L g11911 ( 
.A(n_11399),
.B(n_11006),
.Y(n_11911)
);

OAI22xp5_ASAP7_75t_L g11912 ( 
.A1(n_11622),
.A2(n_11074),
.B1(n_11061),
.B2(n_11047),
.Y(n_11912)
);

OR2x2_ASAP7_75t_L g11913 ( 
.A(n_11312),
.B(n_10943),
.Y(n_11913)
);

INVx2_ASAP7_75t_L g11914 ( 
.A(n_11595),
.Y(n_11914)
);

OR2x2_ASAP7_75t_L g11915 ( 
.A(n_11316),
.B(n_11306),
.Y(n_11915)
);

OR2x2_ASAP7_75t_L g11916 ( 
.A(n_11537),
.B(n_11226),
.Y(n_11916)
);

INVx1_ASAP7_75t_SL g11917 ( 
.A(n_11382),
.Y(n_11917)
);

HB1xp67_ASAP7_75t_L g11918 ( 
.A(n_11486),
.Y(n_11918)
);

NOR2xp67_ASAP7_75t_L g11919 ( 
.A(n_11486),
.B(n_11489),
.Y(n_11919)
);

AND2x2_ASAP7_75t_L g11920 ( 
.A(n_11446),
.B(n_11015),
.Y(n_11920)
);

HB1xp67_ASAP7_75t_L g11921 ( 
.A(n_11489),
.Y(n_11921)
);

OR2x2_ASAP7_75t_L g11922 ( 
.A(n_11296),
.B(n_11022),
.Y(n_11922)
);

NOR3xp33_ASAP7_75t_L g11923 ( 
.A(n_11171),
.B(n_10563),
.C(n_10550),
.Y(n_11923)
);

HB1xp67_ASAP7_75t_L g11924 ( 
.A(n_11229),
.Y(n_11924)
);

AO21x2_ASAP7_75t_L g11925 ( 
.A1(n_11211),
.A2(n_10577),
.B(n_10572),
.Y(n_11925)
);

INVxp67_ASAP7_75t_SL g11926 ( 
.A(n_11211),
.Y(n_11926)
);

NAND3xp33_ASAP7_75t_L g11927 ( 
.A(n_11142),
.B(n_10610),
.C(n_10592),
.Y(n_11927)
);

INVx2_ASAP7_75t_L g11928 ( 
.A(n_11714),
.Y(n_11928)
);

AND2x2_ASAP7_75t_L g11929 ( 
.A(n_11567),
.B(n_11016),
.Y(n_11929)
);

BUFx3_ASAP7_75t_L g11930 ( 
.A(n_11160),
.Y(n_11930)
);

AOI22xp33_ASAP7_75t_SL g11931 ( 
.A1(n_11231),
.A2(n_11190),
.B1(n_11184),
.B2(n_11223),
.Y(n_11931)
);

INVx2_ASAP7_75t_SL g11932 ( 
.A(n_11494),
.Y(n_11932)
);

INVx2_ASAP7_75t_SL g11933 ( 
.A(n_11670),
.Y(n_11933)
);

AND2x2_ASAP7_75t_L g11934 ( 
.A(n_11719),
.B(n_11612),
.Y(n_11934)
);

AND2x2_ASAP7_75t_L g11935 ( 
.A(n_11621),
.B(n_11020),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_11505),
.Y(n_11936)
);

INVx2_ASAP7_75t_L g11937 ( 
.A(n_11715),
.Y(n_11937)
);

OR2x2_ASAP7_75t_L g11938 ( 
.A(n_11303),
.B(n_11125),
.Y(n_11938)
);

INVxp67_ASAP7_75t_SL g11939 ( 
.A(n_11285),
.Y(n_11939)
);

AND2x2_ASAP7_75t_L g11940 ( 
.A(n_11623),
.B(n_11024),
.Y(n_11940)
);

AND2x2_ASAP7_75t_L g11941 ( 
.A(n_11624),
.B(n_10981),
.Y(n_11941)
);

AOI22xp33_ASAP7_75t_L g11942 ( 
.A1(n_11242),
.A2(n_11045),
.B1(n_11043),
.B2(n_11048),
.Y(n_11942)
);

AND2x2_ASAP7_75t_L g11943 ( 
.A(n_11635),
.B(n_10706),
.Y(n_11943)
);

AOI22xp33_ASAP7_75t_L g11944 ( 
.A1(n_11557),
.A2(n_11127),
.B1(n_8207),
.B2(n_8241),
.Y(n_11944)
);

INVxp67_ASAP7_75t_L g11945 ( 
.A(n_11539),
.Y(n_11945)
);

NAND3xp33_ASAP7_75t_SL g11946 ( 
.A(n_11507),
.B(n_8658),
.C(n_8646),
.Y(n_11946)
);

AOI222xp33_ASAP7_75t_L g11947 ( 
.A1(n_11156),
.A2(n_10618),
.B1(n_10611),
.B2(n_10624),
.C1(n_10620),
.C2(n_10614),
.Y(n_11947)
);

INVx1_ASAP7_75t_L g11948 ( 
.A(n_11505),
.Y(n_11948)
);

INVxp67_ASAP7_75t_SL g11949 ( 
.A(n_11286),
.Y(n_11949)
);

INVx2_ASAP7_75t_L g11950 ( 
.A(n_11394),
.Y(n_11950)
);

AND2x2_ASAP7_75t_L g11951 ( 
.A(n_11641),
.B(n_10706),
.Y(n_11951)
);

INVx1_ASAP7_75t_L g11952 ( 
.A(n_11509),
.Y(n_11952)
);

INVx2_ASAP7_75t_L g11953 ( 
.A(n_11549),
.Y(n_11953)
);

INVx2_ASAP7_75t_L g11954 ( 
.A(n_11499),
.Y(n_11954)
);

OAI21xp5_ASAP7_75t_L g11955 ( 
.A1(n_11223),
.A2(n_11127),
.B(n_10630),
.Y(n_11955)
);

INVx3_ASAP7_75t_L g11956 ( 
.A(n_11550),
.Y(n_11956)
);

INVx2_ASAP7_75t_L g11957 ( 
.A(n_11414),
.Y(n_11957)
);

INVx3_ASAP7_75t_SL g11958 ( 
.A(n_11272),
.Y(n_11958)
);

NOR2xp33_ASAP7_75t_L g11959 ( 
.A(n_11561),
.B(n_11135),
.Y(n_11959)
);

CKINVDCx20_ASAP7_75t_R g11960 ( 
.A(n_11356),
.Y(n_11960)
);

BUFx2_ASAP7_75t_SL g11961 ( 
.A(n_11295),
.Y(n_11961)
);

AOI33xp33_ASAP7_75t_L g11962 ( 
.A1(n_11390),
.A2(n_10659),
.A3(n_10643),
.B1(n_10662),
.B2(n_10653),
.B3(n_10629),
.Y(n_11962)
);

INVx2_ASAP7_75t_L g11963 ( 
.A(n_11424),
.Y(n_11963)
);

OAI33xp33_ASAP7_75t_L g11964 ( 
.A1(n_11156),
.A2(n_10676),
.A3(n_10667),
.B1(n_10677),
.B2(n_10670),
.B3(n_10663),
.Y(n_11964)
);

AND2x2_ASAP7_75t_L g11965 ( 
.A(n_11643),
.B(n_10706),
.Y(n_11965)
);

HB1xp67_ASAP7_75t_L g11966 ( 
.A(n_11214),
.Y(n_11966)
);

OAI22xp5_ASAP7_75t_L g11967 ( 
.A1(n_11254),
.A2(n_7777),
.B1(n_7784),
.B2(n_7783),
.Y(n_11967)
);

OR2x2_ASAP7_75t_L g11968 ( 
.A(n_11442),
.B(n_11034),
.Y(n_11968)
);

AND2x2_ASAP7_75t_L g11969 ( 
.A(n_11645),
.B(n_11034),
.Y(n_11969)
);

INVx3_ASAP7_75t_L g11970 ( 
.A(n_11550),
.Y(n_11970)
);

INVx1_ASAP7_75t_L g11971 ( 
.A(n_11270),
.Y(n_11971)
);

HB1xp67_ASAP7_75t_L g11972 ( 
.A(n_11577),
.Y(n_11972)
);

INVx4_ASAP7_75t_L g11973 ( 
.A(n_11451),
.Y(n_11973)
);

INVx1_ASAP7_75t_SL g11974 ( 
.A(n_11718),
.Y(n_11974)
);

AO21x2_ASAP7_75t_L g11975 ( 
.A1(n_11159),
.A2(n_10682),
.B(n_10681),
.Y(n_11975)
);

NAND2xp5_ASAP7_75t_L g11976 ( 
.A(n_11161),
.B(n_10686),
.Y(n_11976)
);

AND2x2_ASAP7_75t_L g11977 ( 
.A(n_11650),
.B(n_11034),
.Y(n_11977)
);

INVx1_ASAP7_75t_L g11978 ( 
.A(n_11274),
.Y(n_11978)
);

NAND2xp5_ASAP7_75t_L g11979 ( 
.A(n_11155),
.B(n_10692),
.Y(n_11979)
);

NAND4xp25_ASAP7_75t_L g11980 ( 
.A(n_11197),
.B(n_10693),
.C(n_10701),
.D(n_10696),
.Y(n_11980)
);

NAND4xp25_ASAP7_75t_SL g11981 ( 
.A(n_11370),
.B(n_10702),
.C(n_10713),
.D(n_10711),
.Y(n_11981)
);

AO21x2_ASAP7_75t_L g11982 ( 
.A1(n_11159),
.A2(n_10723),
.B(n_10717),
.Y(n_11982)
);

AND2x2_ASAP7_75t_L g11983 ( 
.A(n_11651),
.B(n_10728),
.Y(n_11983)
);

INVx1_ASAP7_75t_SL g11984 ( 
.A(n_11482),
.Y(n_11984)
);

BUFx2_ASAP7_75t_L g11985 ( 
.A(n_11685),
.Y(n_11985)
);

BUFx3_ASAP7_75t_L g11986 ( 
.A(n_11283),
.Y(n_11986)
);

OAI221xp5_ASAP7_75t_L g11987 ( 
.A1(n_11245),
.A2(n_10755),
.B1(n_10758),
.B2(n_10741),
.C(n_10738),
.Y(n_11987)
);

NAND2xp5_ASAP7_75t_L g11988 ( 
.A(n_11339),
.B(n_10769),
.Y(n_11988)
);

INVx1_ASAP7_75t_L g11989 ( 
.A(n_11309),
.Y(n_11989)
);

HB1xp67_ASAP7_75t_L g11990 ( 
.A(n_11397),
.Y(n_11990)
);

BUFx2_ASAP7_75t_L g11991 ( 
.A(n_11329),
.Y(n_11991)
);

AND2x2_ASAP7_75t_L g11992 ( 
.A(n_11667),
.B(n_10774),
.Y(n_11992)
);

INVx5_ASAP7_75t_SL g11993 ( 
.A(n_11560),
.Y(n_11993)
);

NAND2xp5_ASAP7_75t_L g11994 ( 
.A(n_11328),
.B(n_11514),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11603),
.B(n_10778),
.Y(n_11995)
);

INVx1_ASAP7_75t_SL g11996 ( 
.A(n_11196),
.Y(n_11996)
);

INVx1_ASAP7_75t_L g11997 ( 
.A(n_11310),
.Y(n_11997)
);

AND2x2_ASAP7_75t_L g11998 ( 
.A(n_11606),
.B(n_10779),
.Y(n_11998)
);

INVx1_ASAP7_75t_L g11999 ( 
.A(n_11545),
.Y(n_11999)
);

AND2x2_ASAP7_75t_L g12000 ( 
.A(n_11611),
.B(n_11351),
.Y(n_12000)
);

HB1xp67_ASAP7_75t_L g12001 ( 
.A(n_11406),
.Y(n_12001)
);

AND2x2_ASAP7_75t_L g12002 ( 
.A(n_11307),
.B(n_10795),
.Y(n_12002)
);

INVx1_ASAP7_75t_L g12003 ( 
.A(n_11545),
.Y(n_12003)
);

OAI221xp5_ASAP7_75t_L g12004 ( 
.A1(n_11320),
.A2(n_10817),
.B1(n_10819),
.B2(n_10810),
.C(n_10804),
.Y(n_12004)
);

OR2x2_ASAP7_75t_L g12005 ( 
.A(n_11257),
.B(n_10687),
.Y(n_12005)
);

AND2x2_ASAP7_75t_L g12006 ( 
.A(n_11319),
.B(n_10822),
.Y(n_12006)
);

NAND2xp5_ASAP7_75t_L g12007 ( 
.A(n_11208),
.B(n_10824),
.Y(n_12007)
);

OAI221xp5_ASAP7_75t_L g12008 ( 
.A1(n_11202),
.A2(n_8119),
.B1(n_8410),
.B2(n_8280),
.C(n_8060),
.Y(n_12008)
);

INVx1_ASAP7_75t_L g12009 ( 
.A(n_11551),
.Y(n_12009)
);

BUFx2_ASAP7_75t_L g12010 ( 
.A(n_11472),
.Y(n_12010)
);

NAND2xp5_ASAP7_75t_L g12011 ( 
.A(n_11324),
.B(n_10687),
.Y(n_12011)
);

INVxp67_ASAP7_75t_SL g12012 ( 
.A(n_11536),
.Y(n_12012)
);

AND2x2_ASAP7_75t_L g12013 ( 
.A(n_11425),
.B(n_10687),
.Y(n_12013)
);

AOI32xp33_ASAP7_75t_L g12014 ( 
.A1(n_11699),
.A2(n_8203),
.A3(n_8222),
.B1(n_8219),
.B2(n_8177),
.Y(n_12014)
);

INVx2_ASAP7_75t_L g12015 ( 
.A(n_11698),
.Y(n_12015)
);

OR2x2_ASAP7_75t_L g12016 ( 
.A(n_11260),
.B(n_10733),
.Y(n_12016)
);

OR2x2_ASAP7_75t_L g12017 ( 
.A(n_11281),
.B(n_10733),
.Y(n_12017)
);

AND2x2_ASAP7_75t_L g12018 ( 
.A(n_11347),
.B(n_11365),
.Y(n_12018)
);

AND2x2_ASAP7_75t_L g12019 ( 
.A(n_11412),
.B(n_10733),
.Y(n_12019)
);

AO21x2_ASAP7_75t_L g12020 ( 
.A1(n_11536),
.A2(n_8974),
.B(n_8973),
.Y(n_12020)
);

AND2x2_ASAP7_75t_L g12021 ( 
.A(n_11279),
.B(n_7834),
.Y(n_12021)
);

OAI31xp33_ASAP7_75t_L g12022 ( 
.A1(n_11265),
.A2(n_7429),
.A3(n_7337),
.B(n_7388),
.Y(n_12022)
);

INVxp67_ASAP7_75t_SL g12023 ( 
.A(n_11551),
.Y(n_12023)
);

INVx1_ASAP7_75t_L g12024 ( 
.A(n_11662),
.Y(n_12024)
);

BUFx3_ASAP7_75t_L g12025 ( 
.A(n_11221),
.Y(n_12025)
);

AND2x2_ASAP7_75t_L g12026 ( 
.A(n_11282),
.B(n_7834),
.Y(n_12026)
);

OR2x6_ASAP7_75t_L g12027 ( 
.A(n_11568),
.B(n_6932),
.Y(n_12027)
);

INVx1_ASAP7_75t_L g12028 ( 
.A(n_11669),
.Y(n_12028)
);

NOR2xp33_ASAP7_75t_L g12029 ( 
.A(n_11642),
.B(n_8659),
.Y(n_12029)
);

INVx1_ASAP7_75t_SL g12030 ( 
.A(n_11224),
.Y(n_12030)
);

INVx2_ASAP7_75t_L g12031 ( 
.A(n_11503),
.Y(n_12031)
);

AND2x2_ASAP7_75t_L g12032 ( 
.A(n_11287),
.B(n_7834),
.Y(n_12032)
);

HB1xp67_ASAP7_75t_L g12033 ( 
.A(n_11630),
.Y(n_12033)
);

NOR2x1_ASAP7_75t_SL g12034 ( 
.A(n_11509),
.B(n_8060),
.Y(n_12034)
);

AND2x2_ASAP7_75t_L g12035 ( 
.A(n_11276),
.B(n_11363),
.Y(n_12035)
);

NAND2xp5_ASAP7_75t_L g12036 ( 
.A(n_11192),
.B(n_8974),
.Y(n_12036)
);

INVx4_ASAP7_75t_L g12037 ( 
.A(n_11466),
.Y(n_12037)
);

OAI33xp33_ASAP7_75t_L g12038 ( 
.A1(n_11458),
.A2(n_8980),
.A3(n_8977),
.B1(n_8984),
.B2(n_8979),
.B3(n_8976),
.Y(n_12038)
);

INVx1_ASAP7_75t_L g12039 ( 
.A(n_11672),
.Y(n_12039)
);

AND2x4_ASAP7_75t_L g12040 ( 
.A(n_11284),
.B(n_8060),
.Y(n_12040)
);

HB1xp67_ASAP7_75t_L g12041 ( 
.A(n_11631),
.Y(n_12041)
);

INVx2_ASAP7_75t_L g12042 ( 
.A(n_11506),
.Y(n_12042)
);

INVx1_ASAP7_75t_SL g12043 ( 
.A(n_11462),
.Y(n_12043)
);

INVx1_ASAP7_75t_L g12044 ( 
.A(n_11674),
.Y(n_12044)
);

AND2x4_ASAP7_75t_SL g12045 ( 
.A(n_11389),
.B(n_7074),
.Y(n_12045)
);

INVx1_ASAP7_75t_L g12046 ( 
.A(n_11321),
.Y(n_12046)
);

OR2x2_ASAP7_75t_L g12047 ( 
.A(n_11318),
.B(n_8976),
.Y(n_12047)
);

AND2x2_ASAP7_75t_L g12048 ( 
.A(n_11368),
.B(n_11376),
.Y(n_12048)
);

NOR2x1_ASAP7_75t_L g12049 ( 
.A(n_11218),
.B(n_6850),
.Y(n_12049)
);

HB1xp67_ASAP7_75t_L g12050 ( 
.A(n_11633),
.Y(n_12050)
);

INVx2_ASAP7_75t_L g12051 ( 
.A(n_11513),
.Y(n_12051)
);

AND2x2_ASAP7_75t_L g12052 ( 
.A(n_11379),
.B(n_11380),
.Y(n_12052)
);

AND2x2_ASAP7_75t_L g12053 ( 
.A(n_11712),
.B(n_9915),
.Y(n_12053)
);

INVx1_ASAP7_75t_L g12054 ( 
.A(n_11325),
.Y(n_12054)
);

INVx2_ASAP7_75t_SL g12055 ( 
.A(n_11677),
.Y(n_12055)
);

NAND2xp5_ASAP7_75t_L g12056 ( 
.A(n_11194),
.B(n_8977),
.Y(n_12056)
);

AO31x2_ASAP7_75t_L g12057 ( 
.A1(n_11166),
.A2(n_9081),
.A3(n_9088),
.B(n_9079),
.Y(n_12057)
);

BUFx2_ASAP7_75t_L g12058 ( 
.A(n_11636),
.Y(n_12058)
);

AOI21xp5_ASAP7_75t_L g12059 ( 
.A1(n_11267),
.A2(n_11218),
.B(n_11317),
.Y(n_12059)
);

INVx4_ASAP7_75t_L g12060 ( 
.A(n_11501),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11566),
.Y(n_12061)
);

NAND2xp5_ASAP7_75t_SL g12062 ( 
.A(n_11407),
.B(n_8060),
.Y(n_12062)
);

AOI22xp5_ASAP7_75t_L g12063 ( 
.A1(n_11576),
.A2(n_7783),
.B1(n_7784),
.B2(n_7777),
.Y(n_12063)
);

INVx2_ASAP7_75t_L g12064 ( 
.A(n_11524),
.Y(n_12064)
);

OAI33xp33_ASAP7_75t_L g12065 ( 
.A1(n_11458),
.A2(n_8989),
.A3(n_8980),
.B1(n_8994),
.B2(n_8984),
.B3(n_8979),
.Y(n_12065)
);

AND2x2_ASAP7_75t_L g12066 ( 
.A(n_11278),
.B(n_9941),
.Y(n_12066)
);

HB1xp67_ASAP7_75t_L g12067 ( 
.A(n_11637),
.Y(n_12067)
);

OR2x2_ASAP7_75t_L g12068 ( 
.A(n_11277),
.B(n_11709),
.Y(n_12068)
);

INVx1_ASAP7_75t_SL g12069 ( 
.A(n_11463),
.Y(n_12069)
);

AND2x2_ASAP7_75t_L g12070 ( 
.A(n_11253),
.B(n_9941),
.Y(n_12070)
);

AND2x2_ASAP7_75t_L g12071 ( 
.A(n_11255),
.B(n_8177),
.Y(n_12071)
);

INVx1_ASAP7_75t_SL g12072 ( 
.A(n_11465),
.Y(n_12072)
);

INVx1_ASAP7_75t_L g12073 ( 
.A(n_11570),
.Y(n_12073)
);

INVx1_ASAP7_75t_L g12074 ( 
.A(n_11530),
.Y(n_12074)
);

AOI22xp5_ASAP7_75t_L g12075 ( 
.A1(n_11300),
.A2(n_7783),
.B1(n_7784),
.B2(n_7777),
.Y(n_12075)
);

INVx3_ASAP7_75t_L g12076 ( 
.A(n_11191),
.Y(n_12076)
);

INVxp67_ASAP7_75t_SL g12077 ( 
.A(n_11191),
.Y(n_12077)
);

INVx1_ASAP7_75t_L g12078 ( 
.A(n_11540),
.Y(n_12078)
);

INVx5_ASAP7_75t_SL g12079 ( 
.A(n_11475),
.Y(n_12079)
);

AND2x2_ASAP7_75t_L g12080 ( 
.A(n_11402),
.B(n_8177),
.Y(n_12080)
);

NAND2xp5_ASAP7_75t_L g12081 ( 
.A(n_11164),
.B(n_8989),
.Y(n_12081)
);

INVx2_ASAP7_75t_L g12082 ( 
.A(n_11525),
.Y(n_12082)
);

INVx2_ASAP7_75t_L g12083 ( 
.A(n_11533),
.Y(n_12083)
);

NAND2xp5_ASAP7_75t_L g12084 ( 
.A(n_11496),
.B(n_8994),
.Y(n_12084)
);

AOI22xp33_ASAP7_75t_L g12085 ( 
.A1(n_11588),
.A2(n_8241),
.B1(n_8454),
.B2(n_8191),
.Y(n_12085)
);

AND2x2_ASAP7_75t_L g12086 ( 
.A(n_11264),
.B(n_8177),
.Y(n_12086)
);

INVx2_ASAP7_75t_L g12087 ( 
.A(n_11535),
.Y(n_12087)
);

INVx1_ASAP7_75t_SL g12088 ( 
.A(n_11520),
.Y(n_12088)
);

INVx5_ASAP7_75t_SL g12089 ( 
.A(n_11487),
.Y(n_12089)
);

NAND2xp5_ASAP7_75t_L g12090 ( 
.A(n_11526),
.B(n_8997),
.Y(n_12090)
);

INVx1_ASAP7_75t_L g12091 ( 
.A(n_11541),
.Y(n_12091)
);

INVx1_ASAP7_75t_L g12092 ( 
.A(n_11542),
.Y(n_12092)
);

INVx1_ASAP7_75t_L g12093 ( 
.A(n_11543),
.Y(n_12093)
);

BUFx2_ASAP7_75t_L g12094 ( 
.A(n_11639),
.Y(n_12094)
);

AND2x2_ASAP7_75t_L g12095 ( 
.A(n_11304),
.B(n_11427),
.Y(n_12095)
);

AND2x2_ASAP7_75t_L g12096 ( 
.A(n_11437),
.B(n_8203),
.Y(n_12096)
);

HB1xp67_ASAP7_75t_L g12097 ( 
.A(n_11640),
.Y(n_12097)
);

NAND2xp5_ASAP7_75t_L g12098 ( 
.A(n_11209),
.B(n_8997),
.Y(n_12098)
);

OR2x2_ASAP7_75t_L g12099 ( 
.A(n_11546),
.B(n_8998),
.Y(n_12099)
);

AND2x2_ASAP7_75t_L g12100 ( 
.A(n_11440),
.B(n_8203),
.Y(n_12100)
);

INVx1_ASAP7_75t_L g12101 ( 
.A(n_11547),
.Y(n_12101)
);

INVx1_ASAP7_75t_L g12102 ( 
.A(n_11548),
.Y(n_12102)
);

AND2x2_ASAP7_75t_L g12103 ( 
.A(n_11444),
.B(n_8203),
.Y(n_12103)
);

AND2x2_ASAP7_75t_L g12104 ( 
.A(n_11459),
.B(n_8219),
.Y(n_12104)
);

INVx5_ASAP7_75t_L g12105 ( 
.A(n_11334),
.Y(n_12105)
);

INVx1_ASAP7_75t_L g12106 ( 
.A(n_11552),
.Y(n_12106)
);

INVx2_ASAP7_75t_L g12107 ( 
.A(n_11480),
.Y(n_12107)
);

OR2x2_ASAP7_75t_L g12108 ( 
.A(n_11555),
.B(n_8998),
.Y(n_12108)
);

AOI22xp33_ASAP7_75t_L g12109 ( 
.A1(n_11225),
.A2(n_8454),
.B1(n_8540),
.B2(n_8191),
.Y(n_12109)
);

NAND2xp5_ASAP7_75t_L g12110 ( 
.A(n_11441),
.B(n_9002),
.Y(n_12110)
);

INVx3_ASAP7_75t_L g12111 ( 
.A(n_11488),
.Y(n_12111)
);

AND2x2_ASAP7_75t_L g12112 ( 
.A(n_11403),
.B(n_8219),
.Y(n_12112)
);

INVx2_ASAP7_75t_L g12113 ( 
.A(n_11323),
.Y(n_12113)
);

AND2x2_ASAP7_75t_L g12114 ( 
.A(n_11409),
.B(n_8219),
.Y(n_12114)
);

CKINVDCx5p33_ASAP7_75t_R g12115 ( 
.A(n_11422),
.Y(n_12115)
);

NAND2xp5_ASAP7_75t_L g12116 ( 
.A(n_11441),
.B(n_9002),
.Y(n_12116)
);

INVx2_ASAP7_75t_L g12117 ( 
.A(n_11327),
.Y(n_12117)
);

INVx2_ASAP7_75t_L g12118 ( 
.A(n_11471),
.Y(n_12118)
);

INVx2_ASAP7_75t_L g12119 ( 
.A(n_11515),
.Y(n_12119)
);

AND2x2_ASAP7_75t_L g12120 ( 
.A(n_11708),
.B(n_8222),
.Y(n_12120)
);

NAND2xp5_ASAP7_75t_L g12121 ( 
.A(n_11527),
.B(n_9004),
.Y(n_12121)
);

INVx1_ASAP7_75t_L g12122 ( 
.A(n_11529),
.Y(n_12122)
);

HB1xp67_ASAP7_75t_L g12123 ( 
.A(n_11646),
.Y(n_12123)
);

AND2x4_ASAP7_75t_L g12124 ( 
.A(n_11421),
.B(n_8119),
.Y(n_12124)
);

AND2x2_ASAP7_75t_L g12125 ( 
.A(n_11531),
.B(n_11431),
.Y(n_12125)
);

NAND2xp5_ASAP7_75t_L g12126 ( 
.A(n_11335),
.B(n_9004),
.Y(n_12126)
);

INVx2_ASAP7_75t_SL g12127 ( 
.A(n_11521),
.Y(n_12127)
);

AND2x2_ASAP7_75t_L g12128 ( 
.A(n_11435),
.B(n_8222),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11607),
.Y(n_12129)
);

OAI211xp5_ASAP7_75t_L g12130 ( 
.A1(n_11186),
.A2(n_11404),
.B(n_11500),
.C(n_11266),
.Y(n_12130)
);

INVx1_ASAP7_75t_L g12131 ( 
.A(n_11330),
.Y(n_12131)
);

OAI21xp33_ASAP7_75t_L g12132 ( 
.A1(n_11461),
.A2(n_9017),
.B(n_9005),
.Y(n_12132)
);

AND2x2_ASAP7_75t_L g12133 ( 
.A(n_11449),
.B(n_8222),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_11331),
.Y(n_12134)
);

INVx2_ASAP7_75t_L g12135 ( 
.A(n_11538),
.Y(n_12135)
);

INVxp67_ASAP7_75t_SL g12136 ( 
.A(n_11428),
.Y(n_12136)
);

INVx2_ASAP7_75t_L g12137 ( 
.A(n_11678),
.Y(n_12137)
);

OAI31xp33_ASAP7_75t_SL g12138 ( 
.A1(n_11222),
.A2(n_7388),
.A3(n_7337),
.B(n_7896),
.Y(n_12138)
);

INVx1_ASAP7_75t_L g12139 ( 
.A(n_11411),
.Y(n_12139)
);

OAI221xp5_ASAP7_75t_L g12140 ( 
.A1(n_11313),
.A2(n_8280),
.B1(n_8418),
.B2(n_8410),
.C(n_8119),
.Y(n_12140)
);

NAND3xp33_ASAP7_75t_L g12141 ( 
.A(n_11616),
.B(n_8280),
.C(n_8119),
.Y(n_12141)
);

OAI21xp5_ASAP7_75t_L g12142 ( 
.A1(n_11293),
.A2(n_7915),
.B(n_7896),
.Y(n_12142)
);

INVx2_ASAP7_75t_L g12143 ( 
.A(n_11694),
.Y(n_12143)
);

AND2x2_ASAP7_75t_L g12144 ( 
.A(n_11569),
.B(n_8222),
.Y(n_12144)
);

AND2x2_ASAP7_75t_L g12145 ( 
.A(n_11711),
.B(n_8228),
.Y(n_12145)
);

AOI22xp33_ASAP7_75t_L g12146 ( 
.A1(n_11648),
.A2(n_8454),
.B1(n_8540),
.B2(n_8191),
.Y(n_12146)
);

AND2x2_ASAP7_75t_L g12147 ( 
.A(n_11655),
.B(n_8228),
.Y(n_12147)
);

AOI211xp5_ASAP7_75t_L g12148 ( 
.A1(n_11256),
.A2(n_8280),
.B(n_8410),
.C(n_8119),
.Y(n_12148)
);

AOI22xp33_ASAP7_75t_L g12149 ( 
.A1(n_11544),
.A2(n_8540),
.B1(n_8721),
.B2(n_8454),
.Y(n_12149)
);

INVx2_ASAP7_75t_SL g12150 ( 
.A(n_11707),
.Y(n_12150)
);

NAND2xp5_ASAP7_75t_L g12151 ( 
.A(n_11381),
.B(n_9005),
.Y(n_12151)
);

NAND2xp5_ASAP7_75t_L g12152 ( 
.A(n_11387),
.B(n_9017),
.Y(n_12152)
);

INVx2_ASAP7_75t_L g12153 ( 
.A(n_11653),
.Y(n_12153)
);

AND2x4_ASAP7_75t_L g12154 ( 
.A(n_11572),
.B(n_8119),
.Y(n_12154)
);

AOI322xp5_ASAP7_75t_L g12155 ( 
.A1(n_11713),
.A2(n_8347),
.A3(n_8218),
.B1(n_8284),
.B2(n_8271),
.C1(n_7372),
.C2(n_7356),
.Y(n_12155)
);

BUFx3_ASAP7_75t_L g12156 ( 
.A(n_11432),
.Y(n_12156)
);

NAND2xp5_ASAP7_75t_L g12157 ( 
.A(n_11433),
.B(n_9019),
.Y(n_12157)
);

AND2x2_ASAP7_75t_L g12158 ( 
.A(n_11362),
.B(n_8228),
.Y(n_12158)
);

INVx2_ASAP7_75t_SL g12159 ( 
.A(n_11654),
.Y(n_12159)
);

AND2x4_ASAP7_75t_L g12160 ( 
.A(n_11657),
.B(n_8280),
.Y(n_12160)
);

AND2x2_ASAP7_75t_L g12161 ( 
.A(n_11366),
.B(n_8228),
.Y(n_12161)
);

INVx1_ASAP7_75t_L g12162 ( 
.A(n_11418),
.Y(n_12162)
);

INVxp67_ASAP7_75t_L g12163 ( 
.A(n_11658),
.Y(n_12163)
);

AOI22xp33_ASAP7_75t_L g12164 ( 
.A1(n_11492),
.A2(n_8540),
.B1(n_8721),
.B2(n_8454),
.Y(n_12164)
);

INVx1_ASAP7_75t_L g12165 ( 
.A(n_11434),
.Y(n_12165)
);

INVx1_ASAP7_75t_L g12166 ( 
.A(n_11436),
.Y(n_12166)
);

INVx2_ASAP7_75t_L g12167 ( 
.A(n_11683),
.Y(n_12167)
);

OAI211xp5_ASAP7_75t_L g12168 ( 
.A1(n_11338),
.A2(n_9786),
.B(n_9499),
.C(n_10254),
.Y(n_12168)
);

AND2x2_ASAP7_75t_L g12169 ( 
.A(n_11371),
.B(n_11377),
.Y(n_12169)
);

INVxp67_ASAP7_75t_SL g12170 ( 
.A(n_11428),
.Y(n_12170)
);

OR2x2_ASAP7_75t_L g12171 ( 
.A(n_11445),
.B(n_9019),
.Y(n_12171)
);

INVx1_ASAP7_75t_L g12172 ( 
.A(n_11477),
.Y(n_12172)
);

AND2x2_ASAP7_75t_L g12173 ( 
.A(n_11378),
.B(n_8228),
.Y(n_12173)
);

OR2x2_ASAP7_75t_L g12174 ( 
.A(n_11333),
.B(n_9020),
.Y(n_12174)
);

OAI31xp33_ASAP7_75t_L g12175 ( 
.A1(n_11332),
.A2(n_8236),
.A3(n_8239),
.B(n_8233),
.Y(n_12175)
);

NAND3xp33_ASAP7_75t_L g12176 ( 
.A(n_11173),
.B(n_8410),
.C(n_8280),
.Y(n_12176)
);

OR2x2_ASAP7_75t_L g12177 ( 
.A(n_11336),
.B(n_9020),
.Y(n_12177)
);

AND2x2_ASAP7_75t_L g12178 ( 
.A(n_11383),
.B(n_8233),
.Y(n_12178)
);

INVx1_ASAP7_75t_L g12179 ( 
.A(n_11484),
.Y(n_12179)
);

OAI21xp33_ASAP7_75t_SL g12180 ( 
.A1(n_11522),
.A2(n_8271),
.B(n_8218),
.Y(n_12180)
);

NAND4xp25_ASAP7_75t_SL g12181 ( 
.A(n_11301),
.B(n_8659),
.C(n_6692),
.D(n_6725),
.Y(n_12181)
);

INVx2_ASAP7_75t_L g12182 ( 
.A(n_11686),
.Y(n_12182)
);

AND2x2_ASAP7_75t_L g12183 ( 
.A(n_11386),
.B(n_8233),
.Y(n_12183)
);

AND2x2_ASAP7_75t_L g12184 ( 
.A(n_11398),
.B(n_8233),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_11688),
.B(n_9283),
.Y(n_12185)
);

INVx2_ASAP7_75t_L g12186 ( 
.A(n_11690),
.Y(n_12186)
);

INVx1_ASAP7_75t_SL g12187 ( 
.A(n_11619),
.Y(n_12187)
);

HB1xp67_ASAP7_75t_L g12188 ( 
.A(n_11620),
.Y(n_12188)
);

OA21x2_ASAP7_75t_L g12189 ( 
.A1(n_11392),
.A2(n_9104),
.B(n_9088),
.Y(n_12189)
);

OAI21xp5_ASAP7_75t_SL g12190 ( 
.A1(n_11280),
.A2(n_11656),
.B(n_11517),
.Y(n_12190)
);

INVx5_ASAP7_75t_SL g12191 ( 
.A(n_11415),
.Y(n_12191)
);

NOR3xp33_ASAP7_75t_SL g12192 ( 
.A(n_11346),
.B(n_7713),
.C(n_7062),
.Y(n_12192)
);

HB1xp67_ASAP7_75t_L g12193 ( 
.A(n_11626),
.Y(n_12193)
);

INVx1_ASAP7_75t_L g12194 ( 
.A(n_11502),
.Y(n_12194)
);

INVx2_ASAP7_75t_L g12195 ( 
.A(n_11695),
.Y(n_12195)
);

AND2x4_ASAP7_75t_SL g12196 ( 
.A(n_11663),
.B(n_7082),
.Y(n_12196)
);

OR2x2_ASAP7_75t_L g12197 ( 
.A(n_11342),
.B(n_9283),
.Y(n_12197)
);

INVx2_ASAP7_75t_L g12198 ( 
.A(n_11697),
.Y(n_12198)
);

AO21x2_ASAP7_75t_L g12199 ( 
.A1(n_11519),
.A2(n_9289),
.B(n_9284),
.Y(n_12199)
);

AND2x4_ASAP7_75t_L g12200 ( 
.A(n_11668),
.B(n_8280),
.Y(n_12200)
);

INVx1_ASAP7_75t_L g12201 ( 
.A(n_11504),
.Y(n_12201)
);

INVx5_ASAP7_75t_L g12202 ( 
.A(n_11649),
.Y(n_12202)
);

HB1xp67_ASAP7_75t_L g12203 ( 
.A(n_11702),
.Y(n_12203)
);

AND2x2_ASAP7_75t_L g12204 ( 
.A(n_11405),
.B(n_8233),
.Y(n_12204)
);

CKINVDCx20_ASAP7_75t_R g12205 ( 
.A(n_11609),
.Y(n_12205)
);

AND2x2_ASAP7_75t_L g12206 ( 
.A(n_11682),
.B(n_8236),
.Y(n_12206)
);

BUFx12f_ASAP7_75t_L g12207 ( 
.A(n_11420),
.Y(n_12207)
);

INVx4_ASAP7_75t_L g12208 ( 
.A(n_11652),
.Y(n_12208)
);

OAI22xp5_ASAP7_75t_SL g12209 ( 
.A1(n_11176),
.A2(n_6719),
.B1(n_7111),
.B2(n_6767),
.Y(n_12209)
);

INVx2_ASAP7_75t_L g12210 ( 
.A(n_11717),
.Y(n_12210)
);

AND2x2_ASAP7_75t_L g12211 ( 
.A(n_11354),
.B(n_8236),
.Y(n_12211)
);

AND2x2_ASAP7_75t_L g12212 ( 
.A(n_11372),
.B(n_8236),
.Y(n_12212)
);

INVx1_ASAP7_75t_L g12213 ( 
.A(n_11512),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_11516),
.Y(n_12214)
);

AND2x4_ASAP7_75t_L g12215 ( 
.A(n_11665),
.B(n_11666),
.Y(n_12215)
);

NAND2xp5_ASAP7_75t_L g12216 ( 
.A(n_11599),
.B(n_9284),
.Y(n_12216)
);

AND2x2_ASAP7_75t_L g12217 ( 
.A(n_11401),
.B(n_8236),
.Y(n_12217)
);

INVx1_ASAP7_75t_L g12218 ( 
.A(n_11344),
.Y(n_12218)
);

AND2x2_ASAP7_75t_L g12219 ( 
.A(n_11498),
.B(n_11564),
.Y(n_12219)
);

OR2x2_ASAP7_75t_L g12220 ( 
.A(n_11350),
.B(n_9289),
.Y(n_12220)
);

INVx2_ASAP7_75t_L g12221 ( 
.A(n_11706),
.Y(n_12221)
);

INVx1_ASAP7_75t_L g12222 ( 
.A(n_11600),
.Y(n_12222)
);

INVx3_ASAP7_75t_L g12223 ( 
.A(n_11352),
.Y(n_12223)
);

AND2x2_ASAP7_75t_L g12224 ( 
.A(n_11679),
.B(n_8239),
.Y(n_12224)
);

AOI211xp5_ASAP7_75t_L g12225 ( 
.A1(n_11341),
.A2(n_8418),
.B(n_8626),
.C(n_8410),
.Y(n_12225)
);

AOI22xp5_ASAP7_75t_L g12226 ( 
.A1(n_11219),
.A2(n_7783),
.B1(n_7784),
.B2(n_7777),
.Y(n_12226)
);

AND2x2_ASAP7_75t_L g12227 ( 
.A(n_11614),
.B(n_8239),
.Y(n_12227)
);

NOR2xp67_ASAP7_75t_SL g12228 ( 
.A(n_11353),
.B(n_7375),
.Y(n_12228)
);

NOR2xp33_ASAP7_75t_SL g12229 ( 
.A(n_11315),
.B(n_7062),
.Y(n_12229)
);

AND2x2_ASAP7_75t_L g12230 ( 
.A(n_11355),
.B(n_8239),
.Y(n_12230)
);

HB1xp67_ASAP7_75t_L g12231 ( 
.A(n_11174),
.Y(n_12231)
);

INVx2_ASAP7_75t_L g12232 ( 
.A(n_11395),
.Y(n_12232)
);

INVx1_ASAP7_75t_L g12233 ( 
.A(n_11605),
.Y(n_12233)
);

OR2x2_ASAP7_75t_L g12234 ( 
.A(n_11610),
.B(n_11613),
.Y(n_12234)
);

AND2x4_ASAP7_75t_L g12235 ( 
.A(n_11720),
.B(n_11518),
.Y(n_12235)
);

INVx2_ASAP7_75t_SL g12236 ( 
.A(n_11511),
.Y(n_12236)
);

AND2x2_ASAP7_75t_L g12237 ( 
.A(n_11632),
.B(n_8239),
.Y(n_12237)
);

AOI22xp33_ASAP7_75t_L g12238 ( 
.A1(n_11233),
.A2(n_8540),
.B1(n_8721),
.B2(n_8454),
.Y(n_12238)
);

AND2x2_ASAP7_75t_L g12239 ( 
.A(n_11618),
.B(n_8256),
.Y(n_12239)
);

NAND2xp5_ASAP7_75t_L g12240 ( 
.A(n_11684),
.B(n_9291),
.Y(n_12240)
);

AND2x2_ASAP7_75t_L g12241 ( 
.A(n_11721),
.B(n_11735),
.Y(n_12241)
);

AND2x4_ASAP7_75t_SL g12242 ( 
.A(n_11733),
.B(n_6750),
.Y(n_12242)
);

AND2x2_ASAP7_75t_L g12243 ( 
.A(n_11721),
.B(n_11701),
.Y(n_12243)
);

AND2x2_ASAP7_75t_L g12244 ( 
.A(n_11741),
.B(n_11594),
.Y(n_12244)
);

INVx1_ASAP7_75t_L g12245 ( 
.A(n_11765),
.Y(n_12245)
);

AND2x2_ASAP7_75t_L g12246 ( 
.A(n_11860),
.B(n_11423),
.Y(n_12246)
);

AND2x2_ASAP7_75t_L g12247 ( 
.A(n_11736),
.B(n_11523),
.Y(n_12247)
);

INVx1_ASAP7_75t_L g12248 ( 
.A(n_11770),
.Y(n_12248)
);

NOR2x1_ASAP7_75t_L g12249 ( 
.A(n_11975),
.B(n_11311),
.Y(n_12249)
);

BUFx2_ASAP7_75t_L g12250 ( 
.A(n_11775),
.Y(n_12250)
);

INVx1_ASAP7_75t_L g12251 ( 
.A(n_11889),
.Y(n_12251)
);

AND2x2_ASAP7_75t_L g12252 ( 
.A(n_11779),
.B(n_11396),
.Y(n_12252)
);

INVx1_ASAP7_75t_L g12253 ( 
.A(n_11782),
.Y(n_12253)
);

HB1xp67_ASAP7_75t_L g12254 ( 
.A(n_11919),
.Y(n_12254)
);

INVx2_ASAP7_75t_SL g12255 ( 
.A(n_12105),
.Y(n_12255)
);

AND2x2_ASAP7_75t_L g12256 ( 
.A(n_11799),
.B(n_11597),
.Y(n_12256)
);

AND2x2_ASAP7_75t_L g12257 ( 
.A(n_11806),
.B(n_11814),
.Y(n_12257)
);

OR2x2_ASAP7_75t_L g12258 ( 
.A(n_11722),
.B(n_11660),
.Y(n_12258)
);

INVx2_ASAP7_75t_SL g12259 ( 
.A(n_12105),
.Y(n_12259)
);

OR2x2_ASAP7_75t_L g12260 ( 
.A(n_11743),
.B(n_11416),
.Y(n_12260)
);

AND2x2_ASAP7_75t_L g12261 ( 
.A(n_11793),
.B(n_11532),
.Y(n_12261)
);

OR2x2_ASAP7_75t_L g12262 ( 
.A(n_11737),
.B(n_11360),
.Y(n_12262)
);

HB1xp67_ASAP7_75t_L g12263 ( 
.A(n_11813),
.Y(n_12263)
);

INVx2_ASAP7_75t_L g12264 ( 
.A(n_12105),
.Y(n_12264)
);

NAND2xp5_ASAP7_75t_L g12265 ( 
.A(n_11729),
.B(n_11691),
.Y(n_12265)
);

AND2x2_ASAP7_75t_L g12266 ( 
.A(n_11725),
.B(n_11481),
.Y(n_12266)
);

NAND2xp5_ASAP7_75t_L g12267 ( 
.A(n_11734),
.B(n_11602),
.Y(n_12267)
);

INVx1_ASAP7_75t_L g12268 ( 
.A(n_11780),
.Y(n_12268)
);

NAND2xp5_ASAP7_75t_L g12269 ( 
.A(n_11838),
.B(n_11608),
.Y(n_12269)
);

OR2x2_ASAP7_75t_L g12270 ( 
.A(n_11745),
.B(n_11361),
.Y(n_12270)
);

INVx1_ASAP7_75t_L g12271 ( 
.A(n_11731),
.Y(n_12271)
);

OR2x2_ASAP7_75t_L g12272 ( 
.A(n_11763),
.B(n_11696),
.Y(n_12272)
);

INVx1_ASAP7_75t_L g12273 ( 
.A(n_11731),
.Y(n_12273)
);

NAND2xp5_ASAP7_75t_L g12274 ( 
.A(n_11991),
.B(n_11625),
.Y(n_12274)
);

NAND2xp5_ASAP7_75t_L g12275 ( 
.A(n_11895),
.B(n_11628),
.Y(n_12275)
);

INVxp67_ASAP7_75t_L g12276 ( 
.A(n_11961),
.Y(n_12276)
);

NAND2xp5_ASAP7_75t_L g12277 ( 
.A(n_11895),
.B(n_11659),
.Y(n_12277)
);

INVx2_ASAP7_75t_L g12278 ( 
.A(n_11827),
.Y(n_12278)
);

INVx1_ASAP7_75t_L g12279 ( 
.A(n_11739),
.Y(n_12279)
);

NAND2xp5_ASAP7_75t_L g12280 ( 
.A(n_11751),
.B(n_11692),
.Y(n_12280)
);

INVx2_ASAP7_75t_L g12281 ( 
.A(n_11775),
.Y(n_12281)
);

AND2x2_ASAP7_75t_L g12282 ( 
.A(n_11748),
.B(n_11468),
.Y(n_12282)
);

NOR2xp33_ASAP7_75t_SL g12283 ( 
.A(n_11733),
.B(n_11580),
.Y(n_12283)
);

INVx1_ASAP7_75t_L g12284 ( 
.A(n_11739),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_11747),
.Y(n_12285)
);

AND2x2_ASAP7_75t_L g12286 ( 
.A(n_11807),
.B(n_11593),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_11747),
.Y(n_12287)
);

NOR2xp33_ASAP7_75t_L g12288 ( 
.A(n_11837),
.B(n_11373),
.Y(n_12288)
);

INVx2_ASAP7_75t_L g12289 ( 
.A(n_11777),
.Y(n_12289)
);

INVxp67_ASAP7_75t_L g12290 ( 
.A(n_11961),
.Y(n_12290)
);

INVx1_ASAP7_75t_L g12291 ( 
.A(n_11824),
.Y(n_12291)
);

AND2x2_ASAP7_75t_L g12292 ( 
.A(n_11828),
.B(n_11693),
.Y(n_12292)
);

INVx2_ASAP7_75t_SL g12293 ( 
.A(n_11777),
.Y(n_12293)
);

AND2x2_ASAP7_75t_L g12294 ( 
.A(n_11819),
.B(n_11700),
.Y(n_12294)
);

AND2x2_ASAP7_75t_L g12295 ( 
.A(n_11832),
.B(n_11479),
.Y(n_12295)
);

INVx1_ASAP7_75t_L g12296 ( 
.A(n_11829),
.Y(n_12296)
);

NAND2xp5_ASAP7_75t_L g12297 ( 
.A(n_11764),
.B(n_12111),
.Y(n_12297)
);

NAND2xp5_ASAP7_75t_L g12298 ( 
.A(n_12111),
.B(n_11388),
.Y(n_12298)
);

HB1xp67_ASAP7_75t_L g12299 ( 
.A(n_11797),
.Y(n_12299)
);

AND2x2_ASAP7_75t_L g12300 ( 
.A(n_11868),
.B(n_11369),
.Y(n_12300)
);

OR2x2_ASAP7_75t_L g12301 ( 
.A(n_11727),
.B(n_11673),
.Y(n_12301)
);

NAND2xp5_ASAP7_75t_L g12302 ( 
.A(n_11926),
.B(n_11374),
.Y(n_12302)
);

OR2x2_ASAP7_75t_L g12303 ( 
.A(n_11974),
.B(n_11483),
.Y(n_12303)
);

OR2x2_ASAP7_75t_L g12304 ( 
.A(n_11851),
.B(n_11290),
.Y(n_12304)
);

AND2x2_ASAP7_75t_L g12305 ( 
.A(n_11871),
.B(n_11297),
.Y(n_12305)
);

NAND2xp5_ASAP7_75t_L g12306 ( 
.A(n_11931),
.B(n_11419),
.Y(n_12306)
);

INVx1_ASAP7_75t_L g12307 ( 
.A(n_11831),
.Y(n_12307)
);

INVx1_ASAP7_75t_L g12308 ( 
.A(n_11834),
.Y(n_12308)
);

INVx2_ASAP7_75t_SL g12309 ( 
.A(n_11817),
.Y(n_12309)
);

INVx1_ASAP7_75t_L g12310 ( 
.A(n_11839),
.Y(n_12310)
);

BUFx2_ASAP7_75t_L g12311 ( 
.A(n_11817),
.Y(n_12311)
);

NAND2xp5_ASAP7_75t_L g12312 ( 
.A(n_11934),
.B(n_11473),
.Y(n_12312)
);

INVx1_ASAP7_75t_L g12313 ( 
.A(n_11847),
.Y(n_12313)
);

NAND2xp5_ASAP7_75t_L g12314 ( 
.A(n_11896),
.B(n_11497),
.Y(n_12314)
);

OR2x2_ASAP7_75t_L g12315 ( 
.A(n_11884),
.B(n_11408),
.Y(n_12315)
);

INVx1_ASAP7_75t_L g12316 ( 
.A(n_11783),
.Y(n_12316)
);

OR2x2_ASAP7_75t_L g12317 ( 
.A(n_11859),
.B(n_11410),
.Y(n_12317)
);

INVx1_ASAP7_75t_L g12318 ( 
.A(n_12203),
.Y(n_12318)
);

INVx1_ASAP7_75t_L g12319 ( 
.A(n_11938),
.Y(n_12319)
);

INVx1_ASAP7_75t_L g12320 ( 
.A(n_12020),
.Y(n_12320)
);

HB1xp67_ASAP7_75t_L g12321 ( 
.A(n_11982),
.Y(n_12321)
);

AND2x2_ASAP7_75t_L g12322 ( 
.A(n_11795),
.B(n_11294),
.Y(n_12322)
);

AND2x2_ASAP7_75t_L g12323 ( 
.A(n_11894),
.B(n_11837),
.Y(n_12323)
);

HB1xp67_ASAP7_75t_L g12324 ( 
.A(n_11925),
.Y(n_12324)
);

NAND2xp5_ASAP7_75t_L g12325 ( 
.A(n_11932),
.B(n_11615),
.Y(n_12325)
);

AND2x4_ASAP7_75t_L g12326 ( 
.A(n_11732),
.B(n_8410),
.Y(n_12326)
);

OR2x2_ASAP7_75t_L g12327 ( 
.A(n_11757),
.B(n_11391),
.Y(n_12327)
);

AND2x2_ASAP7_75t_L g12328 ( 
.A(n_11815),
.B(n_8271),
.Y(n_12328)
);

BUFx2_ASAP7_75t_L g12329 ( 
.A(n_11732),
.Y(n_12329)
);

AND2x4_ASAP7_75t_L g12330 ( 
.A(n_11781),
.B(n_11864),
.Y(n_12330)
);

INVx2_ASAP7_75t_L g12331 ( 
.A(n_11746),
.Y(n_12331)
);

AND2x4_ASAP7_75t_L g12332 ( 
.A(n_11781),
.B(n_8410),
.Y(n_12332)
);

AND2x2_ASAP7_75t_L g12333 ( 
.A(n_11863),
.B(n_8284),
.Y(n_12333)
);

INVx1_ASAP7_75t_L g12334 ( 
.A(n_12033),
.Y(n_12334)
);

INVx1_ASAP7_75t_L g12335 ( 
.A(n_12041),
.Y(n_12335)
);

INVx2_ASAP7_75t_L g12336 ( 
.A(n_11879),
.Y(n_12336)
);

INVx2_ASAP7_75t_L g12337 ( 
.A(n_11879),
.Y(n_12337)
);

INVx1_ASAP7_75t_L g12338 ( 
.A(n_12050),
.Y(n_12338)
);

HB1xp67_ASAP7_75t_L g12339 ( 
.A(n_11906),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_L g12340 ( 
.A(n_11773),
.B(n_11676),
.Y(n_12340)
);

NAND2xp5_ASAP7_75t_L g12341 ( 
.A(n_12095),
.B(n_11676),
.Y(n_12341)
);

INVx1_ASAP7_75t_L g12342 ( 
.A(n_12067),
.Y(n_12342)
);

NAND2xp5_ASAP7_75t_L g12343 ( 
.A(n_11972),
.B(n_11345),
.Y(n_12343)
);

INVx2_ASAP7_75t_L g12344 ( 
.A(n_11879),
.Y(n_12344)
);

OR3x2_ASAP7_75t_L g12345 ( 
.A(n_12234),
.B(n_7964),
.C(n_6974),
.Y(n_12345)
);

INVx3_ASAP7_75t_L g12346 ( 
.A(n_11762),
.Y(n_12346)
);

NAND2xp5_ASAP7_75t_L g12347 ( 
.A(n_11935),
.B(n_11322),
.Y(n_12347)
);

AND2x4_ASAP7_75t_L g12348 ( 
.A(n_11864),
.B(n_8418),
.Y(n_12348)
);

NAND2xp5_ASAP7_75t_L g12349 ( 
.A(n_11940),
.B(n_11289),
.Y(n_12349)
);

AND2x2_ASAP7_75t_L g12350 ( 
.A(n_11877),
.B(n_8284),
.Y(n_12350)
);

INVx2_ASAP7_75t_L g12351 ( 
.A(n_11785),
.Y(n_12351)
);

NAND2xp5_ASAP7_75t_L g12352 ( 
.A(n_11893),
.B(n_11292),
.Y(n_12352)
);

OR2x2_ASAP7_75t_L g12353 ( 
.A(n_11738),
.B(n_11358),
.Y(n_12353)
);

OR2x2_ASAP7_75t_L g12354 ( 
.A(n_11950),
.B(n_11464),
.Y(n_12354)
);

AOI21xp5_ASAP7_75t_L g12355 ( 
.A1(n_12012),
.A2(n_11439),
.B(n_11430),
.Y(n_12355)
);

NOR2xp67_ASAP7_75t_L g12356 ( 
.A(n_11844),
.B(n_11647),
.Y(n_12356)
);

AND2x2_ASAP7_75t_L g12357 ( 
.A(n_11902),
.B(n_8347),
.Y(n_12357)
);

INVx1_ASAP7_75t_L g12358 ( 
.A(n_12097),
.Y(n_12358)
);

NOR2x1_ASAP7_75t_L g12359 ( 
.A(n_12076),
.B(n_11562),
.Y(n_12359)
);

INVx1_ASAP7_75t_L g12360 ( 
.A(n_12123),
.Y(n_12360)
);

INVx2_ASAP7_75t_L g12361 ( 
.A(n_11843),
.Y(n_12361)
);

NOR2x1_ASAP7_75t_L g12362 ( 
.A(n_12076),
.B(n_11562),
.Y(n_12362)
);

NAND2xp5_ASAP7_75t_L g12363 ( 
.A(n_11776),
.B(n_9291),
.Y(n_12363)
);

AND2x4_ASAP7_75t_SL g12364 ( 
.A(n_11820),
.B(n_6783),
.Y(n_12364)
);

INVx1_ASAP7_75t_L g12365 ( 
.A(n_11918),
.Y(n_12365)
);

AND2x2_ASAP7_75t_L g12366 ( 
.A(n_12000),
.B(n_8347),
.Y(n_12366)
);

NOR2x1_ASAP7_75t_L g12367 ( 
.A(n_11956),
.B(n_11970),
.Y(n_12367)
);

HB1xp67_ASAP7_75t_L g12368 ( 
.A(n_11921),
.Y(n_12368)
);

AND2x2_ASAP7_75t_L g12369 ( 
.A(n_12035),
.B(n_9294),
.Y(n_12369)
);

NAND2x1p5_ASAP7_75t_L g12370 ( 
.A(n_11844),
.B(n_7240),
.Y(n_12370)
);

AND2x2_ASAP7_75t_SL g12371 ( 
.A(n_11875),
.B(n_7240),
.Y(n_12371)
);

HB1xp67_ASAP7_75t_L g12372 ( 
.A(n_12202),
.Y(n_12372)
);

NAND2xp5_ASAP7_75t_L g12373 ( 
.A(n_11760),
.B(n_9294),
.Y(n_12373)
);

AND2x4_ASAP7_75t_L g12374 ( 
.A(n_11762),
.B(n_8418),
.Y(n_12374)
);

AND2x2_ASAP7_75t_L g12375 ( 
.A(n_11786),
.B(n_9300),
.Y(n_12375)
);

INVx1_ASAP7_75t_L g12376 ( 
.A(n_11983),
.Y(n_12376)
);

NAND2xp5_ASAP7_75t_L g12377 ( 
.A(n_11796),
.B(n_9300),
.Y(n_12377)
);

NAND2xp5_ASAP7_75t_L g12378 ( 
.A(n_11726),
.B(n_9302),
.Y(n_12378)
);

NOR2xp33_ASAP7_75t_L g12379 ( 
.A(n_11958),
.B(n_11917),
.Y(n_12379)
);

NAND2xp5_ASAP7_75t_L g12380 ( 
.A(n_11990),
.B(n_9302),
.Y(n_12380)
);

AND2x4_ASAP7_75t_L g12381 ( 
.A(n_11866),
.B(n_8418),
.Y(n_12381)
);

AND2x2_ASAP7_75t_L g12382 ( 
.A(n_11790),
.B(n_9304),
.Y(n_12382)
);

HB1xp67_ASAP7_75t_L g12383 ( 
.A(n_12202),
.Y(n_12383)
);

INVx2_ASAP7_75t_L g12384 ( 
.A(n_12034),
.Y(n_12384)
);

OAI22xp33_ASAP7_75t_SL g12385 ( 
.A1(n_11794),
.A2(n_11592),
.B1(n_7783),
.B2(n_7784),
.Y(n_12385)
);

CKINVDCx5p33_ASAP7_75t_R g12386 ( 
.A(n_11930),
.Y(n_12386)
);

INVx4_ASAP7_75t_L g12387 ( 
.A(n_11973),
.Y(n_12387)
);

NAND2xp5_ASAP7_75t_L g12388 ( 
.A(n_12001),
.B(n_9304),
.Y(n_12388)
);

AND2x4_ASAP7_75t_SL g12389 ( 
.A(n_11818),
.B(n_7410),
.Y(n_12389)
);

NAND2xp5_ASAP7_75t_L g12390 ( 
.A(n_11885),
.B(n_9308),
.Y(n_12390)
);

AND2x2_ASAP7_75t_L g12391 ( 
.A(n_11941),
.B(n_9308),
.Y(n_12391)
);

NAND2xp5_ASAP7_75t_L g12392 ( 
.A(n_11857),
.B(n_9313),
.Y(n_12392)
);

BUFx2_ASAP7_75t_L g12393 ( 
.A(n_12023),
.Y(n_12393)
);

INVxp67_ASAP7_75t_SL g12394 ( 
.A(n_11956),
.Y(n_12394)
);

INVx1_ASAP7_75t_L g12395 ( 
.A(n_11992),
.Y(n_12395)
);

AND2x2_ASAP7_75t_L g12396 ( 
.A(n_11929),
.B(n_9313),
.Y(n_12396)
);

NAND2xp5_ASAP7_75t_L g12397 ( 
.A(n_11959),
.B(n_11771),
.Y(n_12397)
);

AND2x2_ASAP7_75t_L g12398 ( 
.A(n_11993),
.B(n_9315),
.Y(n_12398)
);

INVxp67_ASAP7_75t_L g12399 ( 
.A(n_12029),
.Y(n_12399)
);

INVx1_ASAP7_75t_L g12400 ( 
.A(n_11913),
.Y(n_12400)
);

OR2x2_ASAP7_75t_L g12401 ( 
.A(n_11900),
.B(n_11464),
.Y(n_12401)
);

NAND2xp5_ASAP7_75t_L g12402 ( 
.A(n_12127),
.B(n_9315),
.Y(n_12402)
);

AND2x4_ASAP7_75t_L g12403 ( 
.A(n_11842),
.B(n_8418),
.Y(n_12403)
);

INVxp67_ASAP7_75t_L g12404 ( 
.A(n_11744),
.Y(n_12404)
);

AND2x2_ASAP7_75t_L g12405 ( 
.A(n_11993),
.B(n_9318),
.Y(n_12405)
);

INVx1_ASAP7_75t_L g12406 ( 
.A(n_11922),
.Y(n_12406)
);

INVxp67_ASAP7_75t_L g12407 ( 
.A(n_11749),
.Y(n_12407)
);

AND2x2_ASAP7_75t_L g12408 ( 
.A(n_11849),
.B(n_9318),
.Y(n_12408)
);

AND2x2_ASAP7_75t_L g12409 ( 
.A(n_11899),
.B(n_9319),
.Y(n_12409)
);

INVx1_ASAP7_75t_L g12410 ( 
.A(n_11756),
.Y(n_12410)
);

AND2x4_ASAP7_75t_L g12411 ( 
.A(n_11842),
.B(n_8418),
.Y(n_12411)
);

NAND2xp5_ASAP7_75t_L g12412 ( 
.A(n_11778),
.B(n_9319),
.Y(n_12412)
);

AND2x2_ASAP7_75t_L g12413 ( 
.A(n_12048),
.B(n_9320),
.Y(n_12413)
);

INVx1_ASAP7_75t_L g12414 ( 
.A(n_11758),
.Y(n_12414)
);

AND2x2_ASAP7_75t_L g12415 ( 
.A(n_12052),
.B(n_9320),
.Y(n_12415)
);

OR2x2_ASAP7_75t_L g12416 ( 
.A(n_11901),
.B(n_11443),
.Y(n_12416)
);

INVx1_ASAP7_75t_L g12417 ( 
.A(n_11759),
.Y(n_12417)
);

INVx2_ASAP7_75t_L g12418 ( 
.A(n_12034),
.Y(n_12418)
);

INVx1_ASAP7_75t_SL g12419 ( 
.A(n_11872),
.Y(n_12419)
);

AND2x2_ASAP7_75t_L g12420 ( 
.A(n_11911),
.B(n_9326),
.Y(n_12420)
);

AND2x2_ASAP7_75t_L g12421 ( 
.A(n_11920),
.B(n_9326),
.Y(n_12421)
);

NOR3xp33_ASAP7_75t_L g12422 ( 
.A(n_11946),
.B(n_11439),
.C(n_11430),
.Y(n_12422)
);

OR2x2_ASAP7_75t_L g12423 ( 
.A(n_11904),
.B(n_11443),
.Y(n_12423)
);

INVx2_ASAP7_75t_SL g12424 ( 
.A(n_12202),
.Y(n_12424)
);

INVx1_ASAP7_75t_SL g12425 ( 
.A(n_11886),
.Y(n_12425)
);

INVx1_ASAP7_75t_L g12426 ( 
.A(n_11873),
.Y(n_12426)
);

INVx2_ASAP7_75t_SL g12427 ( 
.A(n_11865),
.Y(n_12427)
);

NAND2xp5_ASAP7_75t_L g12428 ( 
.A(n_11788),
.B(n_9331),
.Y(n_12428)
);

NAND2xp5_ASAP7_75t_L g12429 ( 
.A(n_11939),
.B(n_9331),
.Y(n_12429)
);

OR2x2_ASAP7_75t_L g12430 ( 
.A(n_11928),
.B(n_11563),
.Y(n_12430)
);

INVx3_ASAP7_75t_L g12431 ( 
.A(n_11973),
.Y(n_12431)
);

INVx1_ASAP7_75t_L g12432 ( 
.A(n_11962),
.Y(n_12432)
);

INVx3_ASAP7_75t_L g12433 ( 
.A(n_12037),
.Y(n_12433)
);

AND2x4_ASAP7_75t_L g12434 ( 
.A(n_11865),
.B(n_8626),
.Y(n_12434)
);

HB1xp67_ASAP7_75t_L g12435 ( 
.A(n_12013),
.Y(n_12435)
);

AND2x2_ASAP7_75t_L g12436 ( 
.A(n_11883),
.B(n_9335),
.Y(n_12436)
);

OAI21xp5_ASAP7_75t_SL g12437 ( 
.A1(n_11833),
.A2(n_11565),
.B(n_11563),
.Y(n_12437)
);

OAI22xp5_ASAP7_75t_SL g12438 ( 
.A1(n_11888),
.A2(n_11601),
.B1(n_11565),
.B2(n_8626),
.Y(n_12438)
);

NAND2xp5_ASAP7_75t_L g12439 ( 
.A(n_11949),
.B(n_9335),
.Y(n_12439)
);

AND2x2_ASAP7_75t_L g12440 ( 
.A(n_12191),
.B(n_9348),
.Y(n_12440)
);

AND2x2_ASAP7_75t_L g12441 ( 
.A(n_12191),
.B(n_11854),
.Y(n_12441)
);

INVx1_ASAP7_75t_L g12442 ( 
.A(n_12002),
.Y(n_12442)
);

AND2x2_ASAP7_75t_L g12443 ( 
.A(n_11861),
.B(n_9348),
.Y(n_12443)
);

AND2x2_ASAP7_75t_L g12444 ( 
.A(n_11867),
.B(n_9349),
.Y(n_12444)
);

NAND2xp5_ASAP7_75t_SL g12445 ( 
.A(n_11826),
.B(n_8626),
.Y(n_12445)
);

AND2x2_ASAP7_75t_L g12446 ( 
.A(n_11876),
.B(n_11890),
.Y(n_12446)
);

AND2x2_ASAP7_75t_L g12447 ( 
.A(n_12045),
.B(n_9349),
.Y(n_12447)
);

NAND2xp5_ASAP7_75t_L g12448 ( 
.A(n_11730),
.B(n_9350),
.Y(n_12448)
);

AND2x4_ASAP7_75t_L g12449 ( 
.A(n_11914),
.B(n_11954),
.Y(n_12449)
);

AND2x2_ASAP7_75t_L g12450 ( 
.A(n_11963),
.B(n_9350),
.Y(n_12450)
);

INVx2_ASAP7_75t_L g12451 ( 
.A(n_12079),
.Y(n_12451)
);

INVx1_ASAP7_75t_L g12452 ( 
.A(n_12006),
.Y(n_12452)
);

OR2x2_ASAP7_75t_L g12453 ( 
.A(n_11937),
.B(n_11601),
.Y(n_12453)
);

AND2x2_ASAP7_75t_L g12454 ( 
.A(n_11953),
.B(n_9351),
.Y(n_12454)
);

AND2x2_ASAP7_75t_L g12455 ( 
.A(n_12113),
.B(n_9351),
.Y(n_12455)
);

AND2x2_ASAP7_75t_L g12456 ( 
.A(n_12117),
.B(n_9355),
.Y(n_12456)
);

OR2x2_ASAP7_75t_L g12457 ( 
.A(n_11822),
.B(n_9355),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_11848),
.Y(n_12458)
);

NAND2xp5_ASAP7_75t_L g12459 ( 
.A(n_11933),
.B(n_9358),
.Y(n_12459)
);

OR2x2_ASAP7_75t_L g12460 ( 
.A(n_11803),
.B(n_9358),
.Y(n_12460)
);

AND2x2_ASAP7_75t_L g12461 ( 
.A(n_11957),
.B(n_9360),
.Y(n_12461)
);

BUFx2_ASAP7_75t_L g12462 ( 
.A(n_12019),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_11970),
.Y(n_12463)
);

INVx1_ASAP7_75t_L g12464 ( 
.A(n_11995),
.Y(n_12464)
);

INVx1_ASAP7_75t_L g12465 ( 
.A(n_11998),
.Y(n_12465)
);

OR2x2_ASAP7_75t_L g12466 ( 
.A(n_11825),
.B(n_11916),
.Y(n_12466)
);

AND2x2_ASAP7_75t_L g12467 ( 
.A(n_12015),
.B(n_9360),
.Y(n_12467)
);

INVx3_ASAP7_75t_R g12468 ( 
.A(n_12221),
.Y(n_12468)
);

INVx1_ASAP7_75t_L g12469 ( 
.A(n_11723),
.Y(n_12469)
);

INVxp67_ASAP7_75t_SL g12470 ( 
.A(n_11891),
.Y(n_12470)
);

INVx1_ASAP7_75t_L g12471 ( 
.A(n_11728),
.Y(n_12471)
);

OR2x2_ASAP7_75t_L g12472 ( 
.A(n_11915),
.B(n_9366),
.Y(n_12472)
);

OR2x2_ASAP7_75t_L g12473 ( 
.A(n_12068),
.B(n_9366),
.Y(n_12473)
);

INVx1_ASAP7_75t_L g12474 ( 
.A(n_12037),
.Y(n_12474)
);

NAND2xp5_ASAP7_75t_L g12475 ( 
.A(n_12055),
.B(n_9372),
.Y(n_12475)
);

NAND2xp5_ASAP7_75t_L g12476 ( 
.A(n_12150),
.B(n_9372),
.Y(n_12476)
);

AND2x2_ASAP7_75t_L g12477 ( 
.A(n_12031),
.B(n_9379),
.Y(n_12477)
);

OR2x2_ASAP7_75t_L g12478 ( 
.A(n_11750),
.B(n_9379),
.Y(n_12478)
);

NAND2x1p5_ASAP7_75t_L g12479 ( 
.A(n_11986),
.B(n_7240),
.Y(n_12479)
);

INVx1_ASAP7_75t_L g12480 ( 
.A(n_12060),
.Y(n_12480)
);

AND2x2_ASAP7_75t_L g12481 ( 
.A(n_12042),
.B(n_9391),
.Y(n_12481)
);

OR2x2_ASAP7_75t_L g12482 ( 
.A(n_11753),
.B(n_9391),
.Y(n_12482)
);

OR2x2_ASAP7_75t_L g12483 ( 
.A(n_11909),
.B(n_9392),
.Y(n_12483)
);

AND2x2_ASAP7_75t_L g12484 ( 
.A(n_12051),
.B(n_9392),
.Y(n_12484)
);

OR2x2_ASAP7_75t_L g12485 ( 
.A(n_11850),
.B(n_9394),
.Y(n_12485)
);

OR2x2_ASAP7_75t_L g12486 ( 
.A(n_11850),
.B(n_9394),
.Y(n_12486)
);

AND2x2_ASAP7_75t_L g12487 ( 
.A(n_12064),
.B(n_9405),
.Y(n_12487)
);

HB1xp67_ASAP7_75t_L g12488 ( 
.A(n_11969),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_12060),
.Y(n_12489)
);

AND2x2_ASAP7_75t_L g12490 ( 
.A(n_12082),
.B(n_12083),
.Y(n_12490)
);

INVx2_ASAP7_75t_L g12491 ( 
.A(n_12079),
.Y(n_12491)
);

AND2x2_ASAP7_75t_L g12492 ( 
.A(n_12087),
.B(n_9405),
.Y(n_12492)
);

INVx2_ASAP7_75t_L g12493 ( 
.A(n_12089),
.Y(n_12493)
);

AND2x2_ASAP7_75t_L g12494 ( 
.A(n_12107),
.B(n_9407),
.Y(n_12494)
);

NAND2xp5_ASAP7_75t_L g12495 ( 
.A(n_11810),
.B(n_9407),
.Y(n_12495)
);

HB1xp67_ASAP7_75t_L g12496 ( 
.A(n_11977),
.Y(n_12496)
);

INVx1_ASAP7_75t_L g12497 ( 
.A(n_11881),
.Y(n_12497)
);

OR2x2_ASAP7_75t_L g12498 ( 
.A(n_11789),
.B(n_11809),
.Y(n_12498)
);

INVx1_ASAP7_75t_L g12499 ( 
.A(n_12058),
.Y(n_12499)
);

INVx1_ASAP7_75t_L g12500 ( 
.A(n_12094),
.Y(n_12500)
);

NAND2xp5_ASAP7_75t_L g12501 ( 
.A(n_11985),
.B(n_9408),
.Y(n_12501)
);

INVx1_ASAP7_75t_SL g12502 ( 
.A(n_11943),
.Y(n_12502)
);

AND2x2_ASAP7_75t_L g12503 ( 
.A(n_11945),
.B(n_9408),
.Y(n_12503)
);

AND2x2_ASAP7_75t_L g12504 ( 
.A(n_11823),
.B(n_12018),
.Y(n_12504)
);

OR2x2_ASAP7_75t_L g12505 ( 
.A(n_11984),
.B(n_11980),
.Y(n_12505)
);

OR2x2_ASAP7_75t_L g12506 ( 
.A(n_12043),
.B(n_9411),
.Y(n_12506)
);

NOR2xp67_ASAP7_75t_SL g12507 ( 
.A(n_11966),
.B(n_8626),
.Y(n_12507)
);

NAND2xp5_ASAP7_75t_SL g12508 ( 
.A(n_12022),
.B(n_8626),
.Y(n_12508)
);

INVx1_ASAP7_75t_L g12509 ( 
.A(n_12188),
.Y(n_12509)
);

INVx3_ASAP7_75t_R g12510 ( 
.A(n_12017),
.Y(n_12510)
);

AND2x2_ASAP7_75t_L g12511 ( 
.A(n_11792),
.B(n_9411),
.Y(n_12511)
);

INVx2_ASAP7_75t_L g12512 ( 
.A(n_12089),
.Y(n_12512)
);

INVx2_ASAP7_75t_L g12513 ( 
.A(n_12021),
.Y(n_12513)
);

INVx1_ASAP7_75t_L g12514 ( 
.A(n_12193),
.Y(n_12514)
);

AND2x2_ASAP7_75t_L g12515 ( 
.A(n_12239),
.B(n_9414),
.Y(n_12515)
);

NAND2xp5_ASAP7_75t_L g12516 ( 
.A(n_11755),
.B(n_9414),
.Y(n_12516)
);

AND2x2_ASAP7_75t_L g12517 ( 
.A(n_12027),
.B(n_9417),
.Y(n_12517)
);

AND2x2_ASAP7_75t_L g12518 ( 
.A(n_12027),
.B(n_9417),
.Y(n_12518)
);

INVx1_ASAP7_75t_L g12519 ( 
.A(n_12136),
.Y(n_12519)
);

INVx1_ASAP7_75t_L g12520 ( 
.A(n_12170),
.Y(n_12520)
);

NAND2xp5_ASAP7_75t_L g12521 ( 
.A(n_11754),
.B(n_9420),
.Y(n_12521)
);

AND2x2_ASAP7_75t_L g12522 ( 
.A(n_11802),
.B(n_9420),
.Y(n_12522)
);

AND2x2_ASAP7_75t_L g12523 ( 
.A(n_12237),
.B(n_9425),
.Y(n_12523)
);

AND2x2_ASAP7_75t_L g12524 ( 
.A(n_12227),
.B(n_12125),
.Y(n_12524)
);

NOR2xp33_ASAP7_75t_L g12525 ( 
.A(n_11740),
.B(n_7313),
.Y(n_12525)
);

OR2x2_ASAP7_75t_L g12526 ( 
.A(n_12069),
.B(n_9425),
.Y(n_12526)
);

AND2x2_ASAP7_75t_L g12527 ( 
.A(n_12025),
.B(n_9426),
.Y(n_12527)
);

AND2x4_ASAP7_75t_L g12528 ( 
.A(n_12159),
.B(n_8626),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_12185),
.Y(n_12529)
);

NAND2xp5_ASAP7_75t_L g12530 ( 
.A(n_11845),
.B(n_9426),
.Y(n_12530)
);

AND2x2_ASAP7_75t_L g12531 ( 
.A(n_12219),
.B(n_9435),
.Y(n_12531)
);

INVx1_ASAP7_75t_L g12532 ( 
.A(n_12047),
.Y(n_12532)
);

NAND2xp5_ASAP7_75t_L g12533 ( 
.A(n_12118),
.B(n_9435),
.Y(n_12533)
);

AND2x2_ASAP7_75t_L g12534 ( 
.A(n_12211),
.B(n_9437),
.Y(n_12534)
);

OR2x2_ASAP7_75t_L g12535 ( 
.A(n_12072),
.B(n_9437),
.Y(n_12535)
);

NAND2xp5_ASAP7_75t_L g12536 ( 
.A(n_12119),
.B(n_9440),
.Y(n_12536)
);

AND2x4_ASAP7_75t_L g12537 ( 
.A(n_12135),
.B(n_8685),
.Y(n_12537)
);

AND2x2_ASAP7_75t_L g12538 ( 
.A(n_12030),
.B(n_9440),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_12026),
.Y(n_12539)
);

OR2x2_ASAP7_75t_L g12540 ( 
.A(n_12088),
.B(n_9442),
.Y(n_12540)
);

OR2x2_ASAP7_75t_L g12541 ( 
.A(n_11808),
.B(n_9442),
.Y(n_12541)
);

AND2x2_ASAP7_75t_L g12542 ( 
.A(n_12196),
.B(n_9445),
.Y(n_12542)
);

OR2x2_ASAP7_75t_L g12543 ( 
.A(n_11976),
.B(n_9445),
.Y(n_12543)
);

INVx1_ASAP7_75t_L g12544 ( 
.A(n_12099),
.Y(n_12544)
);

INVx1_ASAP7_75t_L g12545 ( 
.A(n_11891),
.Y(n_12545)
);

INVx2_ASAP7_75t_L g12546 ( 
.A(n_12032),
.Y(n_12546)
);

INVx2_ASAP7_75t_L g12547 ( 
.A(n_12189),
.Y(n_12547)
);

AND2x2_ASAP7_75t_L g12548 ( 
.A(n_11924),
.B(n_9447),
.Y(n_12548)
);

INVx1_ASAP7_75t_L g12549 ( 
.A(n_12108),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_11942),
.B(n_9447),
.Y(n_12550)
);

INVx1_ASAP7_75t_L g12551 ( 
.A(n_11840),
.Y(n_12551)
);

AND2x2_ASAP7_75t_L g12552 ( 
.A(n_11784),
.B(n_9448),
.Y(n_12552)
);

INVx1_ASAP7_75t_L g12553 ( 
.A(n_11846),
.Y(n_12553)
);

INVx1_ASAP7_75t_L g12554 ( 
.A(n_12171),
.Y(n_12554)
);

NAND2xp5_ASAP7_75t_L g12555 ( 
.A(n_12049),
.B(n_9448),
.Y(n_12555)
);

NAND2xp5_ASAP7_75t_L g12556 ( 
.A(n_11898),
.B(n_9451),
.Y(n_12556)
);

INVx2_ASAP7_75t_L g12557 ( 
.A(n_12189),
.Y(n_12557)
);

AND2x4_ASAP7_75t_SL g12558 ( 
.A(n_12205),
.B(n_7410),
.Y(n_12558)
);

INVx1_ASAP7_75t_L g12559 ( 
.A(n_12174),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_11999),
.B(n_9451),
.Y(n_12560)
);

INVx2_ASAP7_75t_L g12561 ( 
.A(n_12215),
.Y(n_12561)
);

NOR2xp33_ASAP7_75t_L g12562 ( 
.A(n_11724),
.B(n_12209),
.Y(n_12562)
);

HB1xp67_ASAP7_75t_L g12563 ( 
.A(n_11801),
.Y(n_12563)
);

INVx1_ASAP7_75t_L g12564 ( 
.A(n_12177),
.Y(n_12564)
);

AND2x2_ASAP7_75t_L g12565 ( 
.A(n_11787),
.B(n_9456),
.Y(n_12565)
);

OR2x2_ASAP7_75t_L g12566 ( 
.A(n_11996),
.B(n_9456),
.Y(n_12566)
);

BUFx2_ASAP7_75t_L g12567 ( 
.A(n_12207),
.Y(n_12567)
);

INVx1_ASAP7_75t_L g12568 ( 
.A(n_12197),
.Y(n_12568)
);

NAND2xp5_ASAP7_75t_L g12569 ( 
.A(n_12003),
.B(n_9458),
.Y(n_12569)
);

INVx1_ASAP7_75t_L g12570 ( 
.A(n_12220),
.Y(n_12570)
);

AND2x2_ASAP7_75t_L g12571 ( 
.A(n_12010),
.B(n_9458),
.Y(n_12571)
);

INVx1_ASAP7_75t_L g12572 ( 
.A(n_12084),
.Y(n_12572)
);

AND2x4_ASAP7_75t_L g12573 ( 
.A(n_11742),
.B(n_8685),
.Y(n_12573)
);

INVx2_ASAP7_75t_L g12574 ( 
.A(n_12215),
.Y(n_12574)
);

NAND2xp5_ASAP7_75t_L g12575 ( 
.A(n_12009),
.B(n_12059),
.Y(n_12575)
);

INVx2_ASAP7_75t_L g12576 ( 
.A(n_12154),
.Y(n_12576)
);

AND2x2_ASAP7_75t_L g12577 ( 
.A(n_12224),
.B(n_9475),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_12153),
.Y(n_12578)
);

AND2x2_ASAP7_75t_L g12579 ( 
.A(n_12236),
.B(n_9475),
.Y(n_12579)
);

NAND2xp5_ASAP7_75t_L g12580 ( 
.A(n_11821),
.B(n_9479),
.Y(n_12580)
);

INVx1_ASAP7_75t_L g12581 ( 
.A(n_12167),
.Y(n_12581)
);

AND2x2_ASAP7_75t_L g12582 ( 
.A(n_12156),
.B(n_9479),
.Y(n_12582)
);

AND2x2_ASAP7_75t_L g12583 ( 
.A(n_12232),
.B(n_11897),
.Y(n_12583)
);

HB1xp67_ASAP7_75t_L g12584 ( 
.A(n_11951),
.Y(n_12584)
);

INVx1_ASAP7_75t_L g12585 ( 
.A(n_12182),
.Y(n_12585)
);

AND2x4_ASAP7_75t_L g12586 ( 
.A(n_12208),
.B(n_8685),
.Y(n_12586)
);

OR2x6_ASAP7_75t_L g12587 ( 
.A(n_11752),
.B(n_6939),
.Y(n_12587)
);

AND2x4_ASAP7_75t_L g12588 ( 
.A(n_12208),
.B(n_8685),
.Y(n_12588)
);

AND2x2_ASAP7_75t_L g12589 ( 
.A(n_11965),
.B(n_9482),
.Y(n_12589)
);

AND2x2_ASAP7_75t_L g12590 ( 
.A(n_12192),
.B(n_9482),
.Y(n_12590)
);

INVx1_ASAP7_75t_L g12591 ( 
.A(n_12186),
.Y(n_12591)
);

INVx2_ASAP7_75t_L g12592 ( 
.A(n_12154),
.Y(n_12592)
);

HB1xp67_ASAP7_75t_L g12593 ( 
.A(n_11887),
.Y(n_12593)
);

INVx1_ASAP7_75t_L g12594 ( 
.A(n_12195),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_12200),
.Y(n_12595)
);

AND2x2_ASAP7_75t_L g12596 ( 
.A(n_12137),
.B(n_9483),
.Y(n_12596)
);

INVx2_ASAP7_75t_L g12597 ( 
.A(n_12200),
.Y(n_12597)
);

OR2x2_ASAP7_75t_L g12598 ( 
.A(n_12187),
.B(n_9483),
.Y(n_12598)
);

AND2x2_ASAP7_75t_L g12599 ( 
.A(n_12143),
.B(n_9484),
.Y(n_12599)
);

AND2x2_ASAP7_75t_L g12600 ( 
.A(n_12169),
.B(n_9484),
.Y(n_12600)
);

OAI22xp5_ASAP7_75t_L g12601 ( 
.A1(n_11994),
.A2(n_8721),
.B1(n_8540),
.B2(n_7820),
.Y(n_12601)
);

OR2x2_ASAP7_75t_L g12602 ( 
.A(n_11878),
.B(n_9488),
.Y(n_12602)
);

AND2x2_ASAP7_75t_L g12603 ( 
.A(n_11761),
.B(n_9488),
.Y(n_12603)
);

HB1xp67_ASAP7_75t_L g12604 ( 
.A(n_11887),
.Y(n_12604)
);

INVx1_ASAP7_75t_L g12605 ( 
.A(n_12198),
.Y(n_12605)
);

INVx2_ASAP7_75t_L g12606 ( 
.A(n_12040),
.Y(n_12606)
);

AND2x2_ASAP7_75t_L g12607 ( 
.A(n_11852),
.B(n_9489),
.Y(n_12607)
);

NOR2xp67_ASAP7_75t_L g12608 ( 
.A(n_11858),
.B(n_8256),
.Y(n_12608)
);

INVx2_ASAP7_75t_L g12609 ( 
.A(n_12040),
.Y(n_12609)
);

AND2x2_ASAP7_75t_L g12610 ( 
.A(n_12115),
.B(n_12053),
.Y(n_12610)
);

INVx1_ASAP7_75t_L g12611 ( 
.A(n_12210),
.Y(n_12611)
);

OR2x2_ASAP7_75t_L g12612 ( 
.A(n_11979),
.B(n_9489),
.Y(n_12612)
);

AND2x2_ASAP7_75t_L g12613 ( 
.A(n_11791),
.B(n_9494),
.Y(n_12613)
);

NAND2xp5_ASAP7_75t_L g12614 ( 
.A(n_12223),
.B(n_9494),
.Y(n_12614)
);

INVx1_ASAP7_75t_L g12615 ( 
.A(n_12223),
.Y(n_12615)
);

INVx2_ASAP7_75t_SL g12616 ( 
.A(n_12160),
.Y(n_12616)
);

INVx2_ASAP7_75t_L g12617 ( 
.A(n_12124),
.Y(n_12617)
);

OR2x2_ASAP7_75t_L g12618 ( 
.A(n_11768),
.B(n_9497),
.Y(n_12618)
);

NAND2xp5_ASAP7_75t_L g12619 ( 
.A(n_12190),
.B(n_9497),
.Y(n_12619)
);

NAND2xp5_ASAP7_75t_L g12620 ( 
.A(n_11923),
.B(n_9505),
.Y(n_12620)
);

INVx1_ASAP7_75t_L g12621 ( 
.A(n_12090),
.Y(n_12621)
);

INVx2_ASAP7_75t_L g12622 ( 
.A(n_12124),
.Y(n_12622)
);

INVx2_ASAP7_75t_L g12623 ( 
.A(n_12071),
.Y(n_12623)
);

AND2x2_ASAP7_75t_L g12624 ( 
.A(n_11800),
.B(n_9505),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12046),
.Y(n_12625)
);

INVx2_ASAP7_75t_L g12626 ( 
.A(n_12086),
.Y(n_12626)
);

INVx1_ASAP7_75t_L g12627 ( 
.A(n_12046),
.Y(n_12627)
);

NOR2xp33_ASAP7_75t_L g12628 ( 
.A(n_11853),
.B(n_7513),
.Y(n_12628)
);

INVx1_ASAP7_75t_L g12629 ( 
.A(n_12054),
.Y(n_12629)
);

NAND2xp5_ASAP7_75t_L g12630 ( 
.A(n_12130),
.B(n_9508),
.Y(n_12630)
);

AND2x2_ASAP7_75t_L g12631 ( 
.A(n_12120),
.B(n_9508),
.Y(n_12631)
);

NOR2x1_ASAP7_75t_L g12632 ( 
.A(n_11892),
.B(n_9912),
.Y(n_12632)
);

INVx1_ASAP7_75t_L g12633 ( 
.A(n_12054),
.Y(n_12633)
);

INVx2_ASAP7_75t_L g12634 ( 
.A(n_12160),
.Y(n_12634)
);

INVx2_ASAP7_75t_L g12635 ( 
.A(n_12080),
.Y(n_12635)
);

AND2x2_ASAP7_75t_L g12636 ( 
.A(n_11766),
.B(n_9514),
.Y(n_12636)
);

AND2x2_ASAP7_75t_L g12637 ( 
.A(n_11767),
.B(n_9514),
.Y(n_12637)
);

HB1xp67_ASAP7_75t_L g12638 ( 
.A(n_11887),
.Y(n_12638)
);

NOR2x1p5_ASAP7_75t_L g12639 ( 
.A(n_12081),
.B(n_7410),
.Y(n_12639)
);

INVx1_ASAP7_75t_L g12640 ( 
.A(n_12126),
.Y(n_12640)
);

NAND3xp33_ASAP7_75t_L g12641 ( 
.A(n_11772),
.B(n_8726),
.C(n_8685),
.Y(n_12641)
);

AND2x4_ASAP7_75t_L g12642 ( 
.A(n_11892),
.B(n_8685),
.Y(n_12642)
);

INVx2_ASAP7_75t_L g12643 ( 
.A(n_12112),
.Y(n_12643)
);

OR2x2_ASAP7_75t_L g12644 ( 
.A(n_11798),
.B(n_9515),
.Y(n_12644)
);

AND2x2_ASAP7_75t_L g12645 ( 
.A(n_11774),
.B(n_9515),
.Y(n_12645)
);

NAND2xp5_ASAP7_75t_SL g12646 ( 
.A(n_12235),
.B(n_12229),
.Y(n_12646)
);

AND2x4_ASAP7_75t_L g12647 ( 
.A(n_11936),
.B(n_8685),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_12151),
.Y(n_12648)
);

OR2x2_ASAP7_75t_L g12649 ( 
.A(n_11804),
.B(n_9521),
.Y(n_12649)
);

AND2x2_ASAP7_75t_L g12650 ( 
.A(n_12163),
.B(n_9521),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_12152),
.Y(n_12651)
);

INVx2_ASAP7_75t_L g12652 ( 
.A(n_12114),
.Y(n_12652)
);

INVx1_ASAP7_75t_L g12653 ( 
.A(n_12157),
.Y(n_12653)
);

NAND2xp5_ASAP7_75t_L g12654 ( 
.A(n_11769),
.B(n_9522),
.Y(n_12654)
);

INVx1_ASAP7_75t_L g12655 ( 
.A(n_12121),
.Y(n_12655)
);

NOR2xp33_ASAP7_75t_L g12656 ( 
.A(n_12004),
.B(n_7628),
.Y(n_12656)
);

AND2x2_ASAP7_75t_L g12657 ( 
.A(n_12109),
.B(n_9522),
.Y(n_12657)
);

INVx1_ASAP7_75t_L g12658 ( 
.A(n_12216),
.Y(n_12658)
);

AND2x4_ASAP7_75t_SL g12659 ( 
.A(n_11960),
.B(n_7474),
.Y(n_12659)
);

INVx1_ASAP7_75t_L g12660 ( 
.A(n_12218),
.Y(n_12660)
);

INVx1_ASAP7_75t_L g12661 ( 
.A(n_12218),
.Y(n_12661)
);

INVxp67_ASAP7_75t_L g12662 ( 
.A(n_12228),
.Y(n_12662)
);

INVx1_ASAP7_75t_L g12663 ( 
.A(n_11936),
.Y(n_12663)
);

AND2x4_ASAP7_75t_SL g12664 ( 
.A(n_11989),
.B(n_7474),
.Y(n_12664)
);

INVxp67_ASAP7_75t_L g12665 ( 
.A(n_12231),
.Y(n_12665)
);

AND2x2_ASAP7_75t_L g12666 ( 
.A(n_12146),
.B(n_9532),
.Y(n_12666)
);

AND2x2_ASAP7_75t_L g12667 ( 
.A(n_11997),
.B(n_9532),
.Y(n_12667)
);

INVx1_ASAP7_75t_L g12668 ( 
.A(n_11948),
.Y(n_12668)
);

NAND2xp5_ASAP7_75t_L g12669 ( 
.A(n_11948),
.B(n_9538),
.Y(n_12669)
);

INVx1_ASAP7_75t_L g12670 ( 
.A(n_11952),
.Y(n_12670)
);

NOR2xp33_ASAP7_75t_L g12671 ( 
.A(n_11812),
.B(n_7758),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_11952),
.Y(n_12672)
);

INVx2_ASAP7_75t_SL g12673 ( 
.A(n_12212),
.Y(n_12673)
);

OR2x2_ASAP7_75t_L g12674 ( 
.A(n_12240),
.B(n_9538),
.Y(n_12674)
);

INVx2_ASAP7_75t_SL g12675 ( 
.A(n_12217),
.Y(n_12675)
);

NAND2xp5_ASAP7_75t_L g12676 ( 
.A(n_12074),
.B(n_9542),
.Y(n_12676)
);

HB1xp67_ASAP7_75t_L g12677 ( 
.A(n_12199),
.Y(n_12677)
);

INVx2_ASAP7_75t_L g12678 ( 
.A(n_12096),
.Y(n_12678)
);

NAND2xp5_ASAP7_75t_L g12679 ( 
.A(n_12078),
.B(n_9542),
.Y(n_12679)
);

INVx1_ASAP7_75t_L g12680 ( 
.A(n_12098),
.Y(n_12680)
);

NOR2xp33_ASAP7_75t_L g12681 ( 
.A(n_11870),
.B(n_6939),
.Y(n_12681)
);

BUFx3_ASAP7_75t_L g12682 ( 
.A(n_12131),
.Y(n_12682)
);

INVx1_ASAP7_75t_L g12683 ( 
.A(n_12129),
.Y(n_12683)
);

INVx1_ASAP7_75t_L g12684 ( 
.A(n_12110),
.Y(n_12684)
);

AND2x2_ASAP7_75t_L g12685 ( 
.A(n_12134),
.B(n_9549),
.Y(n_12685)
);

AND2x2_ASAP7_75t_L g12686 ( 
.A(n_12206),
.B(n_9549),
.Y(n_12686)
);

BUFx2_ASAP7_75t_L g12687 ( 
.A(n_12077),
.Y(n_12687)
);

INVx1_ASAP7_75t_L g12688 ( 
.A(n_12116),
.Y(n_12688)
);

OR2x2_ASAP7_75t_L g12689 ( 
.A(n_11912),
.B(n_9551),
.Y(n_12689)
);

NAND2xp5_ASAP7_75t_L g12690 ( 
.A(n_12091),
.B(n_9551),
.Y(n_12690)
);

INVx1_ASAP7_75t_L g12691 ( 
.A(n_11971),
.Y(n_12691)
);

NAND2xp5_ASAP7_75t_L g12692 ( 
.A(n_12092),
.B(n_9555),
.Y(n_12692)
);

INVx1_ASAP7_75t_L g12693 ( 
.A(n_11978),
.Y(n_12693)
);

OR2x2_ASAP7_75t_L g12694 ( 
.A(n_12011),
.B(n_9555),
.Y(n_12694)
);

OR2x2_ASAP7_75t_L g12695 ( 
.A(n_11880),
.B(n_9556),
.Y(n_12695)
);

BUFx2_ASAP7_75t_L g12696 ( 
.A(n_11955),
.Y(n_12696)
);

INVx1_ASAP7_75t_L g12697 ( 
.A(n_12005),
.Y(n_12697)
);

AND2x2_ASAP7_75t_L g12698 ( 
.A(n_12147),
.B(n_9556),
.Y(n_12698)
);

AND2x4_ASAP7_75t_L g12699 ( 
.A(n_11927),
.B(n_8726),
.Y(n_12699)
);

INVx1_ASAP7_75t_L g12700 ( 
.A(n_12016),
.Y(n_12700)
);

BUFx2_ASAP7_75t_L g12701 ( 
.A(n_11968),
.Y(n_12701)
);

AND2x2_ASAP7_75t_L g12702 ( 
.A(n_12066),
.B(n_9558),
.Y(n_12702)
);

NAND2xp5_ASAP7_75t_L g12703 ( 
.A(n_12093),
.B(n_9558),
.Y(n_12703)
);

INVx1_ASAP7_75t_L g12704 ( 
.A(n_11988),
.Y(n_12704)
);

AND2x2_ASAP7_75t_L g12705 ( 
.A(n_12070),
.B(n_9560),
.Y(n_12705)
);

OR2x2_ASAP7_75t_L g12706 ( 
.A(n_12101),
.B(n_9560),
.Y(n_12706)
);

INVx1_ASAP7_75t_L g12707 ( 
.A(n_11947),
.Y(n_12707)
);

INVx1_ASAP7_75t_L g12708 ( 
.A(n_12057),
.Y(n_12708)
);

NAND2xp5_ASAP7_75t_L g12709 ( 
.A(n_12102),
.B(n_12106),
.Y(n_12709)
);

AND2x4_ASAP7_75t_L g12710 ( 
.A(n_11805),
.B(n_8726),
.Y(n_12710)
);

NOR2x1_ASAP7_75t_L g12711 ( 
.A(n_11981),
.B(n_10045),
.Y(n_12711)
);

NAND2xp5_ASAP7_75t_L g12712 ( 
.A(n_12122),
.B(n_9568),
.Y(n_12712)
);

OR2x2_ASAP7_75t_L g12713 ( 
.A(n_12007),
.B(n_9568),
.Y(n_12713)
);

AND2x2_ASAP7_75t_L g12714 ( 
.A(n_12085),
.B(n_9572),
.Y(n_12714)
);

INVx1_ASAP7_75t_L g12715 ( 
.A(n_12367),
.Y(n_12715)
);

INVx1_ASAP7_75t_L g12716 ( 
.A(n_12394),
.Y(n_12716)
);

INVx1_ASAP7_75t_L g12717 ( 
.A(n_12463),
.Y(n_12717)
);

INVx1_ASAP7_75t_L g12718 ( 
.A(n_12299),
.Y(n_12718)
);

OAI33xp33_ASAP7_75t_L g12719 ( 
.A1(n_12497),
.A2(n_12214),
.A3(n_12201),
.B1(n_12213),
.B2(n_12194),
.B3(n_11835),
.Y(n_12719)
);

INVx1_ASAP7_75t_L g12720 ( 
.A(n_12593),
.Y(n_12720)
);

INVxp67_ASAP7_75t_SL g12721 ( 
.A(n_12249),
.Y(n_12721)
);

INVx2_ASAP7_75t_L g12722 ( 
.A(n_12255),
.Y(n_12722)
);

NAND2xp5_ASAP7_75t_L g12723 ( 
.A(n_12346),
.B(n_12329),
.Y(n_12723)
);

INVx1_ASAP7_75t_L g12724 ( 
.A(n_12604),
.Y(n_12724)
);

AND2x2_ASAP7_75t_L g12725 ( 
.A(n_12241),
.B(n_11855),
.Y(n_12725)
);

NAND2xp5_ASAP7_75t_L g12726 ( 
.A(n_12346),
.B(n_11856),
.Y(n_12726)
);

NAND2xp5_ASAP7_75t_L g12727 ( 
.A(n_12293),
.B(n_11862),
.Y(n_12727)
);

INVx1_ASAP7_75t_L g12728 ( 
.A(n_12638),
.Y(n_12728)
);

AND2x2_ASAP7_75t_L g12729 ( 
.A(n_12242),
.B(n_11874),
.Y(n_12729)
);

OAI21xp33_ASAP7_75t_L g12730 ( 
.A1(n_12562),
.A2(n_12379),
.B(n_12283),
.Y(n_12730)
);

NAND2xp5_ASAP7_75t_L g12731 ( 
.A(n_12311),
.B(n_11903),
.Y(n_12731)
);

INVx1_ASAP7_75t_L g12732 ( 
.A(n_12321),
.Y(n_12732)
);

INVx1_ASAP7_75t_L g12733 ( 
.A(n_12324),
.Y(n_12733)
);

AND2x2_ASAP7_75t_L g12734 ( 
.A(n_12257),
.B(n_12172),
.Y(n_12734)
);

INVx1_ASAP7_75t_L g12735 ( 
.A(n_12372),
.Y(n_12735)
);

OR2x2_ASAP7_75t_L g12736 ( 
.A(n_12561),
.B(n_12179),
.Y(n_12736)
);

INVx2_ASAP7_75t_L g12737 ( 
.A(n_12259),
.Y(n_12737)
);

NAND2x1_ASAP7_75t_L g12738 ( 
.A(n_12330),
.B(n_12235),
.Y(n_12738)
);

AND2x4_ASAP7_75t_L g12739 ( 
.A(n_12330),
.B(n_11811),
.Y(n_12739)
);

OAI211xp5_ASAP7_75t_SL g12740 ( 
.A1(n_12432),
.A2(n_12148),
.B(n_11987),
.C(n_12138),
.Y(n_12740)
);

INVx1_ASAP7_75t_L g12741 ( 
.A(n_12383),
.Y(n_12741)
);

OR2x2_ASAP7_75t_L g12742 ( 
.A(n_12574),
.B(n_11905),
.Y(n_12742)
);

NAND2xp5_ASAP7_75t_L g12743 ( 
.A(n_12309),
.B(n_11907),
.Y(n_12743)
);

OR2x2_ASAP7_75t_L g12744 ( 
.A(n_12289),
.B(n_11910),
.Y(n_12744)
);

INVx1_ASAP7_75t_L g12745 ( 
.A(n_12263),
.Y(n_12745)
);

INVx3_ASAP7_75t_R g12746 ( 
.A(n_12250),
.Y(n_12746)
);

OR2x2_ASAP7_75t_L g12747 ( 
.A(n_12419),
.B(n_12425),
.Y(n_12747)
);

OR2x2_ASAP7_75t_L g12748 ( 
.A(n_12466),
.B(n_12165),
.Y(n_12748)
);

INVx1_ASAP7_75t_L g12749 ( 
.A(n_12248),
.Y(n_12749)
);

AOI221xp5_ASAP7_75t_L g12750 ( 
.A1(n_12422),
.A2(n_12696),
.B1(n_12437),
.B2(n_12707),
.C(n_12355),
.Y(n_12750)
);

INVx1_ASAP7_75t_L g12751 ( 
.A(n_12248),
.Y(n_12751)
);

NAND2xp5_ASAP7_75t_L g12752 ( 
.A(n_12502),
.B(n_12214),
.Y(n_12752)
);

AND2x2_ASAP7_75t_L g12753 ( 
.A(n_12364),
.B(n_12166),
.Y(n_12753)
);

OR2x2_ASAP7_75t_L g12754 ( 
.A(n_12253),
.B(n_12139),
.Y(n_12754)
);

NAND2xp5_ASAP7_75t_L g12755 ( 
.A(n_12323),
.B(n_12194),
.Y(n_12755)
);

AND2x6_ASAP7_75t_SL g12756 ( 
.A(n_12397),
.B(n_11816),
.Y(n_12756)
);

NAND2xp5_ASAP7_75t_L g12757 ( 
.A(n_12427),
.B(n_12201),
.Y(n_12757)
);

AND2x2_ASAP7_75t_L g12758 ( 
.A(n_12243),
.B(n_12278),
.Y(n_12758)
);

NAND2xp5_ASAP7_75t_L g12759 ( 
.A(n_12254),
.B(n_12213),
.Y(n_12759)
);

INVx2_ASAP7_75t_L g12760 ( 
.A(n_12387),
.Y(n_12760)
);

INVx1_ASAP7_75t_L g12761 ( 
.A(n_12687),
.Y(n_12761)
);

OR2x2_ASAP7_75t_L g12762 ( 
.A(n_12262),
.B(n_12498),
.Y(n_12762)
);

NAND2xp5_ASAP7_75t_L g12763 ( 
.A(n_12610),
.B(n_12024),
.Y(n_12763)
);

NAND4xp25_ASAP7_75t_L g12764 ( 
.A(n_12671),
.B(n_12141),
.C(n_11869),
.D(n_12063),
.Y(n_12764)
);

INVx1_ASAP7_75t_L g12765 ( 
.A(n_12677),
.Y(n_12765)
);

INVx1_ASAP7_75t_L g12766 ( 
.A(n_12291),
.Y(n_12766)
);

OR2x2_ASAP7_75t_L g12767 ( 
.A(n_12401),
.B(n_12162),
.Y(n_12767)
);

INVx1_ASAP7_75t_L g12768 ( 
.A(n_12296),
.Y(n_12768)
);

INVx1_ASAP7_75t_L g12769 ( 
.A(n_12307),
.Y(n_12769)
);

OR2x2_ASAP7_75t_L g12770 ( 
.A(n_12361),
.B(n_12028),
.Y(n_12770)
);

AND2x2_ASAP7_75t_L g12771 ( 
.A(n_12659),
.B(n_12039),
.Y(n_12771)
);

INVx3_ASAP7_75t_L g12772 ( 
.A(n_12387),
.Y(n_12772)
);

INVx1_ASAP7_75t_L g12773 ( 
.A(n_12308),
.Y(n_12773)
);

AND2x2_ASAP7_75t_L g12774 ( 
.A(n_12244),
.B(n_12044),
.Y(n_12774)
);

INVx1_ASAP7_75t_L g12775 ( 
.A(n_12310),
.Y(n_12775)
);

AND2x2_ASAP7_75t_SL g12776 ( 
.A(n_12371),
.B(n_12393),
.Y(n_12776)
);

OR2x2_ASAP7_75t_L g12777 ( 
.A(n_12315),
.B(n_12061),
.Y(n_12777)
);

NAND2xp5_ASAP7_75t_L g12778 ( 
.A(n_12276),
.B(n_12073),
.Y(n_12778)
);

AND2x2_ASAP7_75t_L g12779 ( 
.A(n_12305),
.B(n_11830),
.Y(n_12779)
);

INVx1_ASAP7_75t_L g12780 ( 
.A(n_12313),
.Y(n_12780)
);

OR2x2_ASAP7_75t_L g12781 ( 
.A(n_12354),
.B(n_11836),
.Y(n_12781)
);

INVx2_ASAP7_75t_SL g12782 ( 
.A(n_12431),
.Y(n_12782)
);

INVxp67_ASAP7_75t_SL g12783 ( 
.A(n_12359),
.Y(n_12783)
);

INVx1_ASAP7_75t_SL g12784 ( 
.A(n_12348),
.Y(n_12784)
);

NAND2xp5_ASAP7_75t_L g12785 ( 
.A(n_12290),
.B(n_11841),
.Y(n_12785)
);

OR2x2_ASAP7_75t_L g12786 ( 
.A(n_12464),
.B(n_12036),
.Y(n_12786)
);

NAND2xp5_ASAP7_75t_L g12787 ( 
.A(n_12424),
.B(n_12336),
.Y(n_12787)
);

AOI22xp33_ASAP7_75t_L g12788 ( 
.A1(n_12707),
.A2(n_12181),
.B1(n_12008),
.B2(n_12140),
.Y(n_12788)
);

OR2x2_ASAP7_75t_L g12789 ( 
.A(n_12465),
.B(n_12056),
.Y(n_12789)
);

AND2x4_ASAP7_75t_L g12790 ( 
.A(n_12264),
.B(n_12222),
.Y(n_12790)
);

AND2x2_ASAP7_75t_L g12791 ( 
.A(n_12261),
.B(n_12233),
.Y(n_12791)
);

INVx2_ASAP7_75t_L g12792 ( 
.A(n_12431),
.Y(n_12792)
);

AND2x2_ASAP7_75t_L g12793 ( 
.A(n_12337),
.B(n_12164),
.Y(n_12793)
);

INVx1_ASAP7_75t_L g12794 ( 
.A(n_12563),
.Y(n_12794)
);

OR2x2_ASAP7_75t_L g12795 ( 
.A(n_12351),
.B(n_12132),
.Y(n_12795)
);

NOR2x1_ASAP7_75t_L g12796 ( 
.A(n_12362),
.B(n_12176),
.Y(n_12796)
);

NAND2xp5_ASAP7_75t_L g12797 ( 
.A(n_12344),
.B(n_12014),
.Y(n_12797)
);

NAND2xp5_ASAP7_75t_L g12798 ( 
.A(n_12281),
.B(n_12339),
.Y(n_12798)
);

HB1xp67_ASAP7_75t_L g12799 ( 
.A(n_12433),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12245),
.Y(n_12800)
);

INVx1_ASAP7_75t_L g12801 ( 
.A(n_12433),
.Y(n_12801)
);

OR2x2_ASAP7_75t_L g12802 ( 
.A(n_12317),
.B(n_12297),
.Y(n_12802)
);

NAND2xp5_ASAP7_75t_L g12803 ( 
.A(n_12368),
.B(n_12230),
.Y(n_12803)
);

OAI21xp33_ASAP7_75t_L g12804 ( 
.A1(n_12525),
.A2(n_12238),
.B(n_12226),
.Y(n_12804)
);

AND2x2_ASAP7_75t_L g12805 ( 
.A(n_12567),
.B(n_12100),
.Y(n_12805)
);

INVx2_ASAP7_75t_L g12806 ( 
.A(n_12328),
.Y(n_12806)
);

OAI22xp33_ASAP7_75t_L g12807 ( 
.A1(n_12353),
.A2(n_12075),
.B1(n_11967),
.B2(n_12142),
.Y(n_12807)
);

NAND2xp5_ASAP7_75t_L g12808 ( 
.A(n_12449),
.B(n_12155),
.Y(n_12808)
);

AND2x4_ASAP7_75t_L g12809 ( 
.A(n_12616),
.B(n_12128),
.Y(n_12809)
);

OR2x2_ASAP7_75t_L g12810 ( 
.A(n_12268),
.B(n_12376),
.Y(n_12810)
);

HB1xp67_ASAP7_75t_L g12811 ( 
.A(n_12356),
.Y(n_12811)
);

NOR2xp33_ASAP7_75t_L g12812 ( 
.A(n_12451),
.B(n_11882),
.Y(n_12812)
);

OR2x2_ASAP7_75t_L g12813 ( 
.A(n_12395),
.B(n_12062),
.Y(n_12813)
);

AND2x2_ASAP7_75t_L g12814 ( 
.A(n_12441),
.B(n_12103),
.Y(n_12814)
);

INVxp67_ASAP7_75t_L g12815 ( 
.A(n_12584),
.Y(n_12815)
);

INVx1_ASAP7_75t_L g12816 ( 
.A(n_12320),
.Y(n_12816)
);

NAND2xp5_ASAP7_75t_L g12817 ( 
.A(n_12449),
.B(n_12133),
.Y(n_12817)
);

INVx2_ASAP7_75t_L g12818 ( 
.A(n_12384),
.Y(n_12818)
);

OR2x2_ASAP7_75t_L g12819 ( 
.A(n_12270),
.B(n_11944),
.Y(n_12819)
);

AND2x2_ASAP7_75t_L g12820 ( 
.A(n_12246),
.B(n_12104),
.Y(n_12820)
);

INVx1_ASAP7_75t_L g12821 ( 
.A(n_12446),
.Y(n_12821)
);

INVx1_ASAP7_75t_L g12822 ( 
.A(n_12490),
.Y(n_12822)
);

AND2x2_ASAP7_75t_L g12823 ( 
.A(n_12524),
.B(n_12144),
.Y(n_12823)
);

INVx1_ASAP7_75t_L g12824 ( 
.A(n_12408),
.Y(n_12824)
);

AND2x2_ASAP7_75t_L g12825 ( 
.A(n_12504),
.B(n_12158),
.Y(n_12825)
);

INVx2_ASAP7_75t_L g12826 ( 
.A(n_12418),
.Y(n_12826)
);

NAND2x1_ASAP7_75t_SL g12827 ( 
.A(n_12332),
.B(n_12145),
.Y(n_12827)
);

NAND2xp5_ASAP7_75t_L g12828 ( 
.A(n_12583),
.B(n_12161),
.Y(n_12828)
);

AND2x2_ASAP7_75t_L g12829 ( 
.A(n_12300),
.B(n_12173),
.Y(n_12829)
);

AND2x2_ASAP7_75t_L g12830 ( 
.A(n_12295),
.B(n_12178),
.Y(n_12830)
);

OR2x6_ASAP7_75t_L g12831 ( 
.A(n_12491),
.B(n_6939),
.Y(n_12831)
);

NAND2xp5_ASAP7_75t_L g12832 ( 
.A(n_12251),
.B(n_12183),
.Y(n_12832)
);

INVxp67_ASAP7_75t_SL g12833 ( 
.A(n_12711),
.Y(n_12833)
);

AND2x4_ASAP7_75t_L g12834 ( 
.A(n_12493),
.B(n_12184),
.Y(n_12834)
);

NAND2xp5_ASAP7_75t_L g12835 ( 
.A(n_12251),
.B(n_12204),
.Y(n_12835)
);

AND2x2_ASAP7_75t_L g12836 ( 
.A(n_12256),
.B(n_12247),
.Y(n_12836)
);

INVx2_ASAP7_75t_L g12837 ( 
.A(n_12512),
.Y(n_12837)
);

NAND2xp5_ASAP7_75t_L g12838 ( 
.A(n_12365),
.B(n_12180),
.Y(n_12838)
);

BUFx2_ASAP7_75t_L g12839 ( 
.A(n_12348),
.Y(n_12839)
);

INVx2_ASAP7_75t_L g12840 ( 
.A(n_12374),
.Y(n_12840)
);

INVx2_ASAP7_75t_L g12841 ( 
.A(n_12374),
.Y(n_12841)
);

INVx1_ASAP7_75t_L g12842 ( 
.A(n_12708),
.Y(n_12842)
);

NAND2xp5_ASAP7_75t_L g12843 ( 
.A(n_12365),
.B(n_12175),
.Y(n_12843)
);

INVx1_ASAP7_75t_L g12844 ( 
.A(n_12708),
.Y(n_12844)
);

INVx2_ASAP7_75t_L g12845 ( 
.A(n_12326),
.Y(n_12845)
);

NAND2xp5_ASAP7_75t_L g12846 ( 
.A(n_12550),
.B(n_12225),
.Y(n_12846)
);

OAI22xp5_ASAP7_75t_L g12847 ( 
.A1(n_12575),
.A2(n_12149),
.B1(n_12168),
.B2(n_8730),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_12589),
.Y(n_12848)
);

AND2x4_ASAP7_75t_L g12849 ( 
.A(n_12282),
.B(n_12057),
.Y(n_12849)
);

AND2x2_ASAP7_75t_L g12850 ( 
.A(n_12252),
.B(n_12057),
.Y(n_12850)
);

AND2x2_ASAP7_75t_L g12851 ( 
.A(n_12292),
.B(n_9572),
.Y(n_12851)
);

AND2x4_ASAP7_75t_L g12852 ( 
.A(n_12294),
.B(n_7210),
.Y(n_12852)
);

OR2x2_ASAP7_75t_L g12853 ( 
.A(n_12442),
.B(n_9576),
.Y(n_12853)
);

OR2x2_ASAP7_75t_L g12854 ( 
.A(n_12452),
.B(n_9576),
.Y(n_12854)
);

INVxp67_ASAP7_75t_L g12855 ( 
.A(n_12681),
.Y(n_12855)
);

AND2x2_ASAP7_75t_L g12856 ( 
.A(n_12266),
.B(n_9577),
.Y(n_12856)
);

OR2x2_ASAP7_75t_L g12857 ( 
.A(n_12505),
.B(n_9577),
.Y(n_12857)
);

NOR2x1p5_ASAP7_75t_L g12858 ( 
.A(n_12269),
.B(n_11908),
.Y(n_12858)
);

OAI21xp5_ASAP7_75t_L g12859 ( 
.A1(n_12704),
.A2(n_11964),
.B(n_7915),
.Y(n_12859)
);

INVx1_ASAP7_75t_L g12860 ( 
.A(n_12702),
.Y(n_12860)
);

OAI21xp33_ASAP7_75t_L g12861 ( 
.A1(n_12306),
.A2(n_9586),
.B(n_9581),
.Y(n_12861)
);

INVx2_ASAP7_75t_L g12862 ( 
.A(n_12326),
.Y(n_12862)
);

INVx1_ASAP7_75t_L g12863 ( 
.A(n_12705),
.Y(n_12863)
);

INVx1_ASAP7_75t_L g12864 ( 
.A(n_12435),
.Y(n_12864)
);

INVx2_ASAP7_75t_L g12865 ( 
.A(n_12333),
.Y(n_12865)
);

AND2x2_ASAP7_75t_L g12866 ( 
.A(n_12286),
.B(n_9581),
.Y(n_12866)
);

INVx1_ASAP7_75t_L g12867 ( 
.A(n_12488),
.Y(n_12867)
);

NAND3xp33_ASAP7_75t_L g12868 ( 
.A(n_12704),
.B(n_8730),
.C(n_8726),
.Y(n_12868)
);

INVx2_ASAP7_75t_SL g12869 ( 
.A(n_12332),
.Y(n_12869)
);

OR2x2_ASAP7_75t_L g12870 ( 
.A(n_12654),
.B(n_9586),
.Y(n_12870)
);

NAND2x1p5_ASAP7_75t_L g12871 ( 
.A(n_12474),
.B(n_12480),
.Y(n_12871)
);

NOR2x1_ASAP7_75t_L g12872 ( 
.A(n_12632),
.B(n_10045),
.Y(n_12872)
);

INVx2_ASAP7_75t_L g12873 ( 
.A(n_12403),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_12496),
.Y(n_12874)
);

NAND2xp5_ASAP7_75t_L g12875 ( 
.A(n_12322),
.B(n_12331),
.Y(n_12875)
);

NAND2xp5_ASAP7_75t_L g12876 ( 
.A(n_12462),
.B(n_9597),
.Y(n_12876)
);

AND2x2_ASAP7_75t_L g12877 ( 
.A(n_12558),
.B(n_9597),
.Y(n_12877)
);

AND2x2_ASAP7_75t_L g12878 ( 
.A(n_12513),
.B(n_9598),
.Y(n_12878)
);

OR2x2_ASAP7_75t_L g12879 ( 
.A(n_12539),
.B(n_9598),
.Y(n_12879)
);

INVx1_ASAP7_75t_L g12880 ( 
.A(n_12489),
.Y(n_12880)
);

NOR2xp33_ASAP7_75t_L g12881 ( 
.A(n_12404),
.B(n_12407),
.Y(n_12881)
);

AND2x2_ASAP7_75t_L g12882 ( 
.A(n_12546),
.B(n_9606),
.Y(n_12882)
);

NOR3xp33_ASAP7_75t_L g12883 ( 
.A(n_12662),
.B(n_12065),
.C(n_12038),
.Y(n_12883)
);

NAND2xp5_ASAP7_75t_L g12884 ( 
.A(n_12519),
.B(n_9606),
.Y(n_12884)
);

AND2x2_ASAP7_75t_L g12885 ( 
.A(n_12389),
.B(n_9608),
.Y(n_12885)
);

AND2x4_ASAP7_75t_L g12886 ( 
.A(n_12673),
.B(n_7210),
.Y(n_12886)
);

NOR2xp33_ASAP7_75t_L g12887 ( 
.A(n_12386),
.B(n_8726),
.Y(n_12887)
);

OR2x2_ASAP7_75t_L g12888 ( 
.A(n_12416),
.B(n_12423),
.Y(n_12888)
);

HB1xp67_ASAP7_75t_L g12889 ( 
.A(n_12608),
.Y(n_12889)
);

AND2x2_ASAP7_75t_L g12890 ( 
.A(n_12678),
.B(n_9608),
.Y(n_12890)
);

AND2x2_ASAP7_75t_L g12891 ( 
.A(n_12635),
.B(n_9614),
.Y(n_12891)
);

NAND2xp5_ASAP7_75t_L g12892 ( 
.A(n_12520),
.B(n_9614),
.Y(n_12892)
);

INVx2_ASAP7_75t_SL g12893 ( 
.A(n_12586),
.Y(n_12893)
);

AND2x4_ASAP7_75t_L g12894 ( 
.A(n_12576),
.B(n_7820),
.Y(n_12894)
);

OR2x2_ASAP7_75t_L g12895 ( 
.A(n_12340),
.B(n_9616),
.Y(n_12895)
);

AND2x4_ASAP7_75t_L g12896 ( 
.A(n_12675),
.B(n_7210),
.Y(n_12896)
);

INVxp67_ASAP7_75t_L g12897 ( 
.A(n_12507),
.Y(n_12897)
);

AND2x2_ASAP7_75t_L g12898 ( 
.A(n_12643),
.B(n_9616),
.Y(n_12898)
);

INVx1_ASAP7_75t_L g12899 ( 
.A(n_12485),
.Y(n_12899)
);

INVx2_ASAP7_75t_L g12900 ( 
.A(n_12403),
.Y(n_12900)
);

INVxp67_ASAP7_75t_L g12901 ( 
.A(n_12507),
.Y(n_12901)
);

INVx2_ASAP7_75t_L g12902 ( 
.A(n_12411),
.Y(n_12902)
);

AND2x2_ASAP7_75t_L g12903 ( 
.A(n_12652),
.B(n_12447),
.Y(n_12903)
);

AND2x2_ASAP7_75t_L g12904 ( 
.A(n_12400),
.B(n_9623),
.Y(n_12904)
);

INVx1_ASAP7_75t_L g12905 ( 
.A(n_12486),
.Y(n_12905)
);

NOR2xp33_ASAP7_75t_L g12906 ( 
.A(n_12399),
.B(n_8726),
.Y(n_12906)
);

NAND2xp5_ASAP7_75t_L g12907 ( 
.A(n_12398),
.B(n_9623),
.Y(n_12907)
);

NAND4xp25_ASAP7_75t_L g12908 ( 
.A(n_12628),
.B(n_12656),
.C(n_12288),
.D(n_12352),
.Y(n_12908)
);

AND2x4_ASAP7_75t_L g12909 ( 
.A(n_12592),
.B(n_7820),
.Y(n_12909)
);

INVx2_ASAP7_75t_L g12910 ( 
.A(n_12411),
.Y(n_12910)
);

OR2x2_ASAP7_75t_L g12911 ( 
.A(n_12378),
.B(n_9625),
.Y(n_12911)
);

HB1xp67_ASAP7_75t_L g12912 ( 
.A(n_12547),
.Y(n_12912)
);

INVx1_ASAP7_75t_SL g12913 ( 
.A(n_12405),
.Y(n_12913)
);

NAND2xp5_ASAP7_75t_L g12914 ( 
.A(n_12470),
.B(n_9625),
.Y(n_12914)
);

INVx2_ASAP7_75t_L g12915 ( 
.A(n_12434),
.Y(n_12915)
);

INVx1_ASAP7_75t_L g12916 ( 
.A(n_12579),
.Y(n_12916)
);

INVx1_ASAP7_75t_L g12917 ( 
.A(n_12271),
.Y(n_12917)
);

NAND2xp5_ASAP7_75t_L g12918 ( 
.A(n_12595),
.B(n_9634),
.Y(n_12918)
);

OR2x2_ASAP7_75t_L g12919 ( 
.A(n_12258),
.B(n_12327),
.Y(n_12919)
);

AND2x2_ASAP7_75t_L g12920 ( 
.A(n_12590),
.B(n_9634),
.Y(n_12920)
);

INVx1_ASAP7_75t_L g12921 ( 
.A(n_12273),
.Y(n_12921)
);

INVx1_ASAP7_75t_L g12922 ( 
.A(n_12279),
.Y(n_12922)
);

INVx2_ASAP7_75t_L g12923 ( 
.A(n_12434),
.Y(n_12923)
);

AND2x2_ASAP7_75t_L g12924 ( 
.A(n_12319),
.B(n_9636),
.Y(n_12924)
);

INVx1_ASAP7_75t_L g12925 ( 
.A(n_12284),
.Y(n_12925)
);

NAND2xp5_ASAP7_75t_L g12926 ( 
.A(n_12597),
.B(n_12440),
.Y(n_12926)
);

NAND2x1_ASAP7_75t_L g12927 ( 
.A(n_12586),
.B(n_10063),
.Y(n_12927)
);

NAND2xp5_ASAP7_75t_L g12928 ( 
.A(n_12606),
.B(n_9636),
.Y(n_12928)
);

BUFx2_ASAP7_75t_L g12929 ( 
.A(n_12588),
.Y(n_12929)
);

INVx1_ASAP7_75t_SL g12930 ( 
.A(n_12430),
.Y(n_12930)
);

AOI22xp5_ASAP7_75t_L g12931 ( 
.A1(n_12438),
.A2(n_8730),
.B1(n_8726),
.B2(n_7553),
.Y(n_12931)
);

INVx1_ASAP7_75t_L g12932 ( 
.A(n_12285),
.Y(n_12932)
);

NOR2xp33_ASAP7_75t_SL g12933 ( 
.A(n_12499),
.B(n_7278),
.Y(n_12933)
);

AND2x4_ASAP7_75t_L g12934 ( 
.A(n_12634),
.B(n_7829),
.Y(n_12934)
);

AND2x4_ASAP7_75t_L g12935 ( 
.A(n_12500),
.B(n_7829),
.Y(n_12935)
);

NAND2xp5_ASAP7_75t_L g12936 ( 
.A(n_12609),
.B(n_9647),
.Y(n_12936)
);

HB1xp67_ASAP7_75t_L g12937 ( 
.A(n_12557),
.Y(n_12937)
);

AND2x4_ASAP7_75t_L g12938 ( 
.A(n_12615),
.B(n_8730),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12287),
.Y(n_12939)
);

INVx2_ASAP7_75t_L g12940 ( 
.A(n_12370),
.Y(n_12940)
);

INVx1_ASAP7_75t_L g12941 ( 
.A(n_12571),
.Y(n_12941)
);

NOR2xp33_ASAP7_75t_L g12942 ( 
.A(n_12301),
.B(n_8730),
.Y(n_12942)
);

AND2x4_ASAP7_75t_SL g12943 ( 
.A(n_12375),
.B(n_7474),
.Y(n_12943)
);

OR2x2_ASAP7_75t_L g12944 ( 
.A(n_12363),
.B(n_9647),
.Y(n_12944)
);

INVx1_ASAP7_75t_L g12945 ( 
.A(n_12396),
.Y(n_12945)
);

NOR2xp67_ASAP7_75t_L g12946 ( 
.A(n_12641),
.B(n_8256),
.Y(n_12946)
);

NAND2xp5_ASAP7_75t_L g12947 ( 
.A(n_12617),
.B(n_9649),
.Y(n_12947)
);

INVx1_ASAP7_75t_L g12948 ( 
.A(n_12391),
.Y(n_12948)
);

INVx1_ASAP7_75t_L g12949 ( 
.A(n_12409),
.Y(n_12949)
);

AND2x2_ASAP7_75t_L g12950 ( 
.A(n_12406),
.B(n_9649),
.Y(n_12950)
);

INVx1_ASAP7_75t_L g12951 ( 
.A(n_12413),
.Y(n_12951)
);

INVx1_ASAP7_75t_L g12952 ( 
.A(n_12415),
.Y(n_12952)
);

INVx2_ASAP7_75t_L g12953 ( 
.A(n_12366),
.Y(n_12953)
);

INVx1_ASAP7_75t_L g12954 ( 
.A(n_12548),
.Y(n_12954)
);

NAND2xp5_ASAP7_75t_L g12955 ( 
.A(n_12622),
.B(n_9664),
.Y(n_12955)
);

INVxp67_ASAP7_75t_L g12956 ( 
.A(n_12341),
.Y(n_12956)
);

INVx1_ASAP7_75t_L g12957 ( 
.A(n_12369),
.Y(n_12957)
);

OR2x2_ASAP7_75t_L g12958 ( 
.A(n_12516),
.B(n_9664),
.Y(n_12958)
);

INVx1_ASAP7_75t_L g12959 ( 
.A(n_12501),
.Y(n_12959)
);

AND2x2_ASAP7_75t_L g12960 ( 
.A(n_12542),
.B(n_9666),
.Y(n_12960)
);

NAND2xp5_ASAP7_75t_L g12961 ( 
.A(n_12316),
.B(n_12458),
.Y(n_12961)
);

INVx1_ASAP7_75t_L g12962 ( 
.A(n_12420),
.Y(n_12962)
);

OR2x2_ASAP7_75t_L g12963 ( 
.A(n_12390),
.B(n_9666),
.Y(n_12963)
);

INVx2_ASAP7_75t_L g12964 ( 
.A(n_12350),
.Y(n_12964)
);

AND2x4_ASAP7_75t_L g12965 ( 
.A(n_12527),
.B(n_8730),
.Y(n_12965)
);

NAND2x1p5_ASAP7_75t_L g12966 ( 
.A(n_12682),
.B(n_12588),
.Y(n_12966)
);

OR2x2_ASAP7_75t_L g12967 ( 
.A(n_12265),
.B(n_9686),
.Y(n_12967)
);

INVx1_ASAP7_75t_L g12968 ( 
.A(n_12421),
.Y(n_12968)
);

NOR2x1p5_ASAP7_75t_L g12969 ( 
.A(n_12274),
.B(n_12280),
.Y(n_12969)
);

AND2x4_ASAP7_75t_L g12970 ( 
.A(n_12509),
.B(n_8730),
.Y(n_12970)
);

OR2x2_ASAP7_75t_L g12971 ( 
.A(n_12453),
.B(n_9687),
.Y(n_12971)
);

INVx2_ASAP7_75t_L g12972 ( 
.A(n_12381),
.Y(n_12972)
);

OR2x2_ASAP7_75t_L g12973 ( 
.A(n_12260),
.B(n_9687),
.Y(n_12973)
);

INVx2_ASAP7_75t_L g12974 ( 
.A(n_12381),
.Y(n_12974)
);

AND2x4_ASAP7_75t_L g12975 ( 
.A(n_12514),
.B(n_12318),
.Y(n_12975)
);

INVxp67_ASAP7_75t_SL g12976 ( 
.A(n_12479),
.Y(n_12976)
);

INVx3_ASAP7_75t_L g12977 ( 
.A(n_12528),
.Y(n_12977)
);

INVx1_ASAP7_75t_L g12978 ( 
.A(n_12473),
.Y(n_12978)
);

OR2x2_ASAP7_75t_L g12979 ( 
.A(n_12521),
.B(n_9689),
.Y(n_12979)
);

INVx2_ASAP7_75t_L g12980 ( 
.A(n_12357),
.Y(n_12980)
);

NOR2xp33_ASAP7_75t_L g12981 ( 
.A(n_12646),
.B(n_6939),
.Y(n_12981)
);

INVx4_ASAP7_75t_L g12982 ( 
.A(n_12587),
.Y(n_12982)
);

NOR2x1_ASAP7_75t_L g12983 ( 
.A(n_12701),
.B(n_10063),
.Y(n_12983)
);

INVxp67_ASAP7_75t_L g12984 ( 
.A(n_12303),
.Y(n_12984)
);

INVx1_ASAP7_75t_L g12985 ( 
.A(n_12538),
.Y(n_12985)
);

NAND2x1p5_ASAP7_75t_L g12986 ( 
.A(n_12334),
.B(n_7278),
.Y(n_12986)
);

AND2x4_ASAP7_75t_L g12987 ( 
.A(n_12335),
.B(n_9689),
.Y(n_12987)
);

INVx1_ASAP7_75t_L g12988 ( 
.A(n_12596),
.Y(n_12988)
);

INVxp67_ASAP7_75t_L g12989 ( 
.A(n_12689),
.Y(n_12989)
);

NOR3xp33_ASAP7_75t_L g12990 ( 
.A(n_12343),
.B(n_7345),
.C(n_7341),
.Y(n_12990)
);

O2A1O1Ixp33_ASAP7_75t_SL g12991 ( 
.A1(n_12445),
.A2(n_9694),
.B(n_9691),
.C(n_8263),
.Y(n_12991)
);

INVx2_ASAP7_75t_L g12992 ( 
.A(n_12537),
.Y(n_12992)
);

INVx2_ASAP7_75t_L g12993 ( 
.A(n_12537),
.Y(n_12993)
);

NOR2xp33_ASAP7_75t_L g12994 ( 
.A(n_12468),
.B(n_6974),
.Y(n_12994)
);

NAND2xp5_ASAP7_75t_L g12995 ( 
.A(n_12382),
.B(n_8256),
.Y(n_12995)
);

NAND2xp5_ASAP7_75t_L g12996 ( 
.A(n_12531),
.B(n_8256),
.Y(n_12996)
);

NAND2xp5_ASAP7_75t_L g12997 ( 
.A(n_12338),
.B(n_8263),
.Y(n_12997)
);

INVx1_ASAP7_75t_L g12998 ( 
.A(n_12599),
.Y(n_12998)
);

INVx1_ASAP7_75t_L g12999 ( 
.A(n_12511),
.Y(n_12999)
);

NAND2x1p5_ASAP7_75t_L g13000 ( 
.A(n_12342),
.B(n_12358),
.Y(n_13000)
);

INVx1_ASAP7_75t_L g13001 ( 
.A(n_12402),
.Y(n_13001)
);

INVx1_ASAP7_75t_L g13002 ( 
.A(n_12459),
.Y(n_13002)
);

INVx1_ASAP7_75t_SL g13003 ( 
.A(n_12664),
.Y(n_13003)
);

AND2x4_ASAP7_75t_L g13004 ( 
.A(n_12639),
.B(n_7251),
.Y(n_13004)
);

INVx2_ASAP7_75t_SL g13005 ( 
.A(n_12528),
.Y(n_13005)
);

AND2x2_ASAP7_75t_L g13006 ( 
.A(n_12623),
.B(n_8263),
.Y(n_13006)
);

NOR2xp33_ASAP7_75t_L g13007 ( 
.A(n_12272),
.B(n_6974),
.Y(n_13007)
);

NAND2xp5_ASAP7_75t_L g13008 ( 
.A(n_12360),
.B(n_8263),
.Y(n_13008)
);

INVx1_ASAP7_75t_L g13009 ( 
.A(n_12475),
.Y(n_13009)
);

HB1xp67_ASAP7_75t_SL g13010 ( 
.A(n_12426),
.Y(n_13010)
);

OR2x2_ASAP7_75t_L g13011 ( 
.A(n_12580),
.B(n_9104),
.Y(n_13011)
);

INVx1_ASAP7_75t_SL g13012 ( 
.A(n_12699),
.Y(n_13012)
);

AND2x2_ASAP7_75t_L g13013 ( 
.A(n_12626),
.B(n_8263),
.Y(n_13013)
);

AND2x2_ASAP7_75t_L g13014 ( 
.A(n_12436),
.B(n_8304),
.Y(n_13014)
);

INVx1_ASAP7_75t_L g13015 ( 
.A(n_12476),
.Y(n_13015)
);

AND2x2_ASAP7_75t_L g13016 ( 
.A(n_12503),
.B(n_8304),
.Y(n_13016)
);

INVx2_ASAP7_75t_SL g13017 ( 
.A(n_12573),
.Y(n_13017)
);

INVx1_ASAP7_75t_L g13018 ( 
.A(n_12380),
.Y(n_13018)
);

NAND2xp5_ASAP7_75t_L g13019 ( 
.A(n_12665),
.B(n_8304),
.Y(n_13019)
);

NOR2xp33_ASAP7_75t_L g13020 ( 
.A(n_12275),
.B(n_6974),
.Y(n_13020)
);

OR2x6_ASAP7_75t_L g13021 ( 
.A(n_12578),
.B(n_7024),
.Y(n_13021)
);

INVx1_ASAP7_75t_L g13022 ( 
.A(n_12388),
.Y(n_13022)
);

AND2x2_ASAP7_75t_L g13023 ( 
.A(n_12587),
.B(n_8304),
.Y(n_13023)
);

INVx2_ASAP7_75t_L g13024 ( 
.A(n_12573),
.Y(n_13024)
);

AND2x2_ASAP7_75t_L g13025 ( 
.A(n_12714),
.B(n_8304),
.Y(n_13025)
);

INVx3_ASAP7_75t_L g13026 ( 
.A(n_12710),
.Y(n_13026)
);

OAI33xp33_ASAP7_75t_L g13027 ( 
.A1(n_12630),
.A2(n_12545),
.A3(n_12670),
.B1(n_12672),
.B2(n_12668),
.B3(n_12663),
.Y(n_13027)
);

INVx1_ASAP7_75t_L g13028 ( 
.A(n_12373),
.Y(n_13028)
);

INVx1_ASAP7_75t_L g13029 ( 
.A(n_12566),
.Y(n_13029)
);

INVx1_ASAP7_75t_SL g13030 ( 
.A(n_12699),
.Y(n_13030)
);

INVx1_ASAP7_75t_L g13031 ( 
.A(n_12600),
.Y(n_13031)
);

INVx2_ASAP7_75t_L g13032 ( 
.A(n_12642),
.Y(n_13032)
);

INVx1_ASAP7_75t_L g13033 ( 
.A(n_12642),
.Y(n_13033)
);

AND2x2_ASAP7_75t_L g13034 ( 
.A(n_12666),
.B(n_8306),
.Y(n_13034)
);

NAND2xp5_ASAP7_75t_L g13035 ( 
.A(n_12647),
.B(n_8306),
.Y(n_13035)
);

INVxp67_ASAP7_75t_L g13036 ( 
.A(n_12298),
.Y(n_13036)
);

AND2x2_ASAP7_75t_L g13037 ( 
.A(n_12657),
.B(n_8306),
.Y(n_13037)
);

AND2x2_ASAP7_75t_L g13038 ( 
.A(n_12277),
.B(n_8306),
.Y(n_13038)
);

INVx1_ASAP7_75t_L g13039 ( 
.A(n_12647),
.Y(n_13039)
);

INVx1_ASAP7_75t_L g13040 ( 
.A(n_12443),
.Y(n_13040)
);

INVx1_ASAP7_75t_L g13041 ( 
.A(n_12444),
.Y(n_13041)
);

O2A1O1Ixp33_ASAP7_75t_L g13042 ( 
.A1(n_12530),
.A2(n_12545),
.B(n_12688),
.C(n_12684),
.Y(n_13042)
);

NAND2xp5_ASAP7_75t_L g13043 ( 
.A(n_12522),
.B(n_8306),
.Y(n_13043)
);

OR2x2_ASAP7_75t_L g13044 ( 
.A(n_12347),
.B(n_12555),
.Y(n_13044)
);

AND2x2_ASAP7_75t_L g13045 ( 
.A(n_12312),
.B(n_8323),
.Y(n_13045)
);

AOI21xp5_ASAP7_75t_L g13046 ( 
.A1(n_12508),
.A2(n_9786),
.B(n_7024),
.Y(n_13046)
);

INVx2_ASAP7_75t_L g13047 ( 
.A(n_12710),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_12472),
.Y(n_13048)
);

AOI22xp5_ASAP7_75t_L g13049 ( 
.A1(n_12601),
.A2(n_7567),
.B1(n_7619),
.B2(n_7553),
.Y(n_13049)
);

INVx2_ASAP7_75t_L g13050 ( 
.A(n_12541),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12450),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12454),
.Y(n_13052)
);

NAND4xp25_ASAP7_75t_L g13053 ( 
.A(n_12349),
.B(n_7278),
.C(n_7508),
.D(n_7345),
.Y(n_13053)
);

INVx1_ASAP7_75t_L g13054 ( 
.A(n_12461),
.Y(n_13054)
);

AND2x2_ASAP7_75t_L g13055 ( 
.A(n_12267),
.B(n_8323),
.Y(n_13055)
);

HB1xp67_ASAP7_75t_L g13056 ( 
.A(n_12510),
.Y(n_13056)
);

OR2x2_ASAP7_75t_L g13057 ( 
.A(n_12483),
.B(n_9110),
.Y(n_13057)
);

NAND2x1p5_ASAP7_75t_L g13058 ( 
.A(n_12581),
.B(n_7278),
.Y(n_13058)
);

AND2x2_ASAP7_75t_L g13059 ( 
.A(n_12517),
.B(n_8323),
.Y(n_13059)
);

AND2x2_ASAP7_75t_L g13060 ( 
.A(n_12518),
.B(n_12582),
.Y(n_13060)
);

NAND2xp5_ASAP7_75t_L g13061 ( 
.A(n_12467),
.B(n_8323),
.Y(n_13061)
);

NOR2xp33_ASAP7_75t_L g13062 ( 
.A(n_12314),
.B(n_7024),
.Y(n_13062)
);

OR2x2_ASAP7_75t_L g13063 ( 
.A(n_12556),
.B(n_9110),
.Y(n_13063)
);

INVx2_ASAP7_75t_L g13064 ( 
.A(n_12598),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12523),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_12477),
.Y(n_13066)
);

INVx1_ASAP7_75t_L g13067 ( 
.A(n_12481),
.Y(n_13067)
);

INVx1_ASAP7_75t_L g13068 ( 
.A(n_12484),
.Y(n_13068)
);

A2O1A1Ixp33_ASAP7_75t_L g13069 ( 
.A1(n_12304),
.A2(n_8323),
.B(n_8384),
.C(n_8375),
.Y(n_13069)
);

NAND2xp5_ASAP7_75t_L g13070 ( 
.A(n_12487),
.B(n_8375),
.Y(n_13070)
);

AND2x2_ASAP7_75t_L g13071 ( 
.A(n_12302),
.B(n_8375),
.Y(n_13071)
);

INVx1_ASAP7_75t_L g13072 ( 
.A(n_12492),
.Y(n_13072)
);

INVx2_ASAP7_75t_L g13073 ( 
.A(n_12457),
.Y(n_13073)
);

INVx1_ASAP7_75t_L g13074 ( 
.A(n_12494),
.Y(n_13074)
);

NAND2xp5_ASAP7_75t_L g13075 ( 
.A(n_12532),
.B(n_8375),
.Y(n_13075)
);

INVx1_ASAP7_75t_L g13076 ( 
.A(n_12377),
.Y(n_13076)
);

AND2x2_ASAP7_75t_L g13077 ( 
.A(n_12585),
.B(n_8375),
.Y(n_13077)
);

AND2x2_ASAP7_75t_L g13078 ( 
.A(n_12591),
.B(n_8384),
.Y(n_13078)
);

AOI21x1_ASAP7_75t_SL g13079 ( 
.A1(n_12325),
.A2(n_5990),
.B(n_5988),
.Y(n_13079)
);

AND2x2_ASAP7_75t_L g13080 ( 
.A(n_12594),
.B(n_8384),
.Y(n_13080)
);

NAND2x1p5_ASAP7_75t_L g13081 ( 
.A(n_12605),
.B(n_7149),
.Y(n_13081)
);

AND2x2_ASAP7_75t_L g13082 ( 
.A(n_12611),
.B(n_8384),
.Y(n_13082)
);

INVx1_ASAP7_75t_L g13083 ( 
.A(n_12533),
.Y(n_13083)
);

NAND2xp5_ASAP7_75t_L g13084 ( 
.A(n_12559),
.B(n_8384),
.Y(n_13084)
);

OAI21xp33_ASAP7_75t_L g13085 ( 
.A1(n_12619),
.A2(n_7020),
.B(n_7004),
.Y(n_13085)
);

NAND2x1_ASAP7_75t_L g13086 ( 
.A(n_12515),
.B(n_12631),
.Y(n_13086)
);

AND2x2_ASAP7_75t_L g13087 ( 
.A(n_12534),
.B(n_8392),
.Y(n_13087)
);

AND2x2_ASAP7_75t_L g13088 ( 
.A(n_12577),
.B(n_8392),
.Y(n_13088)
);

AND2x2_ASAP7_75t_L g13089 ( 
.A(n_12564),
.B(n_8392),
.Y(n_13089)
);

INVx2_ASAP7_75t_L g13090 ( 
.A(n_12460),
.Y(n_13090)
);

NAND2xp5_ASAP7_75t_L g13091 ( 
.A(n_12568),
.B(n_8392),
.Y(n_13091)
);

OR2x2_ASAP7_75t_L g13092 ( 
.A(n_12644),
.B(n_9123),
.Y(n_13092)
);

INVx1_ASAP7_75t_SL g13093 ( 
.A(n_12506),
.Y(n_13093)
);

INVx1_ASAP7_75t_L g13094 ( 
.A(n_12536),
.Y(n_13094)
);

INVx1_ASAP7_75t_L g13095 ( 
.A(n_12526),
.Y(n_13095)
);

NAND2xp5_ASAP7_75t_SL g13096 ( 
.A(n_12385),
.B(n_8392),
.Y(n_13096)
);

OR2x2_ASAP7_75t_L g13097 ( 
.A(n_12649),
.B(n_9123),
.Y(n_13097)
);

INVx1_ASAP7_75t_L g13098 ( 
.A(n_12535),
.Y(n_13098)
);

INVx1_ASAP7_75t_L g13099 ( 
.A(n_12540),
.Y(n_13099)
);

INVx2_ASAP7_75t_L g13100 ( 
.A(n_12478),
.Y(n_13100)
);

AND2x2_ASAP7_75t_L g13101 ( 
.A(n_12570),
.B(n_8414),
.Y(n_13101)
);

INVx1_ASAP7_75t_L g13102 ( 
.A(n_12602),
.Y(n_13102)
);

INVx1_ASAP7_75t_L g13103 ( 
.A(n_12448),
.Y(n_13103)
);

NAND2xp5_ASAP7_75t_L g13104 ( 
.A(n_12544),
.B(n_8414),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12455),
.Y(n_13105)
);

AND2x2_ASAP7_75t_L g13106 ( 
.A(n_12456),
.B(n_8414),
.Y(n_13106)
);

INVx2_ASAP7_75t_L g13107 ( 
.A(n_12482),
.Y(n_13107)
);

NAND2xp5_ASAP7_75t_L g13108 ( 
.A(n_12549),
.B(n_8414),
.Y(n_13108)
);

OAI21xp33_ASAP7_75t_L g13109 ( 
.A1(n_12620),
.A2(n_7020),
.B(n_7004),
.Y(n_13109)
);

AND2x4_ASAP7_75t_L g13110 ( 
.A(n_12554),
.B(n_8414),
.Y(n_13110)
);

OR2x2_ASAP7_75t_L g13111 ( 
.A(n_12495),
.B(n_9127),
.Y(n_13111)
);

INVx2_ASAP7_75t_L g13112 ( 
.A(n_12543),
.Y(n_13112)
);

INVx1_ASAP7_75t_L g13113 ( 
.A(n_12612),
.Y(n_13113)
);

INVxp67_ASAP7_75t_L g13114 ( 
.A(n_12695),
.Y(n_13114)
);

AND2x2_ASAP7_75t_L g13115 ( 
.A(n_12551),
.B(n_8422),
.Y(n_13115)
);

INVx2_ASAP7_75t_L g13116 ( 
.A(n_12618),
.Y(n_13116)
);

AND2x2_ASAP7_75t_L g13117 ( 
.A(n_12553),
.B(n_8422),
.Y(n_13117)
);

NAND2xp5_ASAP7_75t_L g13118 ( 
.A(n_12640),
.B(n_8422),
.Y(n_13118)
);

INVx1_ASAP7_75t_L g13119 ( 
.A(n_12392),
.Y(n_13119)
);

OR2x2_ASAP7_75t_L g13120 ( 
.A(n_12709),
.B(n_9127),
.Y(n_13120)
);

OR2x2_ASAP7_75t_L g13121 ( 
.A(n_12674),
.B(n_9133),
.Y(n_13121)
);

NAND2x1p5_ASAP7_75t_L g13122 ( 
.A(n_12410),
.B(n_7149),
.Y(n_13122)
);

INVx5_ASAP7_75t_L g13123 ( 
.A(n_12772),
.Y(n_13123)
);

INVx2_ASAP7_75t_SL g13124 ( 
.A(n_12827),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_13056),
.Y(n_13125)
);

NOR2xp33_ASAP7_75t_SL g13126 ( 
.A(n_12836),
.B(n_12680),
.Y(n_13126)
);

INVx1_ASAP7_75t_L g13127 ( 
.A(n_12799),
.Y(n_13127)
);

OAI22xp5_ASAP7_75t_L g13128 ( 
.A1(n_12833),
.A2(n_12345),
.B1(n_12417),
.B2(n_12414),
.Y(n_13128)
);

INVx1_ASAP7_75t_L g13129 ( 
.A(n_12723),
.Y(n_13129)
);

INVx2_ASAP7_75t_L g13130 ( 
.A(n_12839),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_12747),
.Y(n_13131)
);

NAND2xp5_ASAP7_75t_L g13132 ( 
.A(n_12782),
.B(n_12469),
.Y(n_13132)
);

INVx1_ASAP7_75t_SL g13133 ( 
.A(n_12762),
.Y(n_13133)
);

NOR2xp33_ASAP7_75t_L g13134 ( 
.A(n_12730),
.B(n_12648),
.Y(n_13134)
);

NOR2xp67_ASAP7_75t_L g13135 ( 
.A(n_12897),
.B(n_12697),
.Y(n_13135)
);

AND2x2_ASAP7_75t_L g13136 ( 
.A(n_12805),
.B(n_12552),
.Y(n_13136)
);

INVx1_ASAP7_75t_L g13137 ( 
.A(n_12912),
.Y(n_13137)
);

INVx1_ASAP7_75t_L g13138 ( 
.A(n_12937),
.Y(n_13138)
);

NOR2x1p5_ASAP7_75t_L g13139 ( 
.A(n_12738),
.B(n_12429),
.Y(n_13139)
);

HB1xp67_ASAP7_75t_L g13140 ( 
.A(n_12783),
.Y(n_13140)
);

INVx3_ASAP7_75t_L g13141 ( 
.A(n_12966),
.Y(n_13141)
);

INVx1_ASAP7_75t_L g13142 ( 
.A(n_12929),
.Y(n_13142)
);

INVx2_ASAP7_75t_L g13143 ( 
.A(n_13000),
.Y(n_13143)
);

NOR2x1p5_ASAP7_75t_SL g13144 ( 
.A(n_12765),
.B(n_12694),
.Y(n_13144)
);

INVx1_ASAP7_75t_L g13145 ( 
.A(n_12811),
.Y(n_13145)
);

OAI32xp33_ASAP7_75t_L g13146 ( 
.A1(n_12883),
.A2(n_12569),
.A3(n_12560),
.B1(n_12669),
.B2(n_12700),
.Y(n_13146)
);

AND2x4_ASAP7_75t_L g13147 ( 
.A(n_12869),
.B(n_12471),
.Y(n_13147)
);

AOI22xp5_ASAP7_75t_L g13148 ( 
.A1(n_12750),
.A2(n_12858),
.B1(n_12740),
.B2(n_12721),
.Y(n_13148)
);

AOI22xp5_ASAP7_75t_L g13149 ( 
.A1(n_12812),
.A2(n_12686),
.B1(n_12698),
.B2(n_12693),
.Y(n_13149)
);

INVx2_ASAP7_75t_L g13150 ( 
.A(n_12977),
.Y(n_13150)
);

NAND2xp5_ASAP7_75t_L g13151 ( 
.A(n_12913),
.B(n_12565),
.Y(n_13151)
);

OAI31xp33_ASAP7_75t_L g13152 ( 
.A1(n_12930),
.A2(n_12627),
.A3(n_12629),
.B(n_12625),
.Y(n_13152)
);

INVx1_ASAP7_75t_L g13153 ( 
.A(n_12720),
.Y(n_13153)
);

INVx1_ASAP7_75t_L g13154 ( 
.A(n_12724),
.Y(n_13154)
);

INVx3_ASAP7_75t_L g13155 ( 
.A(n_12871),
.Y(n_13155)
);

NAND2xp5_ASAP7_75t_L g13156 ( 
.A(n_12739),
.B(n_12650),
.Y(n_13156)
);

HB1xp67_ASAP7_75t_L g13157 ( 
.A(n_12746),
.Y(n_13157)
);

NAND2xp5_ASAP7_75t_L g13158 ( 
.A(n_12739),
.B(n_12651),
.Y(n_13158)
);

NOR2xp33_ASAP7_75t_L g13159 ( 
.A(n_12984),
.B(n_12529),
.Y(n_13159)
);

AOI21xp5_ASAP7_75t_L g13160 ( 
.A1(n_12872),
.A2(n_12439),
.B(n_12614),
.Y(n_13160)
);

INVx2_ASAP7_75t_L g13161 ( 
.A(n_12776),
.Y(n_13161)
);

O2A1O1Ixp5_ASAP7_75t_R g13162 ( 
.A1(n_12808),
.A2(n_12412),
.B(n_12428),
.C(n_12676),
.Y(n_13162)
);

NAND2x2_ASAP7_75t_L g13163 ( 
.A(n_12969),
.B(n_12713),
.Y(n_13163)
);

NAND2xp5_ASAP7_75t_L g13164 ( 
.A(n_12722),
.B(n_12607),
.Y(n_13164)
);

NOR2xp67_ASAP7_75t_L g13165 ( 
.A(n_12901),
.B(n_12633),
.Y(n_13165)
);

NOR2xp33_ASAP7_75t_L g13166 ( 
.A(n_12737),
.B(n_12621),
.Y(n_13166)
);

NOR2xp33_ASAP7_75t_L g13167 ( 
.A(n_12792),
.B(n_12691),
.Y(n_13167)
);

INVx1_ASAP7_75t_L g13168 ( 
.A(n_12728),
.Y(n_13168)
);

INVx1_ASAP7_75t_L g13169 ( 
.A(n_12716),
.Y(n_13169)
);

INVx2_ASAP7_75t_L g13170 ( 
.A(n_12927),
.Y(n_13170)
);

NAND4xp75_ASAP7_75t_SL g13171 ( 
.A(n_12981),
.B(n_12636),
.C(n_12603),
.D(n_12624),
.Y(n_13171)
);

INVx1_ASAP7_75t_L g13172 ( 
.A(n_12926),
.Y(n_13172)
);

NAND3xp33_ASAP7_75t_L g13173 ( 
.A(n_12796),
.B(n_12683),
.C(n_12661),
.Y(n_13173)
);

NAND2xp5_ASAP7_75t_L g13174 ( 
.A(n_12758),
.B(n_12658),
.Y(n_13174)
);

AND2x2_ASAP7_75t_L g13175 ( 
.A(n_12779),
.B(n_12829),
.Y(n_13175)
);

OAI32xp33_ASAP7_75t_L g13176 ( 
.A1(n_12838),
.A2(n_12653),
.A3(n_12655),
.B1(n_12572),
.B2(n_12660),
.Y(n_13176)
);

INVx3_ASAP7_75t_L g13177 ( 
.A(n_12852),
.Y(n_13177)
);

OR3x2_ASAP7_75t_L g13178 ( 
.A(n_12764),
.B(n_12706),
.C(n_12690),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_12875),
.Y(n_13179)
);

A2O1A1Ixp33_ASAP7_75t_L g13180 ( 
.A1(n_13042),
.A2(n_12613),
.B(n_12645),
.C(n_12637),
.Y(n_13180)
);

OAI32xp33_ASAP7_75t_L g13181 ( 
.A1(n_12888),
.A2(n_12703),
.A3(n_12712),
.B1(n_12692),
.B2(n_12679),
.Y(n_13181)
);

NAND2xp67_ASAP7_75t_SL g13182 ( 
.A(n_12850),
.B(n_12667),
.Y(n_13182)
);

INVx1_ASAP7_75t_L g13183 ( 
.A(n_12734),
.Y(n_13183)
);

INVx1_ASAP7_75t_L g13184 ( 
.A(n_12735),
.Y(n_13184)
);

INVx1_ASAP7_75t_SL g13185 ( 
.A(n_13010),
.Y(n_13185)
);

INVx1_ASAP7_75t_L g13186 ( 
.A(n_12741),
.Y(n_13186)
);

INVx1_ASAP7_75t_L g13187 ( 
.A(n_12718),
.Y(n_13187)
);

AND2x2_ASAP7_75t_L g13188 ( 
.A(n_12820),
.B(n_12685),
.Y(n_13188)
);

NAND2xp5_ASAP7_75t_L g13189 ( 
.A(n_13012),
.B(n_8422),
.Y(n_13189)
);

INVx2_ASAP7_75t_L g13190 ( 
.A(n_13026),
.Y(n_13190)
);

AND2x2_ASAP7_75t_L g13191 ( 
.A(n_12814),
.B(n_10070),
.Y(n_13191)
);

INVx1_ASAP7_75t_L g13192 ( 
.A(n_12798),
.Y(n_13192)
);

HB1xp67_ASAP7_75t_L g13193 ( 
.A(n_12983),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_12745),
.Y(n_13194)
);

INVxp67_ASAP7_75t_SL g13195 ( 
.A(n_12889),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_12824),
.Y(n_13196)
);

AOI33xp33_ASAP7_75t_L g13197 ( 
.A1(n_12788),
.A2(n_9143),
.A3(n_9134),
.B1(n_9146),
.B2(n_9142),
.B3(n_9133),
.Y(n_13197)
);

INVx2_ASAP7_75t_L g13198 ( 
.A(n_12972),
.Y(n_13198)
);

INVx1_ASAP7_75t_L g13199 ( 
.A(n_12761),
.Y(n_13199)
);

INVxp33_ASAP7_75t_L g13200 ( 
.A(n_12994),
.Y(n_13200)
);

NAND2x1_ASAP7_75t_SL g13201 ( 
.A(n_12849),
.B(n_10070),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_12974),
.Y(n_13202)
);

INVx3_ASAP7_75t_L g13203 ( 
.A(n_12809),
.Y(n_13203)
);

INVx2_ASAP7_75t_L g13204 ( 
.A(n_13005),
.Y(n_13204)
);

OAI31xp67_ASAP7_75t_L g13205 ( 
.A1(n_12837),
.A2(n_9142),
.A3(n_9143),
.B(n_9134),
.Y(n_13205)
);

NAND4xp25_ASAP7_75t_L g13206 ( 
.A(n_13062),
.B(n_7364),
.C(n_7387),
.D(n_7341),
.Y(n_13206)
);

INVx1_ASAP7_75t_L g13207 ( 
.A(n_12725),
.Y(n_13207)
);

NAND2xp5_ASAP7_75t_L g13208 ( 
.A(n_13030),
.B(n_8422),
.Y(n_13208)
);

INVx2_ASAP7_75t_L g13209 ( 
.A(n_12934),
.Y(n_13209)
);

NAND2xp5_ASAP7_75t_L g13210 ( 
.A(n_12809),
.B(n_8530),
.Y(n_13210)
);

INVx2_ASAP7_75t_SL g13211 ( 
.A(n_12934),
.Y(n_13211)
);

NAND2xp5_ASAP7_75t_L g13212 ( 
.A(n_12784),
.B(n_8530),
.Y(n_13212)
);

NAND2xp5_ASAP7_75t_L g13213 ( 
.A(n_12801),
.B(n_8530),
.Y(n_13213)
);

NAND2xp5_ASAP7_75t_L g13214 ( 
.A(n_12860),
.B(n_12863),
.Y(n_13214)
);

INVx2_ASAP7_75t_L g13215 ( 
.A(n_12893),
.Y(n_13215)
);

XOR2x2_ASAP7_75t_L g13216 ( 
.A(n_12881),
.B(n_7160),
.Y(n_13216)
);

INVx1_ASAP7_75t_L g13217 ( 
.A(n_13033),
.Y(n_13217)
);

AND2x2_ASAP7_75t_L g13218 ( 
.A(n_12830),
.B(n_10098),
.Y(n_13218)
);

AND2x2_ASAP7_75t_L g13219 ( 
.A(n_12825),
.B(n_10098),
.Y(n_13219)
);

AOI22xp5_ASAP7_75t_L g13220 ( 
.A1(n_13003),
.A2(n_7024),
.B1(n_7567),
.B2(n_7553),
.Y(n_13220)
);

AOI22xp5_ASAP7_75t_L g13221 ( 
.A1(n_12953),
.A2(n_7024),
.B1(n_7619),
.B2(n_7567),
.Y(n_13221)
);

OR3x2_ASAP7_75t_L g13222 ( 
.A(n_12908),
.B(n_7964),
.C(n_7024),
.Y(n_13222)
);

AOI22xp5_ASAP7_75t_L g13223 ( 
.A1(n_12964),
.A2(n_7681),
.B1(n_7781),
.B2(n_7619),
.Y(n_13223)
);

NOR2x1p5_ASAP7_75t_SL g13224 ( 
.A(n_12899),
.B(n_9146),
.Y(n_13224)
);

O2A1O1Ixp5_ASAP7_75t_R g13225 ( 
.A1(n_12846),
.A2(n_5990),
.B(n_6035),
.C(n_6026),
.Y(n_13225)
);

NOR2xp33_ASAP7_75t_L g13226 ( 
.A(n_12787),
.B(n_8409),
.Y(n_13226)
);

INVx1_ASAP7_75t_L g13227 ( 
.A(n_13039),
.Y(n_13227)
);

OAI21xp33_ASAP7_75t_SL g13228 ( 
.A1(n_12732),
.A2(n_9148),
.B(n_9147),
.Y(n_13228)
);

BUFx2_ASAP7_75t_L g13229 ( 
.A(n_12756),
.Y(n_13229)
);

AND2x2_ASAP7_75t_L g13230 ( 
.A(n_12823),
.B(n_10113),
.Y(n_13230)
);

NAND2xp5_ASAP7_75t_L g13231 ( 
.A(n_12806),
.B(n_8530),
.Y(n_13231)
);

NAND4xp25_ASAP7_75t_L g13232 ( 
.A(n_12804),
.B(n_7364),
.C(n_7387),
.D(n_7341),
.Y(n_13232)
);

AOI21xp33_ASAP7_75t_L g13233 ( 
.A1(n_12956),
.A2(n_10148),
.B(n_10113),
.Y(n_13233)
);

AND2x2_ASAP7_75t_L g13234 ( 
.A(n_12903),
.B(n_10148),
.Y(n_13234)
);

OAI332xp33_ASAP7_75t_L g13235 ( 
.A1(n_12919),
.A2(n_7713),
.A3(n_7356),
.B1(n_7372),
.B2(n_7266),
.B3(n_7458),
.C1(n_7581),
.C2(n_7530),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_13024),
.Y(n_13236)
);

NOR2x1_ASAP7_75t_L g13237 ( 
.A(n_12715),
.B(n_10152),
.Y(n_13237)
);

INVx1_ASAP7_75t_L g13238 ( 
.A(n_12992),
.Y(n_13238)
);

INVx1_ASAP7_75t_L g13239 ( 
.A(n_12993),
.Y(n_13239)
);

NOR2x1_ASAP7_75t_L g13240 ( 
.A(n_12733),
.B(n_12905),
.Y(n_13240)
);

NAND2xp5_ASAP7_75t_L g13241 ( 
.A(n_12865),
.B(n_8530),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_12866),
.Y(n_13242)
);

AOI32xp33_ASAP7_75t_L g13243 ( 
.A1(n_12807),
.A2(n_8653),
.A3(n_8696),
.B1(n_8602),
.B2(n_8546),
.Y(n_13243)
);

OAI32xp33_ASAP7_75t_L g13244 ( 
.A1(n_12963),
.A2(n_13044),
.A3(n_12843),
.B1(n_12781),
.B2(n_12767),
.Y(n_13244)
);

OR2x2_ASAP7_75t_L g13245 ( 
.A(n_12980),
.B(n_9147),
.Y(n_13245)
);

NAND2xp5_ASAP7_75t_SL g13246 ( 
.A(n_13093),
.B(n_8546),
.Y(n_13246)
);

AND2x2_ASAP7_75t_L g13247 ( 
.A(n_12771),
.B(n_12753),
.Y(n_13247)
);

INVx1_ASAP7_75t_L g13248 ( 
.A(n_12851),
.Y(n_13248)
);

NAND2xp5_ASAP7_75t_SL g13249 ( 
.A(n_12975),
.B(n_12933),
.Y(n_13249)
);

AND2x4_ASAP7_75t_L g13250 ( 
.A(n_13017),
.B(n_8546),
.Y(n_13250)
);

AOI21xp5_ASAP7_75t_L g13251 ( 
.A1(n_12859),
.A2(n_12991),
.B(n_12731),
.Y(n_13251)
);

OAI22xp5_ASAP7_75t_L g13252 ( 
.A1(n_13036),
.A2(n_8546),
.B1(n_8653),
.B2(n_8602),
.Y(n_13252)
);

NAND2xp5_ASAP7_75t_L g13253 ( 
.A(n_12818),
.B(n_8546),
.Y(n_13253)
);

INVx2_ASAP7_75t_SL g13254 ( 
.A(n_12943),
.Y(n_13254)
);

INVx2_ASAP7_75t_L g13255 ( 
.A(n_12894),
.Y(n_13255)
);

NAND2xp5_ASAP7_75t_L g13256 ( 
.A(n_12826),
.B(n_8602),
.Y(n_13256)
);

OAI31xp33_ASAP7_75t_L g13257 ( 
.A1(n_12847),
.A2(n_8602),
.A3(n_8696),
.B(n_8653),
.Y(n_13257)
);

INVx1_ASAP7_75t_L g13258 ( 
.A(n_12856),
.Y(n_13258)
);

INVx1_ASAP7_75t_L g13259 ( 
.A(n_12810),
.Y(n_13259)
);

INVx1_ASAP7_75t_L g13260 ( 
.A(n_12821),
.Y(n_13260)
);

BUFx2_ASAP7_75t_L g13261 ( 
.A(n_12976),
.Y(n_13261)
);

INVx1_ASAP7_75t_L g13262 ( 
.A(n_12822),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_12729),
.B(n_10152),
.Y(n_13263)
);

OAI21xp33_ASAP7_75t_SL g13264 ( 
.A1(n_12794),
.A2(n_9157),
.B(n_9148),
.Y(n_13264)
);

NOR2xp67_ASAP7_75t_SL g13265 ( 
.A(n_12802),
.B(n_7375),
.Y(n_13265)
);

OR2x2_ASAP7_75t_L g13266 ( 
.A(n_12795),
.B(n_9157),
.Y(n_13266)
);

INVx1_ASAP7_75t_L g13267 ( 
.A(n_12864),
.Y(n_13267)
);

INVx2_ASAP7_75t_L g13268 ( 
.A(n_12894),
.Y(n_13268)
);

INVx1_ASAP7_75t_L g13269 ( 
.A(n_12867),
.Y(n_13269)
);

INVxp67_ASAP7_75t_SL g13270 ( 
.A(n_13086),
.Y(n_13270)
);

OR2x2_ASAP7_75t_L g13271 ( 
.A(n_12755),
.B(n_9162),
.Y(n_13271)
);

OR2x2_ASAP7_75t_L g13272 ( 
.A(n_12916),
.B(n_9162),
.Y(n_13272)
);

INVx1_ASAP7_75t_L g13273 ( 
.A(n_12874),
.Y(n_13273)
);

NAND2xp5_ASAP7_75t_L g13274 ( 
.A(n_12815),
.B(n_8602),
.Y(n_13274)
);

INVx2_ASAP7_75t_L g13275 ( 
.A(n_12909),
.Y(n_13275)
);

INVx1_ASAP7_75t_L g13276 ( 
.A(n_12816),
.Y(n_13276)
);

OAI22xp33_ASAP7_75t_L g13277 ( 
.A1(n_12748),
.A2(n_8653),
.B1(n_8708),
.B2(n_8696),
.Y(n_13277)
);

NAND4xp75_ASAP7_75t_SL g13278 ( 
.A(n_13020),
.B(n_10180),
.C(n_10254),
.D(n_10323),
.Y(n_13278)
);

INVx1_ASAP7_75t_L g13279 ( 
.A(n_12842),
.Y(n_13279)
);

AOI32xp33_ASAP7_75t_L g13280 ( 
.A1(n_12793),
.A2(n_8708),
.A3(n_8727),
.B1(n_8696),
.B2(n_8653),
.Y(n_13280)
);

AND2x4_ASAP7_75t_L g13281 ( 
.A(n_13032),
.B(n_12873),
.Y(n_13281)
);

INVx1_ASAP7_75t_L g13282 ( 
.A(n_12844),
.Y(n_13282)
);

NAND2xp5_ASAP7_75t_L g13283 ( 
.A(n_12941),
.B(n_12975),
.Y(n_13283)
);

INVx1_ASAP7_75t_L g13284 ( 
.A(n_12726),
.Y(n_13284)
);

INVxp33_ASAP7_75t_L g13285 ( 
.A(n_12887),
.Y(n_13285)
);

INVx2_ASAP7_75t_L g13286 ( 
.A(n_12909),
.Y(n_13286)
);

INVx2_ASAP7_75t_L g13287 ( 
.A(n_12900),
.Y(n_13287)
);

OR2x2_ASAP7_75t_L g13288 ( 
.A(n_12945),
.B(n_9166),
.Y(n_13288)
);

OAI22xp33_ASAP7_75t_L g13289 ( 
.A1(n_12777),
.A2(n_8696),
.B1(n_8727),
.B2(n_8708),
.Y(n_13289)
);

OA222x2_ASAP7_75t_L g13290 ( 
.A1(n_12989),
.A2(n_8708),
.B1(n_8727),
.B2(n_8779),
.C1(n_8743),
.C2(n_8735),
.Y(n_13290)
);

INVx2_ASAP7_75t_SL g13291 ( 
.A(n_12760),
.Y(n_13291)
);

OR2x6_ASAP7_75t_L g13292 ( 
.A(n_12785),
.B(n_8409),
.Y(n_13292)
);

NAND2x1p5_ASAP7_75t_L g13293 ( 
.A(n_12982),
.B(n_7149),
.Y(n_13293)
);

OR2x2_ASAP7_75t_L g13294 ( 
.A(n_12949),
.B(n_9166),
.Y(n_13294)
);

INVx1_ASAP7_75t_L g13295 ( 
.A(n_12749),
.Y(n_13295)
);

INVx3_ASAP7_75t_L g13296 ( 
.A(n_12886),
.Y(n_13296)
);

OAI32xp33_ASAP7_75t_L g13297 ( 
.A1(n_12813),
.A2(n_8727),
.A3(n_8743),
.B1(n_8735),
.B2(n_8708),
.Y(n_13297)
);

INVx1_ASAP7_75t_L g13298 ( 
.A(n_12751),
.Y(n_13298)
);

NAND2xp5_ASAP7_75t_L g13299 ( 
.A(n_12902),
.B(n_8727),
.Y(n_13299)
);

OR2x2_ASAP7_75t_L g13300 ( 
.A(n_12803),
.B(n_9180),
.Y(n_13300)
);

OAI22xp33_ASAP7_75t_L g13301 ( 
.A1(n_13049),
.A2(n_8735),
.B1(n_8779),
.B2(n_8743),
.Y(n_13301)
);

INVx2_ASAP7_75t_L g13302 ( 
.A(n_12910),
.Y(n_13302)
);

AOI22xp5_ASAP7_75t_L g13303 ( 
.A1(n_12855),
.A2(n_7781),
.B1(n_7681),
.B2(n_8735),
.Y(n_13303)
);

INVx3_ASAP7_75t_L g13304 ( 
.A(n_12896),
.Y(n_13304)
);

INVx2_ASAP7_75t_L g13305 ( 
.A(n_12915),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_12954),
.Y(n_13306)
);

AND2x2_ASAP7_75t_L g13307 ( 
.A(n_12791),
.B(n_12774),
.Y(n_13307)
);

INVx1_ASAP7_75t_L g13308 ( 
.A(n_12757),
.Y(n_13308)
);

NAND2xp5_ASAP7_75t_L g13309 ( 
.A(n_12923),
.B(n_8735),
.Y(n_13309)
);

INVx1_ASAP7_75t_L g13310 ( 
.A(n_12759),
.Y(n_13310)
);

AND2x2_ASAP7_75t_L g13311 ( 
.A(n_13045),
.B(n_10180),
.Y(n_13311)
);

OAI222xp33_ASAP7_75t_L g13312 ( 
.A1(n_12931),
.A2(n_8807),
.B1(n_8779),
.B2(n_8804),
.C1(n_8743),
.C2(n_7895),
.Y(n_13312)
);

INVx1_ASAP7_75t_L g13313 ( 
.A(n_12736),
.Y(n_13313)
);

HB1xp67_ASAP7_75t_L g13314 ( 
.A(n_12986),
.Y(n_13314)
);

INVx4_ASAP7_75t_L g13315 ( 
.A(n_12790),
.Y(n_13315)
);

INVx2_ASAP7_75t_L g13316 ( 
.A(n_12845),
.Y(n_13316)
);

INVx1_ASAP7_75t_L g13317 ( 
.A(n_12743),
.Y(n_13317)
);

INVx1_ASAP7_75t_L g13318 ( 
.A(n_12727),
.Y(n_13318)
);

NOR2xp33_ASAP7_75t_L g13319 ( 
.A(n_12817),
.B(n_8409),
.Y(n_13319)
);

INVx1_ASAP7_75t_L g13320 ( 
.A(n_12742),
.Y(n_13320)
);

INVx2_ASAP7_75t_L g13321 ( 
.A(n_12862),
.Y(n_13321)
);

INVx2_ASAP7_75t_L g13322 ( 
.A(n_12840),
.Y(n_13322)
);

AOI32xp33_ASAP7_75t_L g13323 ( 
.A1(n_12906),
.A2(n_8804),
.A3(n_8807),
.B1(n_8779),
.B2(n_8743),
.Y(n_13323)
);

OAI322xp33_ASAP7_75t_L g13324 ( 
.A1(n_12979),
.A2(n_8779),
.A3(n_8807),
.B1(n_8804),
.B2(n_9180),
.C1(n_9189),
.C2(n_9187),
.Y(n_13324)
);

INVx1_ASAP7_75t_L g13325 ( 
.A(n_12951),
.Y(n_13325)
);

OA222x2_ASAP7_75t_L g13326 ( 
.A1(n_12800),
.A2(n_8804),
.B1(n_8807),
.B2(n_7895),
.C1(n_7411),
.C2(n_6993),
.Y(n_13326)
);

AND2x2_ASAP7_75t_L g13327 ( 
.A(n_12834),
.B(n_10323),
.Y(n_13327)
);

AND2x4_ASAP7_75t_L g13328 ( 
.A(n_13047),
.B(n_8804),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_12952),
.Y(n_13329)
);

INVx1_ASAP7_75t_SL g13330 ( 
.A(n_13060),
.Y(n_13330)
);

INVx1_ASAP7_75t_L g13331 ( 
.A(n_12957),
.Y(n_13331)
);

OAI22xp5_ASAP7_75t_L g13332 ( 
.A1(n_12819),
.A2(n_8807),
.B1(n_7284),
.B2(n_7438),
.Y(n_13332)
);

INVx1_ASAP7_75t_L g13333 ( 
.A(n_12962),
.Y(n_13333)
);

INVx1_ASAP7_75t_SL g13334 ( 
.A(n_12744),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_12968),
.Y(n_13335)
);

NAND2xp5_ASAP7_75t_L g13336 ( 
.A(n_12790),
.B(n_12841),
.Y(n_13336)
);

AOI211xp5_ASAP7_75t_L g13337 ( 
.A1(n_12942),
.A2(n_5793),
.B(n_7020),
.C(n_7004),
.Y(n_13337)
);

INVx1_ASAP7_75t_L g13338 ( 
.A(n_12832),
.Y(n_13338)
);

INVx2_ASAP7_75t_L g13339 ( 
.A(n_13058),
.Y(n_13339)
);

AND2x2_ASAP7_75t_L g13340 ( 
.A(n_13055),
.B(n_10349),
.Y(n_13340)
);

INVx2_ASAP7_75t_SL g13341 ( 
.A(n_12935),
.Y(n_13341)
);

XNOR2x1_ASAP7_75t_L g13342 ( 
.A(n_12770),
.B(n_8721),
.Y(n_13342)
);

INVx1_ASAP7_75t_L g13343 ( 
.A(n_12835),
.Y(n_13343)
);

NAND2xp5_ASAP7_75t_L g13344 ( 
.A(n_12935),
.B(n_9499),
.Y(n_13344)
);

INVx2_ASAP7_75t_L g13345 ( 
.A(n_12831),
.Y(n_13345)
);

OA222x2_ASAP7_75t_L g13346 ( 
.A1(n_12895),
.A2(n_7385),
.B1(n_7353),
.B2(n_7405),
.C1(n_7381),
.C2(n_7251),
.Y(n_13346)
);

OAI22xp33_ASAP7_75t_L g13347 ( 
.A1(n_12763),
.A2(n_7284),
.B1(n_7438),
.B2(n_7149),
.Y(n_13347)
);

INVx1_ASAP7_75t_L g13348 ( 
.A(n_12717),
.Y(n_13348)
);

OR2x2_ASAP7_75t_L g13349 ( 
.A(n_12985),
.B(n_9187),
.Y(n_13349)
);

INVx2_ASAP7_75t_L g13350 ( 
.A(n_12831),
.Y(n_13350)
);

NOR2x1p5_ASAP7_75t_L g13351 ( 
.A(n_12828),
.B(n_7681),
.Y(n_13351)
);

AOI32xp33_ASAP7_75t_L g13352 ( 
.A1(n_13007),
.A2(n_7266),
.A3(n_7080),
.B1(n_7044),
.B2(n_6951),
.Y(n_13352)
);

NAND4xp75_ASAP7_75t_L g13353 ( 
.A(n_12752),
.B(n_10410),
.C(n_10419),
.D(n_10349),
.Y(n_13353)
);

NOR2xp33_ASAP7_75t_SL g13354 ( 
.A(n_13027),
.B(n_13064),
.Y(n_13354)
);

OR2x2_ASAP7_75t_L g13355 ( 
.A(n_12948),
.B(n_9189),
.Y(n_13355)
);

INVx1_ASAP7_75t_L g13356 ( 
.A(n_13031),
.Y(n_13356)
);

INVx1_ASAP7_75t_L g13357 ( 
.A(n_12848),
.Y(n_13357)
);

INVx2_ASAP7_75t_SL g13358 ( 
.A(n_12970),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_13038),
.B(n_10410),
.Y(n_13359)
);

INVx1_ASAP7_75t_SL g13360 ( 
.A(n_12754),
.Y(n_13360)
);

NAND2xp5_ASAP7_75t_L g13361 ( 
.A(n_12999),
.B(n_9499),
.Y(n_13361)
);

OAI322xp33_ASAP7_75t_L g13362 ( 
.A1(n_12961),
.A2(n_9221),
.A3(n_9197),
.B1(n_9228),
.B2(n_9230),
.C1(n_9203),
.C2(n_9190),
.Y(n_13362)
);

AND2x2_ASAP7_75t_L g13363 ( 
.A(n_13071),
.B(n_10419),
.Y(n_13363)
);

AOI32xp33_ASAP7_75t_L g13364 ( 
.A1(n_12990),
.A2(n_7080),
.A3(n_7044),
.B1(n_6951),
.B2(n_6808),
.Y(n_13364)
);

OR2x6_ASAP7_75t_L g13365 ( 
.A(n_12778),
.B(n_12940),
.Y(n_13365)
);

AOI322xp5_ASAP7_75t_L g13366 ( 
.A1(n_12797),
.A2(n_6999),
.A3(n_7190),
.B1(n_7327),
.B2(n_6926),
.C1(n_7458),
.C2(n_7450),
.Y(n_13366)
);

OR2x2_ASAP7_75t_L g13367 ( 
.A(n_13065),
.B(n_9190),
.Y(n_13367)
);

NAND2xp5_ASAP7_75t_L g13368 ( 
.A(n_12970),
.B(n_12988),
.Y(n_13368)
);

INVx1_ASAP7_75t_L g13369 ( 
.A(n_12971),
.Y(n_13369)
);

NAND4xp75_ASAP7_75t_SL g13370 ( 
.A(n_13034),
.B(n_9499),
.C(n_6564),
.D(n_6491),
.Y(n_13370)
);

OAI22xp5_ASAP7_75t_L g13371 ( 
.A1(n_13114),
.A2(n_7438),
.B1(n_7284),
.B2(n_7020),
.Y(n_13371)
);

INVx1_ASAP7_75t_L g13372 ( 
.A(n_12998),
.Y(n_13372)
);

INVx1_ASAP7_75t_L g13373 ( 
.A(n_12978),
.Y(n_13373)
);

INVx1_ASAP7_75t_L g13374 ( 
.A(n_12876),
.Y(n_13374)
);

BUFx2_ASAP7_75t_L g13375 ( 
.A(n_12965),
.Y(n_13375)
);

OAI33xp33_ASAP7_75t_L g13376 ( 
.A1(n_12766),
.A2(n_9228),
.A3(n_9203),
.B1(n_9230),
.B2(n_9221),
.B3(n_9197),
.Y(n_13376)
);

OR2x2_ASAP7_75t_L g13377 ( 
.A(n_12786),
.B(n_9233),
.Y(n_13377)
);

AND2x2_ASAP7_75t_L g13378 ( 
.A(n_13004),
.B(n_9233),
.Y(n_13378)
);

OR2x2_ASAP7_75t_L g13379 ( 
.A(n_12789),
.B(n_9236),
.Y(n_13379)
);

XNOR2x2_ASAP7_75t_L g13380 ( 
.A(n_12914),
.B(n_7450),
.Y(n_13380)
);

XOR2x2_ASAP7_75t_L g13381 ( 
.A(n_12857),
.B(n_7160),
.Y(n_13381)
);

AND2x2_ASAP7_75t_L g13382 ( 
.A(n_13021),
.B(n_9236),
.Y(n_13382)
);

OR2x2_ASAP7_75t_L g13383 ( 
.A(n_12880),
.B(n_9242),
.Y(n_13383)
);

INVx2_ASAP7_75t_L g13384 ( 
.A(n_13122),
.Y(n_13384)
);

INVxp67_ASAP7_75t_L g13385 ( 
.A(n_13089),
.Y(n_13385)
);

NAND2xp5_ASAP7_75t_L g13386 ( 
.A(n_12938),
.B(n_9242),
.Y(n_13386)
);

INVx1_ASAP7_75t_L g13387 ( 
.A(n_12907),
.Y(n_13387)
);

NAND2xp5_ASAP7_75t_L g13388 ( 
.A(n_12938),
.B(n_13040),
.Y(n_13388)
);

HB1xp67_ASAP7_75t_L g13389 ( 
.A(n_13029),
.Y(n_13389)
);

OAI31xp33_ASAP7_75t_L g13390 ( 
.A1(n_13081),
.A2(n_6880),
.A3(n_6915),
.B(n_6884),
.Y(n_13390)
);

OR2x2_ASAP7_75t_L g13391 ( 
.A(n_13041),
.B(n_9244),
.Y(n_13391)
);

AND2x2_ASAP7_75t_L g13392 ( 
.A(n_13021),
.B(n_9244),
.Y(n_13392)
);

NAND2xp5_ASAP7_75t_L g13393 ( 
.A(n_13051),
.B(n_9246),
.Y(n_13393)
);

INVx1_ASAP7_75t_L g13394 ( 
.A(n_13052),
.Y(n_13394)
);

INVx1_ASAP7_75t_L g13395 ( 
.A(n_13054),
.Y(n_13395)
);

NAND2xp5_ASAP7_75t_L g13396 ( 
.A(n_13066),
.B(n_9246),
.Y(n_13396)
);

INVx1_ASAP7_75t_L g13397 ( 
.A(n_13067),
.Y(n_13397)
);

XNOR2xp5_ASAP7_75t_L g13398 ( 
.A(n_13053),
.B(n_7369),
.Y(n_13398)
);

OAI22xp5_ASAP7_75t_L g13399 ( 
.A1(n_13095),
.A2(n_7438),
.B1(n_7284),
.B2(n_7020),
.Y(n_13399)
);

NOR4xp25_ASAP7_75t_L g13400 ( 
.A(n_12768),
.B(n_9255),
.C(n_9268),
.D(n_9249),
.Y(n_13400)
);

AOI22xp5_ASAP7_75t_SL g13401 ( 
.A1(n_13098),
.A2(n_7229),
.B1(n_7213),
.B2(n_7378),
.Y(n_13401)
);

A2O1A1Ixp33_ASAP7_75t_L g13402 ( 
.A1(n_13046),
.A2(n_8409),
.B(n_8496),
.C(n_8777),
.Y(n_13402)
);

AND2x2_ASAP7_75t_L g13403 ( 
.A(n_12920),
.B(n_9249),
.Y(n_13403)
);

AND2x2_ASAP7_75t_L g13404 ( 
.A(n_13068),
.B(n_9255),
.Y(n_13404)
);

OR2x2_ASAP7_75t_L g13405 ( 
.A(n_13072),
.B(n_9268),
.Y(n_13405)
);

INVx2_ASAP7_75t_L g13406 ( 
.A(n_12965),
.Y(n_13406)
);

OAI33xp33_ASAP7_75t_L g13407 ( 
.A1(n_12769),
.A2(n_9296),
.A3(n_9272),
.B1(n_9305),
.B2(n_9295),
.B3(n_9271),
.Y(n_13407)
);

INVx1_ASAP7_75t_L g13408 ( 
.A(n_13074),
.Y(n_13408)
);

OR2x2_ASAP7_75t_L g13409 ( 
.A(n_13105),
.B(n_9271),
.Y(n_13409)
);

INVx1_ASAP7_75t_SL g13410 ( 
.A(n_13101),
.Y(n_13410)
);

NAND2xp5_ASAP7_75t_L g13411 ( 
.A(n_13099),
.B(n_9272),
.Y(n_13411)
);

AOI22xp5_ASAP7_75t_L g13412 ( 
.A1(n_13025),
.A2(n_7781),
.B1(n_8496),
.B2(n_8409),
.Y(n_13412)
);

INVx1_ASAP7_75t_L g13413 ( 
.A(n_12773),
.Y(n_13413)
);

OAI22xp33_ASAP7_75t_L g13414 ( 
.A1(n_13019),
.A2(n_7438),
.B1(n_7020),
.B2(n_7030),
.Y(n_13414)
);

NOR2x1_ASAP7_75t_L g13415 ( 
.A(n_12775),
.B(n_9295),
.Y(n_13415)
);

AND2x2_ASAP7_75t_L g13416 ( 
.A(n_13048),
.B(n_9296),
.Y(n_13416)
);

AOI22xp5_ASAP7_75t_L g13417 ( 
.A1(n_13037),
.A2(n_8496),
.B1(n_7020),
.B2(n_7030),
.Y(n_13417)
);

AOI22xp5_ASAP7_75t_L g13418 ( 
.A1(n_13085),
.A2(n_8496),
.B1(n_7030),
.B2(n_7093),
.Y(n_13418)
);

NAND2x2_ASAP7_75t_L g13419 ( 
.A(n_12973),
.B(n_6425),
.Y(n_13419)
);

AOI322xp5_ASAP7_75t_L g13420 ( 
.A1(n_12780),
.A2(n_7190),
.A3(n_7327),
.B1(n_6999),
.B2(n_7621),
.C1(n_7581),
.C2(n_7530),
.Y(n_13420)
);

AND2x2_ASAP7_75t_L g13421 ( 
.A(n_13073),
.B(n_9305),
.Y(n_13421)
);

OR2x2_ASAP7_75t_L g13422 ( 
.A(n_12967),
.B(n_9307),
.Y(n_13422)
);

OAI211xp5_ASAP7_75t_SL g13423 ( 
.A1(n_13103),
.A2(n_7395),
.B(n_7412),
.C(n_7367),
.Y(n_13423)
);

INVx2_ASAP7_75t_L g13424 ( 
.A(n_13016),
.Y(n_13424)
);

INVx2_ASAP7_75t_L g13425 ( 
.A(n_13014),
.Y(n_13425)
);

A2O1A1Ixp33_ASAP7_75t_L g13426 ( 
.A1(n_12861),
.A2(n_8496),
.B(n_8777),
.C(n_8370),
.Y(n_13426)
);

NOR2xp67_ASAP7_75t_L g13427 ( 
.A(n_12868),
.B(n_9307),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_12960),
.Y(n_13428)
);

INVx1_ASAP7_75t_L g13429 ( 
.A(n_12904),
.Y(n_13429)
);

INVx1_ASAP7_75t_L g13430 ( 
.A(n_12924),
.Y(n_13430)
);

AND2x4_ASAP7_75t_L g13431 ( 
.A(n_13090),
.B(n_9309),
.Y(n_13431)
);

INVx1_ASAP7_75t_L g13432 ( 
.A(n_12950),
.Y(n_13432)
);

HB1xp67_ASAP7_75t_L g13433 ( 
.A(n_13100),
.Y(n_13433)
);

INVx2_ASAP7_75t_SL g13434 ( 
.A(n_13110),
.Y(n_13434)
);

NOR2xp33_ASAP7_75t_SL g13435 ( 
.A(n_12719),
.B(n_7364),
.Y(n_13435)
);

A2O1A1Ixp33_ASAP7_75t_L g13436 ( 
.A1(n_12917),
.A2(n_8496),
.B(n_8777),
.C(n_8370),
.Y(n_13436)
);

OAI22xp33_ASAP7_75t_L g13437 ( 
.A1(n_12997),
.A2(n_7030),
.B1(n_7093),
.B2(n_7004),
.Y(n_13437)
);

NAND2xp5_ASAP7_75t_L g13438 ( 
.A(n_13107),
.B(n_9309),
.Y(n_13438)
);

INVx1_ASAP7_75t_L g13439 ( 
.A(n_13092),
.Y(n_13439)
);

AOI32xp33_ASAP7_75t_L g13440 ( 
.A1(n_12877),
.A2(n_12885),
.A3(n_13023),
.B1(n_13078),
.B2(n_13077),
.Y(n_13440)
);

INVx2_ASAP7_75t_SL g13441 ( 
.A(n_13110),
.Y(n_13441)
);

AOI22xp5_ASAP7_75t_L g13442 ( 
.A1(n_13006),
.A2(n_13013),
.B1(n_12946),
.B2(n_13109),
.Y(n_13442)
);

NOR2x1_ASAP7_75t_L g13443 ( 
.A(n_12921),
.B(n_12922),
.Y(n_13443)
);

NAND2xp5_ASAP7_75t_L g13444 ( 
.A(n_12878),
.B(n_12882),
.Y(n_13444)
);

INVx1_ASAP7_75t_L g13445 ( 
.A(n_13097),
.Y(n_13445)
);

INVx2_ASAP7_75t_SL g13446 ( 
.A(n_13106),
.Y(n_13446)
);

OAI22xp33_ASAP7_75t_SL g13447 ( 
.A1(n_13096),
.A2(n_12879),
.B1(n_12911),
.B2(n_12854),
.Y(n_13447)
);

OA222x2_ASAP7_75t_L g13448 ( 
.A1(n_12925),
.A2(n_7385),
.B1(n_7353),
.B2(n_7405),
.C1(n_7381),
.C2(n_7251),
.Y(n_13448)
);

AND2x2_ASAP7_75t_L g13449 ( 
.A(n_13050),
.B(n_9310),
.Y(n_13449)
);

INVx1_ASAP7_75t_L g13450 ( 
.A(n_12918),
.Y(n_13450)
);

OAI32xp33_ASAP7_75t_L g13451 ( 
.A1(n_13008),
.A2(n_7086),
.A3(n_7087),
.B1(n_7044),
.B2(n_6808),
.Y(n_13451)
);

NAND5xp2_ASAP7_75t_L g13452 ( 
.A(n_13102),
.B(n_7408),
.C(n_7400),
.D(n_7332),
.E(n_7091),
.Y(n_13452)
);

AOI32xp33_ASAP7_75t_L g13453 ( 
.A1(n_13080),
.A2(n_7087),
.A3(n_7120),
.B1(n_7086),
.B2(n_7044),
.Y(n_13453)
);

INVx1_ASAP7_75t_L g13454 ( 
.A(n_12932),
.Y(n_13454)
);

INVx2_ASAP7_75t_SL g13455 ( 
.A(n_13059),
.Y(n_13455)
);

INVx1_ASAP7_75t_L g13456 ( 
.A(n_12939),
.Y(n_13456)
);

NAND4xp75_ASAP7_75t_L g13457 ( 
.A(n_12959),
.B(n_9224),
.C(n_6696),
.D(n_6817),
.Y(n_13457)
);

INVx1_ASAP7_75t_L g13458 ( 
.A(n_12928),
.Y(n_13458)
);

AND2x2_ASAP7_75t_L g13459 ( 
.A(n_13116),
.B(n_13112),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_12936),
.Y(n_13460)
);

OAI31xp33_ASAP7_75t_L g13461 ( 
.A1(n_13113),
.A2(n_6884),
.A3(n_6915),
.B(n_6880),
.Y(n_13461)
);

INVx2_ASAP7_75t_L g13462 ( 
.A(n_13087),
.Y(n_13462)
);

OAI22xp33_ASAP7_75t_L g13463 ( 
.A1(n_12996),
.A2(n_7030),
.B1(n_7093),
.B2(n_7004),
.Y(n_13463)
);

OAI21xp33_ASAP7_75t_L g13464 ( 
.A1(n_13075),
.A2(n_9321),
.B(n_9310),
.Y(n_13464)
);

INVx1_ASAP7_75t_L g13465 ( 
.A(n_12947),
.Y(n_13465)
);

INVx1_ASAP7_75t_L g13466 ( 
.A(n_12955),
.Y(n_13466)
);

NAND2x1_ASAP7_75t_SL g13467 ( 
.A(n_12987),
.B(n_9321),
.Y(n_13467)
);

AOI32xp33_ASAP7_75t_L g13468 ( 
.A1(n_13082),
.A2(n_7120),
.A3(n_7184),
.B1(n_7087),
.B2(n_7086),
.Y(n_13468)
);

INVx2_ASAP7_75t_SL g13469 ( 
.A(n_13115),
.Y(n_13469)
);

NAND2xp5_ASAP7_75t_L g13470 ( 
.A(n_12890),
.B(n_9330),
.Y(n_13470)
);

INVx1_ASAP7_75t_L g13471 ( 
.A(n_12891),
.Y(n_13471)
);

OAI322xp33_ASAP7_75t_L g13472 ( 
.A1(n_12944),
.A2(n_9359),
.A3(n_9341),
.B1(n_9361),
.B2(n_9373),
.C1(n_9346),
.C2(n_9330),
.Y(n_13472)
);

INVx1_ASAP7_75t_L g13473 ( 
.A(n_12898),
.Y(n_13473)
);

O2A1O1Ixp33_ASAP7_75t_L g13474 ( 
.A1(n_12884),
.A2(n_9346),
.B(n_9359),
.C(n_9341),
.Y(n_13474)
);

NAND2xp5_ASAP7_75t_L g13475 ( 
.A(n_13117),
.B(n_9361),
.Y(n_13475)
);

O2A1O1Ixp33_ASAP7_75t_L g13476 ( 
.A1(n_12892),
.A2(n_9374),
.B(n_9378),
.C(n_9373),
.Y(n_13476)
);

INVx1_ASAP7_75t_L g13477 ( 
.A(n_13084),
.Y(n_13477)
);

INVx1_ASAP7_75t_L g13478 ( 
.A(n_13091),
.Y(n_13478)
);

INVx1_ASAP7_75t_L g13479 ( 
.A(n_13104),
.Y(n_13479)
);

OAI31xp33_ASAP7_75t_L g13480 ( 
.A1(n_13069),
.A2(n_6944),
.A3(n_7393),
.B(n_7304),
.Y(n_13480)
);

INVx1_ASAP7_75t_L g13481 ( 
.A(n_13108),
.Y(n_13481)
);

AND2x4_ASAP7_75t_L g13482 ( 
.A(n_12987),
.B(n_9374),
.Y(n_13482)
);

INVx1_ASAP7_75t_L g13483 ( 
.A(n_12853),
.Y(n_13483)
);

AOI22xp5_ASAP7_75t_L g13484 ( 
.A1(n_13088),
.A2(n_13028),
.B1(n_13022),
.B2(n_13018),
.Y(n_13484)
);

NOR2xp33_ASAP7_75t_L g13485 ( 
.A(n_13076),
.B(n_7424),
.Y(n_13485)
);

OR2x2_ASAP7_75t_L g13486 ( 
.A(n_13118),
.B(n_9378),
.Y(n_13486)
);

INVx1_ASAP7_75t_L g13487 ( 
.A(n_12870),
.Y(n_13487)
);

NAND2xp5_ASAP7_75t_L g13488 ( 
.A(n_13083),
.B(n_9384),
.Y(n_13488)
);

INVx2_ASAP7_75t_SL g13489 ( 
.A(n_13057),
.Y(n_13489)
);

OA222x2_ASAP7_75t_L g13490 ( 
.A1(n_12958),
.A2(n_7405),
.B1(n_7381),
.B2(n_7486),
.C1(n_7385),
.C2(n_7353),
.Y(n_13490)
);

INVxp67_ASAP7_75t_SL g13491 ( 
.A(n_13035),
.Y(n_13491)
);

INVx1_ASAP7_75t_L g13492 ( 
.A(n_13011),
.Y(n_13492)
);

A2O1A1Ixp33_ASAP7_75t_L g13493 ( 
.A1(n_13001),
.A2(n_8370),
.B(n_8313),
.C(n_8223),
.Y(n_13493)
);

INVx1_ASAP7_75t_SL g13494 ( 
.A(n_13043),
.Y(n_13494)
);

INVx1_ASAP7_75t_SL g13495 ( 
.A(n_13133),
.Y(n_13495)
);

AND2x2_ASAP7_75t_L g13496 ( 
.A(n_13175),
.B(n_13002),
.Y(n_13496)
);

HB1xp67_ASAP7_75t_L g13497 ( 
.A(n_13123),
.Y(n_13497)
);

XNOR2xp5_ASAP7_75t_L g13498 ( 
.A(n_13148),
.B(n_13342),
.Y(n_13498)
);

INVx1_ASAP7_75t_L g13499 ( 
.A(n_13224),
.Y(n_13499)
);

XNOR2xp5_ASAP7_75t_L g13500 ( 
.A(n_13247),
.B(n_13009),
.Y(n_13500)
);

INVx1_ASAP7_75t_L g13501 ( 
.A(n_13193),
.Y(n_13501)
);

INVx1_ASAP7_75t_L g13502 ( 
.A(n_13203),
.Y(n_13502)
);

INVx1_ASAP7_75t_L g13503 ( 
.A(n_13157),
.Y(n_13503)
);

XNOR2x2_ASAP7_75t_L g13504 ( 
.A(n_13240),
.B(n_13094),
.Y(n_13504)
);

XOR2x2_ASAP7_75t_L g13505 ( 
.A(n_13171),
.B(n_13015),
.Y(n_13505)
);

NOR2xp33_ASAP7_75t_L g13506 ( 
.A(n_13315),
.B(n_13119),
.Y(n_13506)
);

INVx2_ASAP7_75t_L g13507 ( 
.A(n_13201),
.Y(n_13507)
);

INVx2_ASAP7_75t_L g13508 ( 
.A(n_13123),
.Y(n_13508)
);

NAND2xp5_ASAP7_75t_L g13509 ( 
.A(n_13270),
.B(n_13281),
.Y(n_13509)
);

OAI22xp33_ASAP7_75t_L g13510 ( 
.A1(n_13229),
.A2(n_12995),
.B1(n_13070),
.B2(n_13061),
.Y(n_13510)
);

INVx2_ASAP7_75t_L g13511 ( 
.A(n_13123),
.Y(n_13511)
);

INVx1_ASAP7_75t_L g13512 ( 
.A(n_13336),
.Y(n_13512)
);

XOR2x2_ASAP7_75t_L g13513 ( 
.A(n_13485),
.B(n_13120),
.Y(n_13513)
);

INVx1_ASAP7_75t_L g13514 ( 
.A(n_13195),
.Y(n_13514)
);

OA22x2_ASAP7_75t_L g13515 ( 
.A1(n_13220),
.A2(n_13079),
.B1(n_13111),
.B2(n_9388),
.Y(n_13515)
);

XOR2x2_ASAP7_75t_L g13516 ( 
.A(n_13398),
.B(n_13063),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_13156),
.Y(n_13517)
);

INVx2_ASAP7_75t_SL g13518 ( 
.A(n_13155),
.Y(n_13518)
);

XNOR2xp5_ASAP7_75t_L g13519 ( 
.A(n_13185),
.B(n_13121),
.Y(n_13519)
);

OA22x2_ASAP7_75t_L g13520 ( 
.A1(n_13124),
.A2(n_9388),
.B1(n_9390),
.B2(n_9384),
.Y(n_13520)
);

OAI22xp33_ASAP7_75t_L g13521 ( 
.A1(n_13354),
.A2(n_13126),
.B1(n_13163),
.B2(n_13141),
.Y(n_13521)
);

XOR2x2_ASAP7_75t_L g13522 ( 
.A(n_13307),
.B(n_7486),
.Y(n_13522)
);

INVx1_ASAP7_75t_L g13523 ( 
.A(n_13142),
.Y(n_13523)
);

INVx1_ASAP7_75t_SL g13524 ( 
.A(n_13261),
.Y(n_13524)
);

XNOR2xp5_ASAP7_75t_L g13525 ( 
.A(n_13139),
.B(n_7427),
.Y(n_13525)
);

NOR2xp33_ASAP7_75t_L g13526 ( 
.A(n_13423),
.B(n_7525),
.Y(n_13526)
);

XNOR2xp5_ASAP7_75t_L g13527 ( 
.A(n_13131),
.B(n_7519),
.Y(n_13527)
);

XNOR2x1_ASAP7_75t_L g13528 ( 
.A(n_13144),
.B(n_13330),
.Y(n_13528)
);

INVx1_ASAP7_75t_L g13529 ( 
.A(n_13281),
.Y(n_13529)
);

XOR2x2_ASAP7_75t_L g13530 ( 
.A(n_13249),
.B(n_7486),
.Y(n_13530)
);

AO22x1_ASAP7_75t_L g13531 ( 
.A1(n_13147),
.A2(n_9401),
.B1(n_9402),
.B2(n_9390),
.Y(n_13531)
);

XNOR2x1_ASAP7_75t_L g13532 ( 
.A(n_13136),
.B(n_8721),
.Y(n_13532)
);

INVxp67_ASAP7_75t_SL g13533 ( 
.A(n_13380),
.Y(n_13533)
);

INVx2_ASAP7_75t_L g13534 ( 
.A(n_13467),
.Y(n_13534)
);

INVx1_ASAP7_75t_L g13535 ( 
.A(n_13188),
.Y(n_13535)
);

XNOR2xp5_ASAP7_75t_L g13536 ( 
.A(n_13149),
.B(n_7543),
.Y(n_13536)
);

CKINVDCx16_ASAP7_75t_R g13537 ( 
.A(n_13433),
.Y(n_13537)
);

AND2x2_ASAP7_75t_L g13538 ( 
.A(n_13204),
.B(n_13215),
.Y(n_13538)
);

NAND2xp5_ASAP7_75t_L g13539 ( 
.A(n_13130),
.B(n_9401),
.Y(n_13539)
);

INVx1_ASAP7_75t_SL g13540 ( 
.A(n_13360),
.Y(n_13540)
);

XNOR2xp5_ASAP7_75t_L g13541 ( 
.A(n_13216),
.B(n_7611),
.Y(n_13541)
);

OAI22x1_ASAP7_75t_L g13542 ( 
.A1(n_13143),
.A2(n_9409),
.B1(n_9415),
.B2(n_9402),
.Y(n_13542)
);

XOR2x2_ASAP7_75t_L g13543 ( 
.A(n_13134),
.B(n_13226),
.Y(n_13543)
);

XOR2x2_ASAP7_75t_L g13544 ( 
.A(n_13162),
.B(n_7523),
.Y(n_13544)
);

XNOR2x2_ASAP7_75t_L g13545 ( 
.A(n_13173),
.B(n_13443),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_13140),
.Y(n_13546)
);

INVx1_ASAP7_75t_SL g13547 ( 
.A(n_13334),
.Y(n_13547)
);

NAND2xp5_ASAP7_75t_L g13548 ( 
.A(n_13341),
.B(n_9409),
.Y(n_13548)
);

XOR2x2_ASAP7_75t_L g13549 ( 
.A(n_13174),
.B(n_7523),
.Y(n_13549)
);

INVxp67_ASAP7_75t_SL g13550 ( 
.A(n_13389),
.Y(n_13550)
);

NAND2xp33_ASAP7_75t_R g13551 ( 
.A(n_13147),
.B(n_13375),
.Y(n_13551)
);

INVx1_ASAP7_75t_SL g13552 ( 
.A(n_13283),
.Y(n_13552)
);

AOI22xp5_ASAP7_75t_SL g13553 ( 
.A1(n_13259),
.A2(n_7229),
.B1(n_7213),
.B2(n_7634),
.Y(n_13553)
);

INVx2_ASAP7_75t_SL g13554 ( 
.A(n_13211),
.Y(n_13554)
);

XOR2x2_ASAP7_75t_L g13555 ( 
.A(n_13135),
.B(n_7523),
.Y(n_13555)
);

AND2x4_ASAP7_75t_L g13556 ( 
.A(n_13190),
.B(n_7531),
.Y(n_13556)
);

INVx2_ASAP7_75t_L g13557 ( 
.A(n_13170),
.Y(n_13557)
);

INVxp67_ASAP7_75t_L g13558 ( 
.A(n_13435),
.Y(n_13558)
);

XNOR2x2_ASAP7_75t_L g13559 ( 
.A(n_13160),
.B(n_9415),
.Y(n_13559)
);

OA22x2_ASAP7_75t_L g13560 ( 
.A1(n_13221),
.A2(n_9421),
.B1(n_9428),
.B2(n_9419),
.Y(n_13560)
);

OR2x2_ASAP7_75t_L g13561 ( 
.A(n_13125),
.B(n_9419),
.Y(n_13561)
);

AND2x2_ASAP7_75t_L g13562 ( 
.A(n_13150),
.B(n_9421),
.Y(n_13562)
);

INVx1_ASAP7_75t_L g13563 ( 
.A(n_13209),
.Y(n_13563)
);

XOR2x2_ASAP7_75t_L g13564 ( 
.A(n_13151),
.B(n_7531),
.Y(n_13564)
);

NOR2xp33_ASAP7_75t_L g13565 ( 
.A(n_13127),
.B(n_7555),
.Y(n_13565)
);

INVx1_ASAP7_75t_SL g13566 ( 
.A(n_13263),
.Y(n_13566)
);

INVx1_ASAP7_75t_L g13567 ( 
.A(n_13255),
.Y(n_13567)
);

INVxp67_ASAP7_75t_L g13568 ( 
.A(n_13314),
.Y(n_13568)
);

XOR2xp5_ASAP7_75t_L g13569 ( 
.A(n_13178),
.B(n_7640),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_L g13570 ( 
.A(n_13207),
.B(n_9428),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_13268),
.Y(n_13571)
);

INVx1_ASAP7_75t_L g13572 ( 
.A(n_13275),
.Y(n_13572)
);

XNOR2xp5_ASAP7_75t_L g13573 ( 
.A(n_13232),
.B(n_7682),
.Y(n_13573)
);

INVx3_ASAP7_75t_SL g13574 ( 
.A(n_13365),
.Y(n_13574)
);

INVx2_ASAP7_75t_L g13575 ( 
.A(n_13286),
.Y(n_13575)
);

INVx1_ASAP7_75t_L g13576 ( 
.A(n_13183),
.Y(n_13576)
);

XNOR2x2_ASAP7_75t_L g13577 ( 
.A(n_13158),
.B(n_9432),
.Y(n_13577)
);

AOI22xp5_ASAP7_75t_L g13578 ( 
.A1(n_13161),
.A2(n_7752),
.B1(n_8456),
.B2(n_7093),
.Y(n_13578)
);

INVx1_ASAP7_75t_L g13579 ( 
.A(n_13287),
.Y(n_13579)
);

XOR2xp5_ASAP7_75t_L g13580 ( 
.A(n_13222),
.B(n_7698),
.Y(n_13580)
);

INVx1_ASAP7_75t_L g13581 ( 
.A(n_13302),
.Y(n_13581)
);

NOR2xp33_ASAP7_75t_L g13582 ( 
.A(n_13296),
.B(n_7653),
.Y(n_13582)
);

INVx1_ASAP7_75t_SL g13583 ( 
.A(n_13459),
.Y(n_13583)
);

AOI22x1_ASAP7_75t_SL g13584 ( 
.A1(n_13129),
.A2(n_9441),
.B1(n_9444),
.B2(n_9432),
.Y(n_13584)
);

XOR2x2_ASAP7_75t_L g13585 ( 
.A(n_13164),
.B(n_7531),
.Y(n_13585)
);

INVx1_ASAP7_75t_L g13586 ( 
.A(n_13305),
.Y(n_13586)
);

CKINVDCx5p33_ASAP7_75t_R g13587 ( 
.A(n_13365),
.Y(n_13587)
);

INVxp67_ASAP7_75t_L g13588 ( 
.A(n_13167),
.Y(n_13588)
);

XOR2x2_ASAP7_75t_L g13589 ( 
.A(n_13319),
.B(n_13159),
.Y(n_13589)
);

XOR2xp5_ASAP7_75t_L g13590 ( 
.A(n_13128),
.B(n_6425),
.Y(n_13590)
);

INVx1_ASAP7_75t_L g13591 ( 
.A(n_13316),
.Y(n_13591)
);

NAND2xp5_ASAP7_75t_L g13592 ( 
.A(n_13304),
.B(n_9441),
.Y(n_13592)
);

INVx2_ASAP7_75t_SL g13593 ( 
.A(n_13250),
.Y(n_13593)
);

INVx1_ASAP7_75t_SL g13594 ( 
.A(n_13410),
.Y(n_13594)
);

INVx8_ASAP7_75t_L g13595 ( 
.A(n_13177),
.Y(n_13595)
);

INVx1_ASAP7_75t_L g13596 ( 
.A(n_13321),
.Y(n_13596)
);

INVx1_ASAP7_75t_L g13597 ( 
.A(n_13322),
.Y(n_13597)
);

INVxp67_ASAP7_75t_L g13598 ( 
.A(n_13166),
.Y(n_13598)
);

INVx1_ASAP7_75t_L g13599 ( 
.A(n_13198),
.Y(n_13599)
);

NOR2xp33_ASAP7_75t_L g13600 ( 
.A(n_13145),
.B(n_7710),
.Y(n_13600)
);

OA22x2_ASAP7_75t_L g13601 ( 
.A1(n_13303),
.A2(n_9452),
.B1(n_9464),
.B2(n_9444),
.Y(n_13601)
);

INVx5_ASAP7_75t_L g13602 ( 
.A(n_13291),
.Y(n_13602)
);

AND2x2_ASAP7_75t_L g13603 ( 
.A(n_13202),
.B(n_9452),
.Y(n_13603)
);

INVxp67_ASAP7_75t_L g13604 ( 
.A(n_13358),
.Y(n_13604)
);

INVx1_ASAP7_75t_SL g13605 ( 
.A(n_13327),
.Y(n_13605)
);

XNOR2xp5_ASAP7_75t_L g13606 ( 
.A(n_13351),
.B(n_7536),
.Y(n_13606)
);

INVxp33_ASAP7_75t_SL g13607 ( 
.A(n_13265),
.Y(n_13607)
);

INVx4_ASAP7_75t_L g13608 ( 
.A(n_13339),
.Y(n_13608)
);

BUFx3_ASAP7_75t_L g13609 ( 
.A(n_13236),
.Y(n_13609)
);

INVx2_ASAP7_75t_L g13610 ( 
.A(n_13434),
.Y(n_13610)
);

INVxp67_ASAP7_75t_L g13611 ( 
.A(n_13210),
.Y(n_13611)
);

NOR2x1_ASAP7_75t_L g13612 ( 
.A(n_13182),
.B(n_9464),
.Y(n_13612)
);

INVx1_ASAP7_75t_L g13613 ( 
.A(n_13217),
.Y(n_13613)
);

INVx1_ASAP7_75t_L g13614 ( 
.A(n_13227),
.Y(n_13614)
);

INVx2_ASAP7_75t_L g13615 ( 
.A(n_13441),
.Y(n_13615)
);

INVx2_ASAP7_75t_L g13616 ( 
.A(n_13250),
.Y(n_13616)
);

INVx1_ASAP7_75t_L g13617 ( 
.A(n_13137),
.Y(n_13617)
);

XNOR2x2_ASAP7_75t_L g13618 ( 
.A(n_13237),
.B(n_9478),
.Y(n_13618)
);

INVx1_ASAP7_75t_SL g13619 ( 
.A(n_13234),
.Y(n_13619)
);

XOR2xp5_ASAP7_75t_L g13620 ( 
.A(n_13200),
.B(n_6425),
.Y(n_13620)
);

INVx1_ASAP7_75t_SL g13621 ( 
.A(n_13368),
.Y(n_13621)
);

INVxp67_ASAP7_75t_L g13622 ( 
.A(n_13388),
.Y(n_13622)
);

INVx1_ASAP7_75t_L g13623 ( 
.A(n_13138),
.Y(n_13623)
);

INVx1_ASAP7_75t_L g13624 ( 
.A(n_13238),
.Y(n_13624)
);

INVx1_ASAP7_75t_SL g13625 ( 
.A(n_13242),
.Y(n_13625)
);

AND2x2_ASAP7_75t_L g13626 ( 
.A(n_13239),
.B(n_9478),
.Y(n_13626)
);

INVx1_ASAP7_75t_SL g13627 ( 
.A(n_13248),
.Y(n_13627)
);

INVx2_ASAP7_75t_SL g13628 ( 
.A(n_13293),
.Y(n_13628)
);

OA22x2_ASAP7_75t_L g13629 ( 
.A1(n_13223),
.A2(n_9491),
.B1(n_9495),
.B2(n_9480),
.Y(n_13629)
);

INVx2_ASAP7_75t_L g13630 ( 
.A(n_13191),
.Y(n_13630)
);

XOR2xp5_ASAP7_75t_L g13631 ( 
.A(n_13285),
.B(n_6442),
.Y(n_13631)
);

INVxp67_ASAP7_75t_L g13632 ( 
.A(n_13189),
.Y(n_13632)
);

XOR2x2_ASAP7_75t_L g13633 ( 
.A(n_13165),
.B(n_7536),
.Y(n_13633)
);

INVx1_ASAP7_75t_L g13634 ( 
.A(n_13258),
.Y(n_13634)
);

AOI22xp5_ASAP7_75t_L g13635 ( 
.A1(n_13254),
.A2(n_8456),
.B1(n_7093),
.B2(n_7115),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_13132),
.Y(n_13636)
);

INVxp67_ASAP7_75t_L g13637 ( 
.A(n_13208),
.Y(n_13637)
);

INVxp67_ASAP7_75t_L g13638 ( 
.A(n_13212),
.Y(n_13638)
);

INVx1_ASAP7_75t_L g13639 ( 
.A(n_13214),
.Y(n_13639)
);

AOI22xp5_ASAP7_75t_L g13640 ( 
.A1(n_13192),
.A2(n_8456),
.B1(n_7093),
.B2(n_7115),
.Y(n_13640)
);

OAI22x1_ASAP7_75t_L g13641 ( 
.A1(n_13313),
.A2(n_9491),
.B1(n_9495),
.B2(n_9480),
.Y(n_13641)
);

OAI22xp5_ASAP7_75t_L g13642 ( 
.A1(n_13412),
.A2(n_13419),
.B1(n_13199),
.B2(n_13417),
.Y(n_13642)
);

XNOR2x1_ASAP7_75t_L g13643 ( 
.A(n_13345),
.B(n_6442),
.Y(n_13643)
);

INVxp67_ASAP7_75t_L g13644 ( 
.A(n_13320),
.Y(n_13644)
);

INVx2_ASAP7_75t_L g13645 ( 
.A(n_13230),
.Y(n_13645)
);

AND2x2_ASAP7_75t_L g13646 ( 
.A(n_13350),
.B(n_9498),
.Y(n_13646)
);

INVx2_ASAP7_75t_SL g13647 ( 
.A(n_13328),
.Y(n_13647)
);

XNOR2xp5_ASAP7_75t_L g13648 ( 
.A(n_13484),
.B(n_7536),
.Y(n_13648)
);

INVx1_ASAP7_75t_SL g13649 ( 
.A(n_13266),
.Y(n_13649)
);

XNOR2xp5_ASAP7_75t_L g13650 ( 
.A(n_13442),
.B(n_7541),
.Y(n_13650)
);

INVxp67_ASAP7_75t_SL g13651 ( 
.A(n_13415),
.Y(n_13651)
);

INVxp67_ASAP7_75t_L g13652 ( 
.A(n_13184),
.Y(n_13652)
);

INVx1_ASAP7_75t_L g13653 ( 
.A(n_13186),
.Y(n_13653)
);

XNOR2xp5_ASAP7_75t_L g13654 ( 
.A(n_13206),
.B(n_7541),
.Y(n_13654)
);

XOR2x2_ASAP7_75t_L g13655 ( 
.A(n_13444),
.B(n_7541),
.Y(n_13655)
);

NOR2xp33_ASAP7_75t_L g13656 ( 
.A(n_13244),
.B(n_7720),
.Y(n_13656)
);

INVx2_ASAP7_75t_L g13657 ( 
.A(n_13219),
.Y(n_13657)
);

OA22x2_ASAP7_75t_L g13658 ( 
.A1(n_13455),
.A2(n_9501),
.B1(n_9506),
.B2(n_9498),
.Y(n_13658)
);

XOR2x2_ASAP7_75t_L g13659 ( 
.A(n_13179),
.B(n_7565),
.Y(n_13659)
);

AO22x2_ASAP7_75t_L g13660 ( 
.A1(n_13406),
.A2(n_9506),
.B1(n_9511),
.B2(n_9501),
.Y(n_13660)
);

OR2x2_ASAP7_75t_L g13661 ( 
.A(n_13469),
.B(n_9511),
.Y(n_13661)
);

XOR2xp5_ASAP7_75t_L g13662 ( 
.A(n_13172),
.B(n_6442),
.Y(n_13662)
);

XOR2x2_ASAP7_75t_L g13663 ( 
.A(n_13251),
.B(n_7565),
.Y(n_13663)
);

INVx1_ASAP7_75t_L g13664 ( 
.A(n_13429),
.Y(n_13664)
);

XNOR2x2_ASAP7_75t_L g13665 ( 
.A(n_13369),
.B(n_9513),
.Y(n_13665)
);

INVx1_ASAP7_75t_L g13666 ( 
.A(n_13430),
.Y(n_13666)
);

INVx2_ASAP7_75t_L g13667 ( 
.A(n_13328),
.Y(n_13667)
);

HB1xp67_ASAP7_75t_L g13668 ( 
.A(n_13218),
.Y(n_13668)
);

INVx1_ASAP7_75t_L g13669 ( 
.A(n_13432),
.Y(n_13669)
);

INVx1_ASAP7_75t_L g13670 ( 
.A(n_13428),
.Y(n_13670)
);

INVxp67_ASAP7_75t_L g13671 ( 
.A(n_13299),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_13187),
.Y(n_13672)
);

OR2x2_ASAP7_75t_L g13673 ( 
.A(n_13325),
.B(n_9513),
.Y(n_13673)
);

INVx1_ASAP7_75t_L g13674 ( 
.A(n_13194),
.Y(n_13674)
);

XOR2x2_ASAP7_75t_L g13675 ( 
.A(n_13246),
.B(n_7565),
.Y(n_13675)
);

XNOR2x1_ASAP7_75t_L g13676 ( 
.A(n_13494),
.B(n_6488),
.Y(n_13676)
);

INVxp67_ASAP7_75t_L g13677 ( 
.A(n_13309),
.Y(n_13677)
);

XOR2x2_ASAP7_75t_L g13678 ( 
.A(n_13447),
.B(n_7608),
.Y(n_13678)
);

NOR2x1_ASAP7_75t_L g13679 ( 
.A(n_13373),
.B(n_9518),
.Y(n_13679)
);

NOR2x1_ASAP7_75t_R g13680 ( 
.A(n_13317),
.B(n_7726),
.Y(n_13680)
);

INVx1_ASAP7_75t_L g13681 ( 
.A(n_13267),
.Y(n_13681)
);

XOR2xp5_ASAP7_75t_L g13682 ( 
.A(n_13338),
.B(n_6488),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_13269),
.Y(n_13683)
);

OA22x2_ASAP7_75t_L g13684 ( 
.A1(n_13446),
.A2(n_9520),
.B1(n_9524),
.B2(n_9518),
.Y(n_13684)
);

XNOR2x1_ASAP7_75t_L g13685 ( 
.A(n_13292),
.B(n_13425),
.Y(n_13685)
);

NAND2xp5_ASAP7_75t_L g13686 ( 
.A(n_13489),
.B(n_9520),
.Y(n_13686)
);

INVxp67_ASAP7_75t_L g13687 ( 
.A(n_13253),
.Y(n_13687)
);

INVx1_ASAP7_75t_L g13688 ( 
.A(n_13273),
.Y(n_13688)
);

XOR2x2_ASAP7_75t_L g13689 ( 
.A(n_13318),
.B(n_7608),
.Y(n_13689)
);

XNOR2xp5_ASAP7_75t_L g13690 ( 
.A(n_13401),
.B(n_7608),
.Y(n_13690)
);

INVxp67_ASAP7_75t_L g13691 ( 
.A(n_13256),
.Y(n_13691)
);

XNOR2x2_ASAP7_75t_L g13692 ( 
.A(n_13295),
.B(n_9524),
.Y(n_13692)
);

INVx1_ASAP7_75t_L g13693 ( 
.A(n_13329),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_13331),
.Y(n_13694)
);

XOR2x2_ASAP7_75t_L g13695 ( 
.A(n_13343),
.B(n_7637),
.Y(n_13695)
);

XNOR2x1_ASAP7_75t_L g13696 ( 
.A(n_13292),
.B(n_6488),
.Y(n_13696)
);

NOR2x1_ASAP7_75t_L g13697 ( 
.A(n_13483),
.B(n_9530),
.Y(n_13697)
);

INVx1_ASAP7_75t_SL g13698 ( 
.A(n_13245),
.Y(n_13698)
);

NOR2xp33_ASAP7_75t_L g13699 ( 
.A(n_13146),
.B(n_7742),
.Y(n_13699)
);

INVxp67_ASAP7_75t_L g13700 ( 
.A(n_13231),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_13333),
.Y(n_13701)
);

INVx1_ASAP7_75t_L g13702 ( 
.A(n_13335),
.Y(n_13702)
);

XOR2x2_ASAP7_75t_L g13703 ( 
.A(n_13284),
.B(n_7637),
.Y(n_13703)
);

INVx2_ASAP7_75t_SL g13704 ( 
.A(n_13431),
.Y(n_13704)
);

NAND2xp5_ASAP7_75t_L g13705 ( 
.A(n_13180),
.B(n_9530),
.Y(n_13705)
);

INVx2_ASAP7_75t_L g13706 ( 
.A(n_13311),
.Y(n_13706)
);

AOI22xp5_ASAP7_75t_SL g13707 ( 
.A1(n_13385),
.A2(n_7497),
.B1(n_7574),
.B2(n_7464),
.Y(n_13707)
);

INVx1_ASAP7_75t_L g13708 ( 
.A(n_13356),
.Y(n_13708)
);

INVx2_ASAP7_75t_SL g13709 ( 
.A(n_13431),
.Y(n_13709)
);

INVx1_ASAP7_75t_L g13710 ( 
.A(n_13357),
.Y(n_13710)
);

XNOR2xp5_ASAP7_75t_L g13711 ( 
.A(n_13381),
.B(n_7637),
.Y(n_13711)
);

OA22x2_ASAP7_75t_L g13712 ( 
.A1(n_13169),
.A2(n_9535),
.B1(n_9536),
.B2(n_9531),
.Y(n_13712)
);

OR2x2_ASAP7_75t_L g13713 ( 
.A(n_13260),
.B(n_9531),
.Y(n_13713)
);

BUFx3_ASAP7_75t_L g13714 ( 
.A(n_13262),
.Y(n_13714)
);

INVx2_ASAP7_75t_L g13715 ( 
.A(n_13359),
.Y(n_13715)
);

OAI22x1_ASAP7_75t_L g13716 ( 
.A1(n_13424),
.A2(n_9536),
.B1(n_9540),
.B2(n_9535),
.Y(n_13716)
);

AND2x2_ASAP7_75t_L g13717 ( 
.A(n_13462),
.B(n_9540),
.Y(n_13717)
);

XNOR2xp5_ASAP7_75t_L g13718 ( 
.A(n_13196),
.B(n_7639),
.Y(n_13718)
);

NOR2xp33_ASAP7_75t_L g13719 ( 
.A(n_13176),
.B(n_7364),
.Y(n_13719)
);

INVx1_ASAP7_75t_L g13720 ( 
.A(n_13306),
.Y(n_13720)
);

OAI22x1_ASAP7_75t_L g13721 ( 
.A1(n_13310),
.A2(n_9548),
.B1(n_9552),
.B2(n_9544),
.Y(n_13721)
);

NOR2xp33_ASAP7_75t_L g13722 ( 
.A(n_13181),
.B(n_7387),
.Y(n_13722)
);

NOR2xp33_ASAP7_75t_L g13723 ( 
.A(n_13439),
.B(n_7387),
.Y(n_13723)
);

OA22x2_ASAP7_75t_L g13724 ( 
.A1(n_13418),
.A2(n_9548),
.B1(n_9552),
.B2(n_9544),
.Y(n_13724)
);

INVxp67_ASAP7_75t_L g13725 ( 
.A(n_13241),
.Y(n_13725)
);

INVx2_ASAP7_75t_L g13726 ( 
.A(n_13340),
.Y(n_13726)
);

OA22x2_ASAP7_75t_L g13727 ( 
.A1(n_13445),
.A2(n_9566),
.B1(n_9570),
.B2(n_9565),
.Y(n_13727)
);

HB1xp67_ASAP7_75t_L g13728 ( 
.A(n_13427),
.Y(n_13728)
);

XOR2x2_ASAP7_75t_L g13729 ( 
.A(n_13308),
.B(n_13274),
.Y(n_13729)
);

INVxp67_ASAP7_75t_L g13730 ( 
.A(n_13213),
.Y(n_13730)
);

XNOR2xp5_ASAP7_75t_L g13731 ( 
.A(n_13372),
.B(n_7639),
.Y(n_13731)
);

NAND2xp5_ASAP7_75t_L g13732 ( 
.A(n_13152),
.B(n_9565),
.Y(n_13732)
);

NAND2xp5_ASAP7_75t_L g13733 ( 
.A(n_13440),
.B(n_9566),
.Y(n_13733)
);

XNOR2xp5_ASAP7_75t_L g13734 ( 
.A(n_13394),
.B(n_7639),
.Y(n_13734)
);

AND2x2_ASAP7_75t_L g13735 ( 
.A(n_13395),
.B(n_9570),
.Y(n_13735)
);

INVx1_ASAP7_75t_L g13736 ( 
.A(n_13416),
.Y(n_13736)
);

NOR2x1_ASAP7_75t_L g13737 ( 
.A(n_13298),
.B(n_9575),
.Y(n_13737)
);

XOR2x2_ASAP7_75t_L g13738 ( 
.A(n_13471),
.B(n_7662),
.Y(n_13738)
);

NAND2xp5_ASAP7_75t_L g13739 ( 
.A(n_13473),
.B(n_9575),
.Y(n_13739)
);

AOI22xp5_ASAP7_75t_L g13740 ( 
.A1(n_13332),
.A2(n_8456),
.B1(n_7093),
.B2(n_7115),
.Y(n_13740)
);

HB1xp67_ASAP7_75t_L g13741 ( 
.A(n_13482),
.Y(n_13741)
);

INVx1_ASAP7_75t_SL g13742 ( 
.A(n_13421),
.Y(n_13742)
);

OA22x2_ASAP7_75t_L g13743 ( 
.A1(n_13397),
.A2(n_9595),
.B1(n_9599),
.B2(n_9580),
.Y(n_13743)
);

XNOR2x1_ASAP7_75t_L g13744 ( 
.A(n_13408),
.B(n_6488),
.Y(n_13744)
);

INVxp67_ASAP7_75t_L g13745 ( 
.A(n_13404),
.Y(n_13745)
);

AND2x2_ASAP7_75t_L g13746 ( 
.A(n_13492),
.B(n_9580),
.Y(n_13746)
);

XNOR2xp5_ASAP7_75t_L g13747 ( 
.A(n_13378),
.B(n_7662),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_13449),
.B(n_9595),
.Y(n_13748)
);

OR2x2_ASAP7_75t_L g13749 ( 
.A(n_13300),
.B(n_9599),
.Y(n_13749)
);

INVx1_ASAP7_75t_SL g13750 ( 
.A(n_13377),
.Y(n_13750)
);

XOR2x2_ASAP7_75t_L g13751 ( 
.A(n_13370),
.B(n_7662),
.Y(n_13751)
);

XNOR2xp5_ASAP7_75t_L g13752 ( 
.A(n_13348),
.B(n_7686),
.Y(n_13752)
);

NAND2xp5_ASAP7_75t_L g13753 ( 
.A(n_13153),
.B(n_9600),
.Y(n_13753)
);

XNOR2xp5_ASAP7_75t_L g13754 ( 
.A(n_13382),
.B(n_7686),
.Y(n_13754)
);

INVx1_ASAP7_75t_SL g13755 ( 
.A(n_13379),
.Y(n_13755)
);

XNOR2xp5_ASAP7_75t_L g13756 ( 
.A(n_13392),
.B(n_13487),
.Y(n_13756)
);

XNOR2xp5_ASAP7_75t_L g13757 ( 
.A(n_13413),
.B(n_7464),
.Y(n_13757)
);

INVx2_ASAP7_75t_L g13758 ( 
.A(n_13363),
.Y(n_13758)
);

INVx1_ASAP7_75t_L g13759 ( 
.A(n_13288),
.Y(n_13759)
);

NAND2xp5_ASAP7_75t_L g13760 ( 
.A(n_13154),
.B(n_9600),
.Y(n_13760)
);

INVx1_ASAP7_75t_L g13761 ( 
.A(n_13294),
.Y(n_13761)
);

INVx2_ASAP7_75t_L g13762 ( 
.A(n_13482),
.Y(n_13762)
);

INVx2_ASAP7_75t_SL g13763 ( 
.A(n_13367),
.Y(n_13763)
);

INVx1_ASAP7_75t_L g13764 ( 
.A(n_13355),
.Y(n_13764)
);

HB1xp67_ASAP7_75t_L g13765 ( 
.A(n_13278),
.Y(n_13765)
);

INVx2_ASAP7_75t_L g13766 ( 
.A(n_13422),
.Y(n_13766)
);

INVx2_ASAP7_75t_L g13767 ( 
.A(n_13383),
.Y(n_13767)
);

INVx1_ASAP7_75t_L g13768 ( 
.A(n_13168),
.Y(n_13768)
);

INVx2_ASAP7_75t_L g13769 ( 
.A(n_13272),
.Y(n_13769)
);

OA22x2_ASAP7_75t_L g13770 ( 
.A1(n_13384),
.A2(n_9607),
.B1(n_9619),
.B2(n_9602),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_13349),
.Y(n_13771)
);

INVxp67_ASAP7_75t_L g13772 ( 
.A(n_13271),
.Y(n_13772)
);

AND2x2_ASAP7_75t_L g13773 ( 
.A(n_13491),
.B(n_9602),
.Y(n_13773)
);

XOR2x2_ASAP7_75t_L g13774 ( 
.A(n_13438),
.B(n_13411),
.Y(n_13774)
);

INVx1_ASAP7_75t_L g13775 ( 
.A(n_13391),
.Y(n_13775)
);

INVx2_ASAP7_75t_SL g13776 ( 
.A(n_13405),
.Y(n_13776)
);

NOR2xp33_ASAP7_75t_L g13777 ( 
.A(n_13387),
.B(n_7491),
.Y(n_13777)
);

INVx1_ASAP7_75t_L g13778 ( 
.A(n_13409),
.Y(n_13778)
);

INVx2_ASAP7_75t_L g13779 ( 
.A(n_13403),
.Y(n_13779)
);

AND2x4_ASAP7_75t_L g13780 ( 
.A(n_13477),
.B(n_13478),
.Y(n_13780)
);

INVx2_ASAP7_75t_L g13781 ( 
.A(n_13353),
.Y(n_13781)
);

AND2x2_ASAP7_75t_L g13782 ( 
.A(n_13346),
.B(n_9607),
.Y(n_13782)
);

INVx1_ASAP7_75t_L g13783 ( 
.A(n_13279),
.Y(n_13783)
);

OA22x2_ASAP7_75t_L g13784 ( 
.A1(n_13454),
.A2(n_9620),
.B1(n_9635),
.B2(n_9619),
.Y(n_13784)
);

INVx2_ASAP7_75t_L g13785 ( 
.A(n_13486),
.Y(n_13785)
);

AND2x2_ASAP7_75t_L g13786 ( 
.A(n_13479),
.B(n_9620),
.Y(n_13786)
);

NAND2xp5_ASAP7_75t_L g13787 ( 
.A(n_13456),
.B(n_9635),
.Y(n_13787)
);

INVxp67_ASAP7_75t_L g13788 ( 
.A(n_13393),
.Y(n_13788)
);

INVx2_ASAP7_75t_SL g13789 ( 
.A(n_13396),
.Y(n_13789)
);

INVx1_ASAP7_75t_SL g13790 ( 
.A(n_13361),
.Y(n_13790)
);

INVx1_ASAP7_75t_L g13791 ( 
.A(n_13282),
.Y(n_13791)
);

AND2x2_ASAP7_75t_L g13792 ( 
.A(n_13481),
.B(n_9638),
.Y(n_13792)
);

INVx2_ASAP7_75t_SL g13793 ( 
.A(n_13470),
.Y(n_13793)
);

INVxp67_ASAP7_75t_SL g13794 ( 
.A(n_13386),
.Y(n_13794)
);

XOR2x2_ASAP7_75t_L g13795 ( 
.A(n_13450),
.B(n_7686),
.Y(n_13795)
);

INVx1_ASAP7_75t_SL g13796 ( 
.A(n_13475),
.Y(n_13796)
);

XOR2x2_ASAP7_75t_L g13797 ( 
.A(n_13458),
.B(n_7775),
.Y(n_13797)
);

XNOR2xp5_ASAP7_75t_L g13798 ( 
.A(n_13301),
.B(n_13374),
.Y(n_13798)
);

NAND2xp5_ASAP7_75t_L g13799 ( 
.A(n_13460),
.B(n_13465),
.Y(n_13799)
);

OAI22xp33_ASAP7_75t_SL g13800 ( 
.A1(n_13276),
.A2(n_9641),
.B1(n_9643),
.B2(n_9638),
.Y(n_13800)
);

INVx2_ASAP7_75t_L g13801 ( 
.A(n_13344),
.Y(n_13801)
);

INVx1_ASAP7_75t_L g13802 ( 
.A(n_13488),
.Y(n_13802)
);

XOR2x2_ASAP7_75t_L g13803 ( 
.A(n_13466),
.B(n_7775),
.Y(n_13803)
);

XNOR2xp5_ASAP7_75t_L g13804 ( 
.A(n_13400),
.B(n_7775),
.Y(n_13804)
);

XNOR2x2_ASAP7_75t_L g13805 ( 
.A(n_13252),
.B(n_9641),
.Y(n_13805)
);

NOR2xp33_ASAP7_75t_L g13806 ( 
.A(n_13235),
.B(n_7491),
.Y(n_13806)
);

AOI22xp33_ASAP7_75t_L g13807 ( 
.A1(n_13595),
.A2(n_13574),
.B1(n_13503),
.B2(n_13518),
.Y(n_13807)
);

INVx1_ASAP7_75t_L g13808 ( 
.A(n_13497),
.Y(n_13808)
);

AOI22xp5_ASAP7_75t_L g13809 ( 
.A1(n_13587),
.A2(n_13347),
.B1(n_13371),
.B2(n_13399),
.Y(n_13809)
);

OAI22xp5_ASAP7_75t_L g13810 ( 
.A1(n_13537),
.A2(n_13402),
.B1(n_13337),
.B2(n_13364),
.Y(n_13810)
);

NAND2xp5_ASAP7_75t_L g13811 ( 
.A(n_13602),
.B(n_13595),
.Y(n_13811)
);

INVx4_ASAP7_75t_L g13812 ( 
.A(n_13602),
.Y(n_13812)
);

OAI21x1_ASAP7_75t_L g13813 ( 
.A1(n_13499),
.A2(n_13476),
.B(n_13474),
.Y(n_13813)
);

AND2x4_ASAP7_75t_L g13814 ( 
.A(n_13602),
.B(n_13225),
.Y(n_13814)
);

INVx1_ASAP7_75t_SL g13815 ( 
.A(n_13528),
.Y(n_13815)
);

CKINVDCx16_ASAP7_75t_R g13816 ( 
.A(n_13551),
.Y(n_13816)
);

AND2x2_ASAP7_75t_L g13817 ( 
.A(n_13538),
.B(n_13448),
.Y(n_13817)
);

INVx2_ASAP7_75t_L g13818 ( 
.A(n_13618),
.Y(n_13818)
);

NAND2xp5_ASAP7_75t_L g13819 ( 
.A(n_13529),
.B(n_13197),
.Y(n_13819)
);

AOI22xp33_ASAP7_75t_SL g13820 ( 
.A1(n_13545),
.A2(n_13297),
.B1(n_13451),
.B2(n_13326),
.Y(n_13820)
);

NOR2xp33_ASAP7_75t_L g13821 ( 
.A(n_13604),
.B(n_13228),
.Y(n_13821)
);

INVxp67_ASAP7_75t_L g13822 ( 
.A(n_13582),
.Y(n_13822)
);

INVx1_ASAP7_75t_SL g13823 ( 
.A(n_13509),
.Y(n_13823)
);

AOI22xp5_ASAP7_75t_L g13824 ( 
.A1(n_13526),
.A2(n_13414),
.B1(n_13376),
.B2(n_13407),
.Y(n_13824)
);

OR2x2_ASAP7_75t_L g13825 ( 
.A(n_13524),
.B(n_13452),
.Y(n_13825)
);

INVx1_ASAP7_75t_L g13826 ( 
.A(n_13741),
.Y(n_13826)
);

INVx4_ASAP7_75t_L g13827 ( 
.A(n_13508),
.Y(n_13827)
);

AOI22xp33_ASAP7_75t_L g13828 ( 
.A1(n_13607),
.A2(n_13461),
.B1(n_13233),
.B2(n_13390),
.Y(n_13828)
);

INVx1_ASAP7_75t_SL g13829 ( 
.A(n_13495),
.Y(n_13829)
);

INVx2_ASAP7_75t_SL g13830 ( 
.A(n_13555),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_13668),
.Y(n_13831)
);

INVx1_ASAP7_75t_L g13832 ( 
.A(n_13550),
.Y(n_13832)
);

NAND2xp33_ASAP7_75t_SL g13833 ( 
.A(n_13782),
.B(n_13490),
.Y(n_13833)
);

AOI22xp33_ASAP7_75t_SL g13834 ( 
.A1(n_13533),
.A2(n_13264),
.B1(n_13205),
.B2(n_13480),
.Y(n_13834)
);

AND2x2_ASAP7_75t_L g13835 ( 
.A(n_13610),
.B(n_13366),
.Y(n_13835)
);

OAI22xp5_ASAP7_75t_L g13836 ( 
.A1(n_13558),
.A2(n_13243),
.B1(n_13426),
.B2(n_13352),
.Y(n_13836)
);

INVx2_ASAP7_75t_L g13837 ( 
.A(n_13511),
.Y(n_13837)
);

INVx1_ASAP7_75t_SL g13838 ( 
.A(n_13547),
.Y(n_13838)
);

CKINVDCx14_ASAP7_75t_R g13839 ( 
.A(n_13500),
.Y(n_13839)
);

NAND2xp5_ASAP7_75t_L g13840 ( 
.A(n_13554),
.B(n_13257),
.Y(n_13840)
);

INVx1_ASAP7_75t_L g13841 ( 
.A(n_13519),
.Y(n_13841)
);

NAND2xp5_ASAP7_75t_L g13842 ( 
.A(n_13502),
.B(n_13420),
.Y(n_13842)
);

INVx1_ASAP7_75t_SL g13843 ( 
.A(n_13540),
.Y(n_13843)
);

INVx1_ASAP7_75t_L g13844 ( 
.A(n_13651),
.Y(n_13844)
);

AND2x2_ASAP7_75t_L g13845 ( 
.A(n_13615),
.B(n_13496),
.Y(n_13845)
);

INVx1_ASAP7_75t_L g13846 ( 
.A(n_13593),
.Y(n_13846)
);

OR2x2_ASAP7_75t_L g13847 ( 
.A(n_13583),
.B(n_13621),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_13616),
.Y(n_13848)
);

INVx1_ASAP7_75t_L g13849 ( 
.A(n_13704),
.Y(n_13849)
);

AND2x2_ASAP7_75t_L g13850 ( 
.A(n_13535),
.B(n_13290),
.Y(n_13850)
);

INVx2_ASAP7_75t_L g13851 ( 
.A(n_13633),
.Y(n_13851)
);

INVx1_ASAP7_75t_L g13852 ( 
.A(n_13709),
.Y(n_13852)
);

INVx1_ASAP7_75t_L g13853 ( 
.A(n_13514),
.Y(n_13853)
);

INVx1_ASAP7_75t_SL g13854 ( 
.A(n_13566),
.Y(n_13854)
);

AOI21xp5_ASAP7_75t_L g13855 ( 
.A1(n_13521),
.A2(n_13277),
.B(n_13289),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_13552),
.B(n_13464),
.Y(n_13856)
);

AND2x2_ASAP7_75t_L g13857 ( 
.A(n_13594),
.B(n_13436),
.Y(n_13857)
);

INVx1_ASAP7_75t_L g13858 ( 
.A(n_13504),
.Y(n_13858)
);

NAND2xp5_ASAP7_75t_L g13859 ( 
.A(n_13619),
.B(n_13575),
.Y(n_13859)
);

INVx1_ASAP7_75t_L g13860 ( 
.A(n_13527),
.Y(n_13860)
);

INVx1_ASAP7_75t_SL g13861 ( 
.A(n_13649),
.Y(n_13861)
);

INVx2_ASAP7_75t_L g13862 ( 
.A(n_13522),
.Y(n_13862)
);

OR2x2_ASAP7_75t_L g13863 ( 
.A(n_13605),
.B(n_13437),
.Y(n_13863)
);

OR2x2_ASAP7_75t_L g13864 ( 
.A(n_13630),
.B(n_13463),
.Y(n_13864)
);

AND2x4_ASAP7_75t_SL g13865 ( 
.A(n_13608),
.B(n_7491),
.Y(n_13865)
);

INVx5_ASAP7_75t_L g13866 ( 
.A(n_13609),
.Y(n_13866)
);

OAI22xp5_ASAP7_75t_L g13867 ( 
.A1(n_13568),
.A2(n_13453),
.B1(n_13468),
.B2(n_13280),
.Y(n_13867)
);

AOI22xp33_ASAP7_75t_L g13868 ( 
.A1(n_13656),
.A2(n_13324),
.B1(n_13362),
.B2(n_13472),
.Y(n_13868)
);

INVx1_ASAP7_75t_SL g13869 ( 
.A(n_13678),
.Y(n_13869)
);

INVx1_ASAP7_75t_SL g13870 ( 
.A(n_13663),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_13647),
.Y(n_13871)
);

INVx1_ASAP7_75t_L g13872 ( 
.A(n_13756),
.Y(n_13872)
);

INVx1_ASAP7_75t_SL g13873 ( 
.A(n_13625),
.Y(n_13873)
);

INVx2_ASAP7_75t_L g13874 ( 
.A(n_13530),
.Y(n_13874)
);

INVx2_ASAP7_75t_L g13875 ( 
.A(n_13507),
.Y(n_13875)
);

BUFx2_ASAP7_75t_L g13876 ( 
.A(n_13559),
.Y(n_13876)
);

INVx2_ASAP7_75t_L g13877 ( 
.A(n_13564),
.Y(n_13877)
);

BUFx3_ASAP7_75t_L g13878 ( 
.A(n_13714),
.Y(n_13878)
);

INVx1_ASAP7_75t_L g13879 ( 
.A(n_13665),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_13667),
.Y(n_13880)
);

AND2x2_ASAP7_75t_L g13881 ( 
.A(n_13556),
.B(n_13457),
.Y(n_13881)
);

HB1xp67_ASAP7_75t_L g13882 ( 
.A(n_13525),
.Y(n_13882)
);

INVx2_ASAP7_75t_L g13883 ( 
.A(n_13660),
.Y(n_13883)
);

INVx1_ASAP7_75t_L g13884 ( 
.A(n_13728),
.Y(n_13884)
);

NAND2xp5_ASAP7_75t_SL g13885 ( 
.A(n_13553),
.B(n_13323),
.Y(n_13885)
);

AND2x2_ASAP7_75t_L g13886 ( 
.A(n_13600),
.B(n_13565),
.Y(n_13886)
);

INVx2_ASAP7_75t_L g13887 ( 
.A(n_13660),
.Y(n_13887)
);

INVx1_ASAP7_75t_SL g13888 ( 
.A(n_13627),
.Y(n_13888)
);

INVx1_ASAP7_75t_L g13889 ( 
.A(n_13645),
.Y(n_13889)
);

INVx2_ASAP7_75t_L g13890 ( 
.A(n_13549),
.Y(n_13890)
);

BUFx3_ASAP7_75t_L g13891 ( 
.A(n_13563),
.Y(n_13891)
);

OAI22xp5_ASAP7_75t_L g13892 ( 
.A1(n_13569),
.A2(n_13493),
.B1(n_9644),
.B2(n_9653),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_13657),
.Y(n_13893)
);

INVx1_ASAP7_75t_L g13894 ( 
.A(n_13612),
.Y(n_13894)
);

INVx1_ASAP7_75t_L g13895 ( 
.A(n_13546),
.Y(n_13895)
);

NOR2xp33_ASAP7_75t_SL g13896 ( 
.A(n_13742),
.B(n_13312),
.Y(n_13896)
);

NAND2xp5_ASAP7_75t_L g13897 ( 
.A(n_13567),
.B(n_9643),
.Y(n_13897)
);

AND2x2_ASAP7_75t_L g13898 ( 
.A(n_13523),
.B(n_9644),
.Y(n_13898)
);

OR2x2_ASAP7_75t_L g13899 ( 
.A(n_13571),
.B(n_9653),
.Y(n_13899)
);

INVx2_ASAP7_75t_L g13900 ( 
.A(n_13577),
.Y(n_13900)
);

NOR2x1_ASAP7_75t_L g13901 ( 
.A(n_13762),
.B(n_9654),
.Y(n_13901)
);

NOR2xp33_ASAP7_75t_SL g13902 ( 
.A(n_13680),
.B(n_7491),
.Y(n_13902)
);

NAND2xp5_ASAP7_75t_L g13903 ( 
.A(n_13572),
.B(n_9654),
.Y(n_13903)
);

INVx1_ASAP7_75t_SL g13904 ( 
.A(n_13750),
.Y(n_13904)
);

AND2x4_ASAP7_75t_L g13905 ( 
.A(n_13776),
.B(n_9659),
.Y(n_13905)
);

INVxp67_ASAP7_75t_SL g13906 ( 
.A(n_13697),
.Y(n_13906)
);

INVx4_ASAP7_75t_L g13907 ( 
.A(n_13780),
.Y(n_13907)
);

HB1xp67_ASAP7_75t_L g13908 ( 
.A(n_13804),
.Y(n_13908)
);

INVx2_ASAP7_75t_SL g13909 ( 
.A(n_13676),
.Y(n_13909)
);

NAND2xp5_ASAP7_75t_L g13910 ( 
.A(n_13557),
.B(n_9659),
.Y(n_13910)
);

OR2x2_ASAP7_75t_L g13911 ( 
.A(n_13706),
.B(n_9667),
.Y(n_13911)
);

AND2x2_ASAP7_75t_L g13912 ( 
.A(n_13699),
.B(n_9667),
.Y(n_13912)
);

AOI21xp5_ASAP7_75t_L g13913 ( 
.A1(n_13536),
.A2(n_9675),
.B(n_9670),
.Y(n_13913)
);

NOR2xp33_ASAP7_75t_L g13914 ( 
.A(n_13622),
.B(n_13745),
.Y(n_13914)
);

INVx1_ASAP7_75t_SL g13915 ( 
.A(n_13755),
.Y(n_13915)
);

INVx2_ASAP7_75t_L g13916 ( 
.A(n_13585),
.Y(n_13916)
);

AOI22xp5_ASAP7_75t_L g13917 ( 
.A1(n_13806),
.A2(n_8456),
.B1(n_7115),
.B2(n_7148),
.Y(n_13917)
);

AND2x2_ASAP7_75t_L g13918 ( 
.A(n_13512),
.B(n_9670),
.Y(n_13918)
);

INVx1_ASAP7_75t_L g13919 ( 
.A(n_13715),
.Y(n_13919)
);

INVx1_ASAP7_75t_SL g13920 ( 
.A(n_13698),
.Y(n_13920)
);

AND2x2_ASAP7_75t_L g13921 ( 
.A(n_13779),
.B(n_9675),
.Y(n_13921)
);

AND2x2_ASAP7_75t_L g13922 ( 
.A(n_13579),
.B(n_9679),
.Y(n_13922)
);

OR2x2_ASAP7_75t_L g13923 ( 
.A(n_13726),
.B(n_9679),
.Y(n_13923)
);

INVx1_ASAP7_75t_SL g13924 ( 
.A(n_13584),
.Y(n_13924)
);

AND2x2_ASAP7_75t_L g13925 ( 
.A(n_13581),
.B(n_9695),
.Y(n_13925)
);

HB1xp67_ASAP7_75t_L g13926 ( 
.A(n_13757),
.Y(n_13926)
);

INVx1_ASAP7_75t_L g13927 ( 
.A(n_13758),
.Y(n_13927)
);

BUFx2_ASAP7_75t_L g13928 ( 
.A(n_13501),
.Y(n_13928)
);

AOI22x1_ASAP7_75t_L g13929 ( 
.A1(n_13590),
.A2(n_9695),
.B1(n_7383),
.B2(n_7436),
.Y(n_13929)
);

NAND2xp5_ASAP7_75t_L g13930 ( 
.A(n_13586),
.B(n_13591),
.Y(n_13930)
);

OAI21xp5_ASAP7_75t_L g13931 ( 
.A1(n_13644),
.A2(n_8167),
.B(n_8148),
.Y(n_13931)
);

INVx1_ASAP7_75t_SL g13932 ( 
.A(n_13544),
.Y(n_13932)
);

AOI221xp5_ASAP7_75t_L g13933 ( 
.A1(n_13781),
.A2(n_13765),
.B1(n_13510),
.B2(n_13719),
.C(n_13642),
.Y(n_13933)
);

NAND2xp5_ASAP7_75t_L g13934 ( 
.A(n_13596),
.B(n_8078),
.Y(n_13934)
);

AOI22xp5_ASAP7_75t_L g13935 ( 
.A1(n_13580),
.A2(n_8456),
.B1(n_7115),
.B2(n_7148),
.Y(n_13935)
);

INVxp67_ASAP7_75t_SL g13936 ( 
.A(n_13679),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_13732),
.Y(n_13937)
);

AND2x2_ASAP7_75t_SL g13938 ( 
.A(n_13506),
.B(n_13597),
.Y(n_13938)
);

INVx1_ASAP7_75t_L g13939 ( 
.A(n_13692),
.Y(n_13939)
);

BUFx2_ASAP7_75t_L g13940 ( 
.A(n_13769),
.Y(n_13940)
);

AND2x2_ASAP7_75t_L g13941 ( 
.A(n_13599),
.B(n_8775),
.Y(n_13941)
);

INVx1_ASAP7_75t_SL g13942 ( 
.A(n_13685),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_13517),
.B(n_8775),
.Y(n_13943)
);

HB1xp67_ASAP7_75t_L g13944 ( 
.A(n_13757),
.Y(n_13944)
);

INVx2_ASAP7_75t_L g13945 ( 
.A(n_13655),
.Y(n_13945)
);

CKINVDCx14_ASAP7_75t_R g13946 ( 
.A(n_13498),
.Y(n_13946)
);

OA21x2_ASAP7_75t_L g13947 ( 
.A1(n_13759),
.A2(n_8130),
.B(n_8123),
.Y(n_13947)
);

HB1xp67_ASAP7_75t_L g13948 ( 
.A(n_13648),
.Y(n_13948)
);

NOR2x1_ASAP7_75t_L g13949 ( 
.A(n_13761),
.B(n_7558),
.Y(n_13949)
);

INVx2_ASAP7_75t_SL g13950 ( 
.A(n_13675),
.Y(n_13950)
);

NOR2xp33_ASAP7_75t_L g13951 ( 
.A(n_13736),
.B(n_7558),
.Y(n_13951)
);

NAND2xp5_ASAP7_75t_L g13952 ( 
.A(n_13763),
.B(n_8078),
.Y(n_13952)
);

INVx2_ASAP7_75t_L g13953 ( 
.A(n_13738),
.Y(n_13953)
);

OR2x2_ASAP7_75t_L g13954 ( 
.A(n_13634),
.B(n_13670),
.Y(n_13954)
);

HB1xp67_ASAP7_75t_L g13955 ( 
.A(n_13718),
.Y(n_13955)
);

INVx1_ASAP7_75t_L g13956 ( 
.A(n_13731),
.Y(n_13956)
);

INVx1_ASAP7_75t_SL g13957 ( 
.A(n_13696),
.Y(n_13957)
);

AND2x2_ASAP7_75t_L g13958 ( 
.A(n_13576),
.B(n_8775),
.Y(n_13958)
);

OR2x2_ASAP7_75t_L g13959 ( 
.A(n_13592),
.B(n_8079),
.Y(n_13959)
);

AOI22xp33_ASAP7_75t_L g13960 ( 
.A1(n_13631),
.A2(n_7559),
.B1(n_7560),
.B2(n_7558),
.Y(n_13960)
);

INVx1_ASAP7_75t_L g13961 ( 
.A(n_13734),
.Y(n_13961)
);

INVx1_ASAP7_75t_L g13962 ( 
.A(n_13774),
.Y(n_13962)
);

OR2x2_ASAP7_75t_L g13963 ( 
.A(n_13617),
.B(n_8079),
.Y(n_13963)
);

AND2x4_ASAP7_75t_L g13964 ( 
.A(n_13767),
.B(n_7558),
.Y(n_13964)
);

INVx1_ASAP7_75t_L g13965 ( 
.A(n_13661),
.Y(n_13965)
);

AOI22xp33_ASAP7_75t_L g13966 ( 
.A1(n_13623),
.A2(n_7560),
.B1(n_7564),
.B2(n_7559),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_13598),
.B(n_8456),
.Y(n_13967)
);

AND2x2_ASAP7_75t_L g13968 ( 
.A(n_13588),
.B(n_8456),
.Y(n_13968)
);

AND2x4_ASAP7_75t_L g13969 ( 
.A(n_13628),
.B(n_13764),
.Y(n_13969)
);

INVx1_ASAP7_75t_L g13970 ( 
.A(n_13534),
.Y(n_13970)
);

INVx1_ASAP7_75t_L g13971 ( 
.A(n_13548),
.Y(n_13971)
);

OR2x2_ASAP7_75t_L g13972 ( 
.A(n_13624),
.B(n_13766),
.Y(n_13972)
);

INVx2_ASAP7_75t_L g13973 ( 
.A(n_13751),
.Y(n_13973)
);

OR2x2_ASAP7_75t_L g13974 ( 
.A(n_13664),
.B(n_8082),
.Y(n_13974)
);

INVx3_ASAP7_75t_L g13975 ( 
.A(n_13659),
.Y(n_13975)
);

INVx1_ASAP7_75t_L g13976 ( 
.A(n_13561),
.Y(n_13976)
);

NAND2xp5_ASAP7_75t_L g13977 ( 
.A(n_13541),
.B(n_8082),
.Y(n_13977)
);

OR2x2_ASAP7_75t_L g13978 ( 
.A(n_13666),
.B(n_8086),
.Y(n_13978)
);

INVx1_ASAP7_75t_L g13979 ( 
.A(n_13520),
.Y(n_13979)
);

BUFx2_ASAP7_75t_L g13980 ( 
.A(n_13771),
.Y(n_13980)
);

AOI22xp33_ASAP7_75t_L g13981 ( 
.A1(n_13620),
.A2(n_7560),
.B1(n_7564),
.B2(n_7559),
.Y(n_13981)
);

BUFx2_ASAP7_75t_L g13982 ( 
.A(n_13775),
.Y(n_13982)
);

INVx2_ASAP7_75t_L g13983 ( 
.A(n_13532),
.Y(n_13983)
);

INVx1_ASAP7_75t_SL g13984 ( 
.A(n_13744),
.Y(n_13984)
);

INVx1_ASAP7_75t_SL g13985 ( 
.A(n_13695),
.Y(n_13985)
);

INVx1_ASAP7_75t_SL g13986 ( 
.A(n_13703),
.Y(n_13986)
);

INVx1_ASAP7_75t_L g13987 ( 
.A(n_13752),
.Y(n_13987)
);

NAND2xp5_ASAP7_75t_L g13988 ( 
.A(n_13650),
.B(n_13778),
.Y(n_13988)
);

INVx1_ASAP7_75t_L g13989 ( 
.A(n_13705),
.Y(n_13989)
);

HB1xp67_ASAP7_75t_L g13990 ( 
.A(n_13690),
.Y(n_13990)
);

OR2x2_ASAP7_75t_L g13991 ( 
.A(n_13669),
.B(n_8086),
.Y(n_13991)
);

AND2x2_ASAP7_75t_L g13992 ( 
.A(n_13796),
.B(n_8456),
.Y(n_13992)
);

CKINVDCx16_ASAP7_75t_R g13993 ( 
.A(n_13662),
.Y(n_13993)
);

NAND2xp5_ASAP7_75t_L g13994 ( 
.A(n_13754),
.B(n_8092),
.Y(n_13994)
);

NAND2xp5_ASAP7_75t_L g13995 ( 
.A(n_13613),
.B(n_13614),
.Y(n_13995)
);

AND2x2_ASAP7_75t_L g13996 ( 
.A(n_13636),
.B(n_8456),
.Y(n_13996)
);

INVx3_ASAP7_75t_SL g13997 ( 
.A(n_13589),
.Y(n_13997)
);

BUFx3_ASAP7_75t_L g13998 ( 
.A(n_13643),
.Y(n_13998)
);

OR2x2_ASAP7_75t_L g13999 ( 
.A(n_13733),
.B(n_8092),
.Y(n_13999)
);

INVx1_ASAP7_75t_L g14000 ( 
.A(n_13603),
.Y(n_14000)
);

AND2x2_ASAP7_75t_L g14001 ( 
.A(n_13646),
.B(n_8456),
.Y(n_14001)
);

NOR2x1_ASAP7_75t_L g14002 ( 
.A(n_13693),
.B(n_7559),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13626),
.Y(n_14003)
);

INVx1_ASAP7_75t_L g14004 ( 
.A(n_13717),
.Y(n_14004)
);

INVxp67_ASAP7_75t_L g14005 ( 
.A(n_13722),
.Y(n_14005)
);

INVx1_ASAP7_75t_SL g14006 ( 
.A(n_13689),
.Y(n_14006)
);

OR2x2_ASAP7_75t_L g14007 ( 
.A(n_13539),
.B(n_8093),
.Y(n_14007)
);

INVx1_ASAP7_75t_SL g14008 ( 
.A(n_13795),
.Y(n_14008)
);

OR2x2_ASAP7_75t_L g14009 ( 
.A(n_13789),
.B(n_8093),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_13773),
.Y(n_14010)
);

NAND2xp5_ASAP7_75t_L g14011 ( 
.A(n_13747),
.B(n_13711),
.Y(n_14011)
);

AOI222xp33_ASAP7_75t_L g14012 ( 
.A1(n_13652),
.A2(n_6146),
.B1(n_6032),
.B2(n_7115),
.C1(n_7148),
.C2(n_7030),
.Y(n_14012)
);

OR2x2_ASAP7_75t_L g14013 ( 
.A(n_13653),
.B(n_8098),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_13562),
.Y(n_14014)
);

CKINVDCx16_ASAP7_75t_R g14015 ( 
.A(n_13682),
.Y(n_14015)
);

NAND2xp5_ASAP7_75t_L g14016 ( 
.A(n_13790),
.B(n_8098),
.Y(n_14016)
);

INVx2_ASAP7_75t_L g14017 ( 
.A(n_13513),
.Y(n_14017)
);

HB1xp67_ASAP7_75t_L g14018 ( 
.A(n_13737),
.Y(n_14018)
);

INVx2_ASAP7_75t_L g14019 ( 
.A(n_13797),
.Y(n_14019)
);

INVx3_ASAP7_75t_L g14020 ( 
.A(n_13803),
.Y(n_14020)
);

INVx1_ASAP7_75t_L g14021 ( 
.A(n_13686),
.Y(n_14021)
);

INVx1_ASAP7_75t_SL g14022 ( 
.A(n_13505),
.Y(n_14022)
);

BUFx2_ASAP7_75t_L g14023 ( 
.A(n_13746),
.Y(n_14023)
);

BUFx2_ASAP7_75t_L g14024 ( 
.A(n_13772),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_13729),
.Y(n_14025)
);

AOI22xp33_ASAP7_75t_L g14026 ( 
.A1(n_13639),
.A2(n_7564),
.B1(n_7572),
.B2(n_7560),
.Y(n_14026)
);

AND2x2_ASAP7_75t_L g14027 ( 
.A(n_13785),
.B(n_8456),
.Y(n_14027)
);

AND2x2_ASAP7_75t_L g14028 ( 
.A(n_13793),
.B(n_6944),
.Y(n_14028)
);

INVx2_ASAP7_75t_L g14029 ( 
.A(n_13805),
.Y(n_14029)
);

AND2x2_ASAP7_75t_L g14030 ( 
.A(n_13632),
.B(n_13637),
.Y(n_14030)
);

INVx3_ASAP7_75t_SL g14031 ( 
.A(n_13543),
.Y(n_14031)
);

INVx1_ASAP7_75t_SL g14032 ( 
.A(n_13516),
.Y(n_14032)
);

NAND2xp5_ASAP7_75t_SL g14033 ( 
.A(n_13707),
.B(n_7030),
.Y(n_14033)
);

AND2x2_ASAP7_75t_L g14034 ( 
.A(n_13638),
.B(n_7402),
.Y(n_14034)
);

NOR2xp33_ASAP7_75t_L g14035 ( 
.A(n_13672),
.B(n_7564),
.Y(n_14035)
);

AND2x2_ASAP7_75t_L g14036 ( 
.A(n_13606),
.B(n_7402),
.Y(n_14036)
);

OR2x2_ASAP7_75t_L g14037 ( 
.A(n_13674),
.B(n_8100),
.Y(n_14037)
);

INVx1_ASAP7_75t_L g14038 ( 
.A(n_13735),
.Y(n_14038)
);

INVx4_ASAP7_75t_L g14039 ( 
.A(n_13694),
.Y(n_14039)
);

INVx2_ASAP7_75t_L g14040 ( 
.A(n_13658),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_13673),
.Y(n_14041)
);

NOR2x1_ASAP7_75t_L g14042 ( 
.A(n_13701),
.B(n_7572),
.Y(n_14042)
);

OAI21x1_ASAP7_75t_L g14043 ( 
.A1(n_13770),
.A2(n_8132),
.B(n_8130),
.Y(n_14043)
);

INVx2_ASAP7_75t_L g14044 ( 
.A(n_13684),
.Y(n_14044)
);

INVx1_ASAP7_75t_L g14045 ( 
.A(n_13713),
.Y(n_14045)
);

INVx1_ASAP7_75t_SL g14046 ( 
.A(n_13749),
.Y(n_14046)
);

INVx1_ASAP7_75t_L g14047 ( 
.A(n_13743),
.Y(n_14047)
);

INVx1_ASAP7_75t_L g14048 ( 
.A(n_13712),
.Y(n_14048)
);

AND2x2_ASAP7_75t_L g14049 ( 
.A(n_13681),
.B(n_7449),
.Y(n_14049)
);

HB1xp67_ASAP7_75t_L g14050 ( 
.A(n_13641),
.Y(n_14050)
);

AND2x2_ASAP7_75t_L g14051 ( 
.A(n_13683),
.B(n_7449),
.Y(n_14051)
);

INVx1_ASAP7_75t_L g14052 ( 
.A(n_13784),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13688),
.B(n_7455),
.Y(n_14053)
);

OR2x2_ASAP7_75t_L g14054 ( 
.A(n_13768),
.B(n_8100),
.Y(n_14054)
);

NAND2xp5_ASAP7_75t_L g14055 ( 
.A(n_13702),
.B(n_8102),
.Y(n_14055)
);

CKINVDCx16_ASAP7_75t_R g14056 ( 
.A(n_13798),
.Y(n_14056)
);

INVx1_ASAP7_75t_L g14057 ( 
.A(n_13708),
.Y(n_14057)
);

NAND2xp5_ASAP7_75t_L g14058 ( 
.A(n_13710),
.B(n_8102),
.Y(n_14058)
);

INVx2_ASAP7_75t_SL g14059 ( 
.A(n_13727),
.Y(n_14059)
);

INVx1_ASAP7_75t_L g14060 ( 
.A(n_13720),
.Y(n_14060)
);

AND2x2_ASAP7_75t_L g14061 ( 
.A(n_13723),
.B(n_7455),
.Y(n_14061)
);

BUFx3_ASAP7_75t_L g14062 ( 
.A(n_13783),
.Y(n_14062)
);

OR2x2_ASAP7_75t_L g14063 ( 
.A(n_13570),
.B(n_8114),
.Y(n_14063)
);

INVx2_ASAP7_75t_L g14064 ( 
.A(n_13748),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_L g14065 ( 
.A(n_13791),
.B(n_8114),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13794),
.B(n_7086),
.Y(n_14066)
);

A2O1A1Ixp33_ASAP7_75t_SL g14067 ( 
.A1(n_13801),
.A2(n_7120),
.B(n_7184),
.C(n_7087),
.Y(n_14067)
);

INVx1_ASAP7_75t_SL g14068 ( 
.A(n_13786),
.Y(n_14068)
);

NAND2xp5_ASAP7_75t_L g14069 ( 
.A(n_13792),
.B(n_8115),
.Y(n_14069)
);

NAND2xp5_ASAP7_75t_L g14070 ( 
.A(n_13802),
.B(n_8115),
.Y(n_14070)
);

HB1xp67_ASAP7_75t_L g14071 ( 
.A(n_13542),
.Y(n_14071)
);

BUFx3_ASAP7_75t_L g14072 ( 
.A(n_13777),
.Y(n_14072)
);

INVx1_ASAP7_75t_L g14073 ( 
.A(n_13753),
.Y(n_14073)
);

CKINVDCx16_ASAP7_75t_R g14074 ( 
.A(n_13799),
.Y(n_14074)
);

AND2x2_ASAP7_75t_L g14075 ( 
.A(n_13573),
.B(n_7120),
.Y(n_14075)
);

AND2x2_ASAP7_75t_L g14076 ( 
.A(n_13788),
.B(n_7184),
.Y(n_14076)
);

INVx1_ASAP7_75t_L g14077 ( 
.A(n_13760),
.Y(n_14077)
);

AND2x2_ASAP7_75t_L g14078 ( 
.A(n_13654),
.B(n_7184),
.Y(n_14078)
);

INVx1_ASAP7_75t_SL g14079 ( 
.A(n_13739),
.Y(n_14079)
);

INVx1_ASAP7_75t_L g14080 ( 
.A(n_13787),
.Y(n_14080)
);

INVx1_ASAP7_75t_L g14081 ( 
.A(n_13515),
.Y(n_14081)
);

INVx1_ASAP7_75t_L g14082 ( 
.A(n_13560),
.Y(n_14082)
);

INVx1_ASAP7_75t_SL g14083 ( 
.A(n_13629),
.Y(n_14083)
);

INVx1_ASAP7_75t_L g14084 ( 
.A(n_13601),
.Y(n_14084)
);

INVx1_ASAP7_75t_L g14085 ( 
.A(n_13611),
.Y(n_14085)
);

INVx1_ASAP7_75t_SL g14086 ( 
.A(n_13721),
.Y(n_14086)
);

NOR2x1_ASAP7_75t_L g14087 ( 
.A(n_13730),
.B(n_7572),
.Y(n_14087)
);

AND2x2_ASAP7_75t_L g14088 ( 
.A(n_13671),
.B(n_8130),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13677),
.Y(n_14089)
);

OR2x2_ASAP7_75t_L g14090 ( 
.A(n_13700),
.B(n_8121),
.Y(n_14090)
);

INVx1_ASAP7_75t_SL g14091 ( 
.A(n_13578),
.Y(n_14091)
);

HB1xp67_ASAP7_75t_L g14092 ( 
.A(n_13531),
.Y(n_14092)
);

AOI222xp33_ASAP7_75t_L g14093 ( 
.A1(n_13725),
.A2(n_6146),
.B1(n_6032),
.B2(n_7148),
.C1(n_7444),
.C2(n_7115),
.Y(n_14093)
);

INVx1_ASAP7_75t_SL g14094 ( 
.A(n_13635),
.Y(n_14094)
);

NAND2xp5_ASAP7_75t_L g14095 ( 
.A(n_13687),
.B(n_8121),
.Y(n_14095)
);

BUFx2_ASAP7_75t_L g14096 ( 
.A(n_13724),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_13691),
.Y(n_14097)
);

INVx1_ASAP7_75t_SL g14098 ( 
.A(n_13716),
.Y(n_14098)
);

INVx1_ASAP7_75t_SL g14099 ( 
.A(n_13640),
.Y(n_14099)
);

INVxp67_ASAP7_75t_L g14100 ( 
.A(n_13740),
.Y(n_14100)
);

OR2x2_ASAP7_75t_L g14101 ( 
.A(n_13800),
.B(n_8122),
.Y(n_14101)
);

INVx1_ASAP7_75t_L g14102 ( 
.A(n_13812),
.Y(n_14102)
);

AND2x2_ASAP7_75t_L g14103 ( 
.A(n_13816),
.B(n_8132),
.Y(n_14103)
);

AOI22xp5_ASAP7_75t_L g14104 ( 
.A1(n_13839),
.A2(n_7444),
.B1(n_7529),
.B2(n_7148),
.Y(n_14104)
);

INVx1_ASAP7_75t_SL g14105 ( 
.A(n_13811),
.Y(n_14105)
);

INVx1_ASAP7_75t_L g14106 ( 
.A(n_14018),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_SL g14107 ( 
.A(n_13866),
.B(n_7148),
.Y(n_14107)
);

NAND2xp5_ASAP7_75t_L g14108 ( 
.A(n_13858),
.B(n_8132),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_14092),
.Y(n_14109)
);

OAI221xp5_ASAP7_75t_SL g14110 ( 
.A1(n_13828),
.A2(n_7331),
.B1(n_7646),
.B2(n_7671),
.C(n_7621),
.Y(n_14110)
);

OAI32xp33_ASAP7_75t_SL g14111 ( 
.A1(n_13834),
.A2(n_9224),
.A3(n_9371),
.B1(n_9467),
.B2(n_9317),
.Y(n_14111)
);

OAI22xp33_ASAP7_75t_L g14112 ( 
.A1(n_14056),
.A2(n_7489),
.B1(n_7577),
.B2(n_7459),
.Y(n_14112)
);

OR2x2_ASAP7_75t_L g14113 ( 
.A(n_13907),
.B(n_8122),
.Y(n_14113)
);

NAND2xp5_ASAP7_75t_L g14114 ( 
.A(n_14022),
.B(n_8143),
.Y(n_14114)
);

INVxp67_ASAP7_75t_L g14115 ( 
.A(n_13833),
.Y(n_14115)
);

OAI21xp33_ASAP7_75t_L g14116 ( 
.A1(n_13902),
.A2(n_7444),
.B(n_7148),
.Y(n_14116)
);

NAND2xp5_ASAP7_75t_L g14117 ( 
.A(n_13866),
.B(n_13826),
.Y(n_14117)
);

NOR2xp33_ASAP7_75t_L g14118 ( 
.A(n_13907),
.B(n_7572),
.Y(n_14118)
);

OAI31xp33_ASAP7_75t_L g14119 ( 
.A1(n_13876),
.A2(n_6837),
.A3(n_6746),
.B(n_6817),
.Y(n_14119)
);

INVx1_ASAP7_75t_L g14120 ( 
.A(n_13845),
.Y(n_14120)
);

INVx1_ASAP7_75t_L g14121 ( 
.A(n_13906),
.Y(n_14121)
);

INVx1_ASAP7_75t_L g14122 ( 
.A(n_13866),
.Y(n_14122)
);

NAND3xp33_ASAP7_75t_L g14123 ( 
.A(n_13933),
.B(n_7529),
.C(n_7444),
.Y(n_14123)
);

INVxp67_ASAP7_75t_L g14124 ( 
.A(n_13821),
.Y(n_14124)
);

INVxp67_ASAP7_75t_L g14125 ( 
.A(n_13896),
.Y(n_14125)
);

OAI21xp33_ASAP7_75t_L g14126 ( 
.A1(n_13807),
.A2(n_7529),
.B(n_7444),
.Y(n_14126)
);

OAI22xp33_ASAP7_75t_L g14127 ( 
.A1(n_14031),
.A2(n_7459),
.B1(n_7577),
.B2(n_7489),
.Y(n_14127)
);

AOI21xp33_ASAP7_75t_SL g14128 ( 
.A1(n_13997),
.A2(n_9224),
.B(n_8214),
.Y(n_14128)
);

NAND2xp5_ASAP7_75t_L g14129 ( 
.A(n_13829),
.B(n_8143),
.Y(n_14129)
);

INVx1_ASAP7_75t_L g14130 ( 
.A(n_14071),
.Y(n_14130)
);

OR2x2_ASAP7_75t_L g14131 ( 
.A(n_13815),
.B(n_8125),
.Y(n_14131)
);

NOR2xp33_ASAP7_75t_L g14132 ( 
.A(n_13838),
.B(n_7645),
.Y(n_14132)
);

OAI21xp5_ASAP7_75t_L g14133 ( 
.A1(n_13855),
.A2(n_8214),
.B(n_8206),
.Y(n_14133)
);

INVx1_ASAP7_75t_L g14134 ( 
.A(n_14023),
.Y(n_14134)
);

INVx1_ASAP7_75t_L g14135 ( 
.A(n_13894),
.Y(n_14135)
);

OAI22xp33_ASAP7_75t_L g14136 ( 
.A1(n_14074),
.A2(n_14032),
.B1(n_13843),
.B2(n_13942),
.Y(n_14136)
);

NAND2xp5_ASAP7_75t_L g14137 ( 
.A(n_13808),
.B(n_8143),
.Y(n_14137)
);

HB1xp67_ASAP7_75t_L g14138 ( 
.A(n_13817),
.Y(n_14138)
);

AND2x2_ASAP7_75t_L g14139 ( 
.A(n_13846),
.B(n_8154),
.Y(n_14139)
);

INVx1_ASAP7_75t_L g14140 ( 
.A(n_14050),
.Y(n_14140)
);

NOR2xp33_ASAP7_75t_L g14141 ( 
.A(n_13854),
.B(n_7645),
.Y(n_14141)
);

INVx1_ASAP7_75t_L g14142 ( 
.A(n_13928),
.Y(n_14142)
);

OR2x2_ASAP7_75t_L g14143 ( 
.A(n_13859),
.B(n_8125),
.Y(n_14143)
);

AND2x2_ASAP7_75t_L g14144 ( 
.A(n_13871),
.B(n_8154),
.Y(n_14144)
);

OAI32xp33_ASAP7_75t_L g14145 ( 
.A1(n_14083),
.A2(n_7689),
.A3(n_7688),
.B1(n_7645),
.B2(n_8325),
.Y(n_14145)
);

A2O1A1Ixp33_ASAP7_75t_SL g14146 ( 
.A1(n_13946),
.A2(n_6491),
.B(n_6564),
.C(n_8154),
.Y(n_14146)
);

AOI221xp5_ASAP7_75t_L g14147 ( 
.A1(n_13836),
.A2(n_7534),
.B1(n_7576),
.B2(n_7529),
.C(n_7444),
.Y(n_14147)
);

AOI33xp33_ASAP7_75t_L g14148 ( 
.A1(n_13820),
.A2(n_7730),
.A3(n_7718),
.B1(n_7724),
.B2(n_7702),
.B3(n_6817),
.Y(n_14148)
);

INVxp67_ASAP7_75t_L g14149 ( 
.A(n_13980),
.Y(n_14149)
);

NAND3xp33_ASAP7_75t_L g14150 ( 
.A(n_13831),
.B(n_7529),
.C(n_7444),
.Y(n_14150)
);

A2O1A1Ixp33_ASAP7_75t_L g14151 ( 
.A1(n_13879),
.A2(n_8214),
.B(n_7759),
.C(n_7589),
.Y(n_14151)
);

OAI22xp33_ASAP7_75t_L g14152 ( 
.A1(n_13873),
.A2(n_7534),
.B1(n_7576),
.B2(n_7529),
.Y(n_14152)
);

A2O1A1Ixp33_ASAP7_75t_L g14153 ( 
.A1(n_13939),
.A2(n_7759),
.B(n_7589),
.C(n_6696),
.Y(n_14153)
);

INVx1_ASAP7_75t_L g14154 ( 
.A(n_13982),
.Y(n_14154)
);

XOR2x2_ASAP7_75t_L g14155 ( 
.A(n_14025),
.B(n_7433),
.Y(n_14155)
);

INVx5_ASAP7_75t_L g14156 ( 
.A(n_13827),
.Y(n_14156)
);

INVx1_ASAP7_75t_L g14157 ( 
.A(n_13936),
.Y(n_14157)
);

NOR4xp25_ASAP7_75t_SL g14158 ( 
.A(n_14096),
.B(n_8128),
.C(n_8134),
.D(n_8133),
.Y(n_14158)
);

OAI31xp33_ASAP7_75t_L g14159 ( 
.A1(n_13888),
.A2(n_6837),
.A3(n_6746),
.B(n_6696),
.Y(n_14159)
);

OAI31xp33_ASAP7_75t_L g14160 ( 
.A1(n_13861),
.A2(n_13915),
.A3(n_13904),
.B(n_13920),
.Y(n_14160)
);

AOI21xp33_ASAP7_75t_L g14161 ( 
.A1(n_13847),
.A2(n_9224),
.B(n_7383),
.Y(n_14161)
);

OAI211xp5_ASAP7_75t_L g14162 ( 
.A1(n_13809),
.A2(n_7688),
.B(n_7689),
.C(n_7645),
.Y(n_14162)
);

NAND3xp33_ASAP7_75t_L g14163 ( 
.A(n_13832),
.B(n_7534),
.C(n_7529),
.Y(n_14163)
);

AOI22xp33_ASAP7_75t_SL g14164 ( 
.A1(n_13940),
.A2(n_7574),
.B1(n_7615),
.B2(n_7497),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_13883),
.Y(n_14165)
);

A2O1A1Ixp33_ASAP7_75t_SL g14166 ( 
.A1(n_13914),
.A2(n_6491),
.B(n_6564),
.C(n_8155),
.Y(n_14166)
);

NAND3xp33_ASAP7_75t_L g14167 ( 
.A(n_13844),
.B(n_7576),
.C(n_7534),
.Y(n_14167)
);

INVx1_ASAP7_75t_L g14168 ( 
.A(n_13887),
.Y(n_14168)
);

NAND2x1_ASAP7_75t_L g14169 ( 
.A(n_13905),
.B(n_6726),
.Y(n_14169)
);

OAI21xp33_ASAP7_75t_L g14170 ( 
.A1(n_13835),
.A2(n_7576),
.B(n_7534),
.Y(n_14170)
);

OAI32xp33_ASAP7_75t_L g14171 ( 
.A1(n_13924),
.A2(n_7688),
.A3(n_7689),
.B1(n_8328),
.B2(n_8325),
.Y(n_14171)
);

NAND2xp5_ASAP7_75t_L g14172 ( 
.A(n_13969),
.B(n_8155),
.Y(n_14172)
);

HB1xp67_ASAP7_75t_L g14173 ( 
.A(n_13814),
.Y(n_14173)
);

INVxp67_ASAP7_75t_L g14174 ( 
.A(n_13849),
.Y(n_14174)
);

XNOR2x1_ASAP7_75t_L g14175 ( 
.A(n_13932),
.B(n_7615),
.Y(n_14175)
);

INVx1_ASAP7_75t_L g14176 ( 
.A(n_13852),
.Y(n_14176)
);

OAI21xp33_ASAP7_75t_L g14177 ( 
.A1(n_13842),
.A2(n_7576),
.B(n_7534),
.Y(n_14177)
);

INVx1_ASAP7_75t_L g14178 ( 
.A(n_13969),
.Y(n_14178)
);

INVx1_ASAP7_75t_L g14179 ( 
.A(n_13848),
.Y(n_14179)
);

AOI211xp5_ASAP7_75t_SL g14180 ( 
.A1(n_14005),
.A2(n_7780),
.B(n_6302),
.C(n_6449),
.Y(n_14180)
);

NAND3xp33_ASAP7_75t_SL g14181 ( 
.A(n_13823),
.B(n_5896),
.C(n_7688),
.Y(n_14181)
);

NOR3xp33_ASAP7_75t_L g14182 ( 
.A(n_13993),
.B(n_7689),
.C(n_6231),
.Y(n_14182)
);

INVx1_ASAP7_75t_L g14183 ( 
.A(n_13837),
.Y(n_14183)
);

INVx1_ASAP7_75t_L g14184 ( 
.A(n_13827),
.Y(n_14184)
);

NAND2xp5_ASAP7_75t_L g14185 ( 
.A(n_13880),
.B(n_14029),
.Y(n_14185)
);

OAI21xp5_ASAP7_75t_L g14186 ( 
.A1(n_13822),
.A2(n_8313),
.B(n_8223),
.Y(n_14186)
);

AND2x4_ASAP7_75t_L g14187 ( 
.A(n_13878),
.B(n_8155),
.Y(n_14187)
);

INVx1_ASAP7_75t_L g14188 ( 
.A(n_13891),
.Y(n_14188)
);

NOR2x1_ASAP7_75t_L g14189 ( 
.A(n_13818),
.B(n_8156),
.Y(n_14189)
);

OAI21xp33_ASAP7_75t_L g14190 ( 
.A1(n_13868),
.A2(n_7576),
.B(n_7534),
.Y(n_14190)
);

AND2x2_ASAP7_75t_L g14191 ( 
.A(n_14028),
.B(n_8156),
.Y(n_14191)
);

NAND2xp5_ASAP7_75t_L g14192 ( 
.A(n_14010),
.B(n_8156),
.Y(n_14192)
);

INVx1_ASAP7_75t_L g14193 ( 
.A(n_14024),
.Y(n_14193)
);

INVx1_ASAP7_75t_SL g14194 ( 
.A(n_13814),
.Y(n_14194)
);

A2O1A1Ixp33_ASAP7_75t_L g14195 ( 
.A1(n_13900),
.A2(n_7759),
.B(n_7589),
.C(n_6746),
.Y(n_14195)
);

INVx2_ASAP7_75t_L g14196 ( 
.A(n_13972),
.Y(n_14196)
);

AOI221xp5_ASAP7_75t_L g14197 ( 
.A1(n_13810),
.A2(n_7661),
.B1(n_7691),
.B2(n_7655),
.C(n_7576),
.Y(n_14197)
);

OR2x2_ASAP7_75t_L g14198 ( 
.A(n_14068),
.B(n_8128),
.Y(n_14198)
);

OAI32xp33_ASAP7_75t_L g14199 ( 
.A1(n_14081),
.A2(n_8331),
.A3(n_8333),
.B1(n_8328),
.B2(n_8325),
.Y(n_14199)
);

AOI21xp33_ASAP7_75t_SL g14200 ( 
.A1(n_14015),
.A2(n_8313),
.B(n_8223),
.Y(n_14200)
);

CKINVDCx16_ASAP7_75t_R g14201 ( 
.A(n_13998),
.Y(n_14201)
);

INVx1_ASAP7_75t_L g14202 ( 
.A(n_14049),
.Y(n_14202)
);

NAND2xp5_ASAP7_75t_L g14203 ( 
.A(n_13889),
.B(n_8160),
.Y(n_14203)
);

AND2x2_ASAP7_75t_L g14204 ( 
.A(n_14034),
.B(n_8160),
.Y(n_14204)
);

INVxp67_ASAP7_75t_L g14205 ( 
.A(n_13850),
.Y(n_14205)
);

NAND3xp33_ASAP7_75t_L g14206 ( 
.A(n_13841),
.B(n_7661),
.C(n_7655),
.Y(n_14206)
);

OAI211xp5_ASAP7_75t_SL g14207 ( 
.A1(n_13872),
.A2(n_7330),
.B(n_7358),
.C(n_7298),
.Y(n_14207)
);

NOR2xp33_ASAP7_75t_L g14208 ( 
.A(n_14039),
.B(n_7375),
.Y(n_14208)
);

INVx2_ASAP7_75t_L g14209 ( 
.A(n_13938),
.Y(n_14209)
);

NAND2xp5_ASAP7_75t_SL g14210 ( 
.A(n_14017),
.B(n_7655),
.Y(n_14210)
);

INVx1_ASAP7_75t_L g14211 ( 
.A(n_14051),
.Y(n_14211)
);

INVx1_ASAP7_75t_L g14212 ( 
.A(n_14053),
.Y(n_14212)
);

NAND2xp5_ASAP7_75t_L g14213 ( 
.A(n_13893),
.B(n_8160),
.Y(n_14213)
);

INVxp33_ASAP7_75t_L g14214 ( 
.A(n_13926),
.Y(n_14214)
);

OAI32xp33_ASAP7_75t_L g14215 ( 
.A1(n_13970),
.A2(n_13875),
.A3(n_14084),
.B1(n_14082),
.B2(n_14098),
.Y(n_14215)
);

AOI222xp33_ASAP7_75t_L g14216 ( 
.A1(n_14086),
.A2(n_7661),
.B1(n_7691),
.B2(n_7655),
.C1(n_7185),
.C2(n_6882),
.Y(n_14216)
);

AOI221xp5_ASAP7_75t_L g14217 ( 
.A1(n_13867),
.A2(n_7691),
.B1(n_7661),
.B2(n_7655),
.C(n_6882),
.Y(n_14217)
);

OAI22xp5_ASAP7_75t_L g14218 ( 
.A1(n_13917),
.A2(n_6726),
.B1(n_6735),
.B2(n_6727),
.Y(n_14218)
);

OAI22xp5_ASAP7_75t_L g14219 ( 
.A1(n_13960),
.A2(n_6726),
.B1(n_6735),
.B2(n_6727),
.Y(n_14219)
);

INVx1_ASAP7_75t_SL g14220 ( 
.A(n_13865),
.Y(n_14220)
);

INVx1_ASAP7_75t_L g14221 ( 
.A(n_13901),
.Y(n_14221)
);

OAI221xp5_ASAP7_75t_L g14222 ( 
.A1(n_13824),
.A2(n_6735),
.B1(n_6760),
.B2(n_6727),
.C(n_6726),
.Y(n_14222)
);

OAI31xp33_ASAP7_75t_L g14223 ( 
.A1(n_13869),
.A2(n_6837),
.A3(n_6868),
.B(n_6865),
.Y(n_14223)
);

NAND2xp5_ASAP7_75t_L g14224 ( 
.A(n_13919),
.B(n_8161),
.Y(n_14224)
);

INVx1_ASAP7_75t_L g14225 ( 
.A(n_13954),
.Y(n_14225)
);

INVx1_ASAP7_75t_L g14226 ( 
.A(n_13927),
.Y(n_14226)
);

INVx1_ASAP7_75t_L g14227 ( 
.A(n_14066),
.Y(n_14227)
);

AOI22xp33_ASAP7_75t_L g14228 ( 
.A1(n_13973),
.A2(n_7436),
.B1(n_7442),
.B2(n_7383),
.Y(n_14228)
);

NAND2xp5_ASAP7_75t_SL g14229 ( 
.A(n_13964),
.B(n_7655),
.Y(n_14229)
);

AOI21xp5_ASAP7_75t_SL g14230 ( 
.A1(n_14059),
.A2(n_5500),
.B(n_7655),
.Y(n_14230)
);

OR2x2_ASAP7_75t_L g14231 ( 
.A(n_14064),
.B(n_8133),
.Y(n_14231)
);

OAI221xp5_ASAP7_75t_L g14232 ( 
.A1(n_13966),
.A2(n_6735),
.B1(n_6760),
.B2(n_6727),
.C(n_6726),
.Y(n_14232)
);

INVxp67_ASAP7_75t_L g14233 ( 
.A(n_13944),
.Y(n_14233)
);

INVx2_ASAP7_75t_L g14234 ( 
.A(n_13905),
.Y(n_14234)
);

INVx1_ASAP7_75t_L g14235 ( 
.A(n_13856),
.Y(n_14235)
);

INVx1_ASAP7_75t_L g14236 ( 
.A(n_13813),
.Y(n_14236)
);

NAND2x1_ASAP7_75t_L g14237 ( 
.A(n_13949),
.B(n_6727),
.Y(n_14237)
);

O2A1O1Ixp5_ASAP7_75t_L g14238 ( 
.A1(n_13885),
.A2(n_7759),
.B(n_7964),
.C(n_8161),
.Y(n_14238)
);

XOR2x2_ASAP7_75t_L g14239 ( 
.A(n_13825),
.B(n_7780),
.Y(n_14239)
);

OAI21xp5_ASAP7_75t_SL g14240 ( 
.A1(n_13935),
.A2(n_7691),
.B(n_7661),
.Y(n_14240)
);

AOI321xp33_ASAP7_75t_L g14241 ( 
.A1(n_13892),
.A2(n_7214),
.A3(n_7223),
.B1(n_5896),
.B2(n_7267),
.C(n_7258),
.Y(n_14241)
);

INVx1_ASAP7_75t_L g14242 ( 
.A(n_13884),
.Y(n_14242)
);

INVx1_ASAP7_75t_L g14243 ( 
.A(n_13895),
.Y(n_14243)
);

NAND2xp5_ASAP7_75t_L g14244 ( 
.A(n_14000),
.B(n_8161),
.Y(n_14244)
);

NAND2xp5_ASAP7_75t_L g14245 ( 
.A(n_14003),
.B(n_8164),
.Y(n_14245)
);

NOR4xp25_ASAP7_75t_L g14246 ( 
.A(n_13979),
.B(n_8140),
.C(n_8144),
.D(n_8134),
.Y(n_14246)
);

O2A1O1Ixp33_ASAP7_75t_L g14247 ( 
.A1(n_13908),
.A2(n_6865),
.B(n_7128),
.C(n_6868),
.Y(n_14247)
);

OR2x2_ASAP7_75t_L g14248 ( 
.A(n_14046),
.B(n_8140),
.Y(n_14248)
);

OAI22xp5_ASAP7_75t_L g14249 ( 
.A1(n_13981),
.A2(n_14026),
.B1(n_13870),
.B2(n_13962),
.Y(n_14249)
);

INVx1_ASAP7_75t_SL g14250 ( 
.A(n_13964),
.Y(n_14250)
);

NAND2xp5_ASAP7_75t_L g14251 ( 
.A(n_14036),
.B(n_8164),
.Y(n_14251)
);

OAI211xp5_ASAP7_75t_L g14252 ( 
.A1(n_13840),
.A2(n_7691),
.B(n_7661),
.C(n_6882),
.Y(n_14252)
);

NAND2xp33_ASAP7_75t_R g14253 ( 
.A(n_13857),
.B(n_7625),
.Y(n_14253)
);

INVx1_ASAP7_75t_L g14254 ( 
.A(n_13819),
.Y(n_14254)
);

INVx1_ASAP7_75t_L g14255 ( 
.A(n_13911),
.Y(n_14255)
);

INVx1_ASAP7_75t_L g14256 ( 
.A(n_13923),
.Y(n_14256)
);

A2O1A1Ixp33_ASAP7_75t_L g14257 ( 
.A1(n_14035),
.A2(n_6865),
.B(n_7128),
.C(n_6868),
.Y(n_14257)
);

NAND2xp5_ASAP7_75t_SL g14258 ( 
.A(n_13965),
.B(n_7661),
.Y(n_14258)
);

INVx2_ASAP7_75t_L g14259 ( 
.A(n_14062),
.Y(n_14259)
);

INVx2_ASAP7_75t_SL g14260 ( 
.A(n_14087),
.Y(n_14260)
);

AND2x2_ASAP7_75t_L g14261 ( 
.A(n_13886),
.B(n_14078),
.Y(n_14261)
);

OAI22xp5_ASAP7_75t_L g14262 ( 
.A1(n_13985),
.A2(n_6735),
.B1(n_6772),
.B2(n_6760),
.Y(n_14262)
);

NAND2xp5_ASAP7_75t_L g14263 ( 
.A(n_14038),
.B(n_13976),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_13853),
.Y(n_14264)
);

AOI22xp5_ASAP7_75t_L g14265 ( 
.A1(n_13909),
.A2(n_14006),
.B1(n_14008),
.B2(n_13986),
.Y(n_14265)
);

OAI21xp5_ASAP7_75t_SL g14266 ( 
.A1(n_13984),
.A2(n_7691),
.B(n_6882),
.Y(n_14266)
);

NAND2xp5_ASAP7_75t_L g14267 ( 
.A(n_14014),
.B(n_8164),
.Y(n_14267)
);

INVx1_ASAP7_75t_L g14268 ( 
.A(n_13899),
.Y(n_14268)
);

AOI22xp5_ASAP7_75t_L g14269 ( 
.A1(n_13830),
.A2(n_7691),
.B1(n_6882),
.B2(n_7168),
.Y(n_14269)
);

INVx1_ASAP7_75t_L g14270 ( 
.A(n_13921),
.Y(n_14270)
);

INVx1_ASAP7_75t_L g14271 ( 
.A(n_13898),
.Y(n_14271)
);

INVx1_ASAP7_75t_SL g14272 ( 
.A(n_13881),
.Y(n_14272)
);

AOI22xp33_ASAP7_75t_L g14273 ( 
.A1(n_13990),
.A2(n_7442),
.B1(n_7461),
.B2(n_7436),
.Y(n_14273)
);

NAND2xp5_ASAP7_75t_L g14274 ( 
.A(n_14004),
.B(n_8168),
.Y(n_14274)
);

INVx2_ASAP7_75t_L g14275 ( 
.A(n_13958),
.Y(n_14275)
);

AOI22xp5_ASAP7_75t_L g14276 ( 
.A1(n_13950),
.A2(n_6882),
.B1(n_7168),
.B2(n_6791),
.Y(n_14276)
);

INVx1_ASAP7_75t_L g14277 ( 
.A(n_13988),
.Y(n_14277)
);

NAND2xp5_ASAP7_75t_L g14278 ( 
.A(n_14041),
.B(n_8168),
.Y(n_14278)
);

OAI32xp33_ASAP7_75t_L g14279 ( 
.A1(n_13863),
.A2(n_8333),
.A3(n_8338),
.B1(n_8331),
.B2(n_8328),
.Y(n_14279)
);

INVx1_ASAP7_75t_L g14280 ( 
.A(n_14040),
.Y(n_14280)
);

OAI22xp33_ASAP7_75t_L g14281 ( 
.A1(n_14091),
.A2(n_7168),
.B1(n_7185),
.B2(n_6791),
.Y(n_14281)
);

INVx1_ASAP7_75t_L g14282 ( 
.A(n_14044),
.Y(n_14282)
);

INVx2_ASAP7_75t_L g14283 ( 
.A(n_13941),
.Y(n_14283)
);

INVxp67_ASAP7_75t_SL g14284 ( 
.A(n_14002),
.Y(n_14284)
);

NAND2xp5_ASAP7_75t_L g14285 ( 
.A(n_14045),
.B(n_8168),
.Y(n_14285)
);

INVx1_ASAP7_75t_L g14286 ( 
.A(n_13910),
.Y(n_14286)
);

AOI21xp33_ASAP7_75t_SL g14287 ( 
.A1(n_14047),
.A2(n_7228),
.B(n_7128),
.Y(n_14287)
);

AOI21xp5_ASAP7_75t_L g14288 ( 
.A1(n_14011),
.A2(n_8176),
.B(n_8172),
.Y(n_14288)
);

INVx2_ASAP7_75t_L g14289 ( 
.A(n_13947),
.Y(n_14289)
);

INVx2_ASAP7_75t_L g14290 ( 
.A(n_13947),
.Y(n_14290)
);

HB1xp67_ASAP7_75t_L g14291 ( 
.A(n_14042),
.Y(n_14291)
);

AOI22xp5_ASAP7_75t_L g14292 ( 
.A1(n_13957),
.A2(n_7168),
.B1(n_7185),
.B2(n_6791),
.Y(n_14292)
);

INVx1_ASAP7_75t_L g14293 ( 
.A(n_13930),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_13922),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_13925),
.Y(n_14295)
);

AND2x4_ASAP7_75t_L g14296 ( 
.A(n_13912),
.B(n_8172),
.Y(n_14296)
);

OAI32xp33_ASAP7_75t_L g14297 ( 
.A1(n_14048),
.A2(n_14052),
.A3(n_13864),
.B1(n_13995),
.B2(n_13937),
.Y(n_14297)
);

INVxp67_ASAP7_75t_L g14298 ( 
.A(n_13951),
.Y(n_14298)
);

OAI322xp33_ASAP7_75t_L g14299 ( 
.A1(n_14100),
.A2(n_7741),
.A3(n_7671),
.B1(n_7788),
.B2(n_7727),
.C1(n_7646),
.C2(n_7042),
.Y(n_14299)
);

INVx1_ASAP7_75t_L g14300 ( 
.A(n_13955),
.Y(n_14300)
);

NOR2xp33_ASAP7_75t_L g14301 ( 
.A(n_14079),
.B(n_13989),
.Y(n_14301)
);

OAI21xp33_ASAP7_75t_SL g14302 ( 
.A1(n_14033),
.A2(n_8176),
.B(n_8172),
.Y(n_14302)
);

AOI22xp5_ASAP7_75t_L g14303 ( 
.A1(n_13860),
.A2(n_7168),
.B1(n_7185),
.B2(n_6791),
.Y(n_14303)
);

INVx1_ASAP7_75t_L g14304 ( 
.A(n_14076),
.Y(n_14304)
);

NOR3xp33_ASAP7_75t_L g14305 ( 
.A(n_13882),
.B(n_6231),
.C(n_6230),
.Y(n_14305)
);

O2A1O1Ixp33_ASAP7_75t_L g14306 ( 
.A1(n_13948),
.A2(n_7228),
.B(n_7254),
.C(n_7247),
.Y(n_14306)
);

AOI22xp33_ASAP7_75t_L g14307 ( 
.A1(n_13975),
.A2(n_7461),
.B1(n_7575),
.B2(n_7442),
.Y(n_14307)
);

NOR2xp33_ASAP7_75t_L g14308 ( 
.A(n_14020),
.B(n_7461),
.Y(n_14308)
);

OAI32xp33_ASAP7_75t_L g14309 ( 
.A1(n_13977),
.A2(n_8338),
.A3(n_8340),
.B1(n_8333),
.B2(n_8331),
.Y(n_14309)
);

NAND2xp5_ASAP7_75t_L g14310 ( 
.A(n_14061),
.B(n_8176),
.Y(n_14310)
);

NAND2xp5_ASAP7_75t_SL g14311 ( 
.A(n_13943),
.B(n_6791),
.Y(n_14311)
);

INVx1_ASAP7_75t_L g14312 ( 
.A(n_13897),
.Y(n_14312)
);

XNOR2xp5_ASAP7_75t_L g14313 ( 
.A(n_13929),
.B(n_6533),
.Y(n_14313)
);

INVx1_ASAP7_75t_SL g14314 ( 
.A(n_13992),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_13903),
.Y(n_14315)
);

OAI32xp33_ASAP7_75t_L g14316 ( 
.A1(n_14094),
.A2(n_8345),
.A3(n_8350),
.B1(n_8340),
.B2(n_8338),
.Y(n_14316)
);

INVx1_ASAP7_75t_L g14317 ( 
.A(n_13918),
.Y(n_14317)
);

NAND2xp5_ASAP7_75t_L g14318 ( 
.A(n_14075),
.B(n_14057),
.Y(n_14318)
);

INVx1_ASAP7_75t_L g14319 ( 
.A(n_14060),
.Y(n_14319)
);

OAI322xp33_ASAP7_75t_L g14320 ( 
.A1(n_14099),
.A2(n_7741),
.A3(n_7788),
.B1(n_7727),
.B2(n_7042),
.C1(n_7019),
.C2(n_6958),
.Y(n_14320)
);

XNOR2x1_ASAP7_75t_L g14321 ( 
.A(n_13877),
.B(n_6533),
.Y(n_14321)
);

OAI22xp5_ASAP7_75t_L g14322 ( 
.A1(n_13874),
.A2(n_6760),
.B1(n_6793),
.B2(n_6772),
.Y(n_14322)
);

INVx2_ASAP7_75t_L g14323 ( 
.A(n_14043),
.Y(n_14323)
);

AOI322xp5_ASAP7_75t_L g14324 ( 
.A1(n_13956),
.A2(n_13987),
.A3(n_13961),
.B1(n_13916),
.B2(n_13945),
.C1(n_13890),
.C2(n_13851),
.Y(n_14324)
);

NAND2xp5_ASAP7_75t_L g14325 ( 
.A(n_14027),
.B(n_8182),
.Y(n_14325)
);

OR2x2_ASAP7_75t_L g14326 ( 
.A(n_13994),
.B(n_8144),
.Y(n_14326)
);

AOI22xp5_ASAP7_75t_SL g14327 ( 
.A1(n_14030),
.A2(n_7168),
.B1(n_7185),
.B2(n_6791),
.Y(n_14327)
);

O2A1O1Ixp33_ASAP7_75t_L g14328 ( 
.A1(n_13953),
.A2(n_7228),
.B(n_7254),
.C(n_7247),
.Y(n_14328)
);

AOI22xp5_ASAP7_75t_L g14329 ( 
.A1(n_13862),
.A2(n_7225),
.B1(n_7362),
.B2(n_7185),
.Y(n_14329)
);

NAND2xp5_ASAP7_75t_L g14330 ( 
.A(n_14088),
.B(n_8182),
.Y(n_14330)
);

AND2x2_ASAP7_75t_L g14331 ( 
.A(n_13967),
.B(n_13968),
.Y(n_14331)
);

INVx1_ASAP7_75t_L g14332 ( 
.A(n_13952),
.Y(n_14332)
);

NAND2xp5_ASAP7_75t_L g14333 ( 
.A(n_14085),
.B(n_8182),
.Y(n_14333)
);

OR4x1_ASAP7_75t_L g14334 ( 
.A(n_14089),
.B(n_7254),
.C(n_7263),
.D(n_7247),
.Y(n_14334)
);

OAI21xp5_ASAP7_75t_L g14335 ( 
.A1(n_13913),
.A2(n_7346),
.B(n_7263),
.Y(n_14335)
);

AND2x4_ASAP7_75t_L g14336 ( 
.A(n_14072),
.B(n_8183),
.Y(n_14336)
);

O2A1O1Ixp33_ASAP7_75t_L g14337 ( 
.A1(n_14019),
.A2(n_7263),
.B(n_7386),
.C(n_7346),
.Y(n_14337)
);

INVxp33_ASAP7_75t_L g14338 ( 
.A(n_13983),
.Y(n_14338)
);

NOR2x1_ASAP7_75t_R g14339 ( 
.A(n_14097),
.B(n_7575),
.Y(n_14339)
);

NAND2xp5_ASAP7_75t_L g14340 ( 
.A(n_14178),
.B(n_13996),
.Y(n_14340)
);

AOI321xp33_ASAP7_75t_SL g14341 ( 
.A1(n_14272),
.A2(n_13963),
.A3(n_14021),
.B1(n_13971),
.B2(n_13991),
.C(n_13978),
.Y(n_14341)
);

INVx2_ASAP7_75t_L g14342 ( 
.A(n_14156),
.Y(n_14342)
);

AOI222xp33_ASAP7_75t_L g14343 ( 
.A1(n_14115),
.A2(n_14001),
.B1(n_14080),
.B2(n_14077),
.C1(n_14073),
.C2(n_14095),
.Y(n_14343)
);

INVx1_ASAP7_75t_L g14344 ( 
.A(n_14156),
.Y(n_14344)
);

NAND2xp5_ASAP7_75t_L g14345 ( 
.A(n_14138),
.B(n_14016),
.Y(n_14345)
);

OR2x2_ASAP7_75t_L g14346 ( 
.A(n_14194),
.B(n_13999),
.Y(n_14346)
);

INVx1_ASAP7_75t_L g14347 ( 
.A(n_14156),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_14173),
.Y(n_14348)
);

NOR2xp33_ASAP7_75t_L g14349 ( 
.A(n_14207),
.B(n_14090),
.Y(n_14349)
);

INVx1_ASAP7_75t_L g14350 ( 
.A(n_14117),
.Y(n_14350)
);

INVx1_ASAP7_75t_L g14351 ( 
.A(n_14184),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_14122),
.Y(n_14352)
);

NAND2xp5_ASAP7_75t_SL g14353 ( 
.A(n_14136),
.B(n_14012),
.Y(n_14353)
);

A2O1A1Ixp33_ASAP7_75t_L g14354 ( 
.A1(n_14160),
.A2(n_14101),
.B(n_13934),
.C(n_14009),
.Y(n_14354)
);

OR2x2_ASAP7_75t_L g14355 ( 
.A(n_14130),
.B(n_14069),
.Y(n_14355)
);

AND2x4_ASAP7_75t_SL g14356 ( 
.A(n_14193),
.B(n_13974),
.Y(n_14356)
);

INVx1_ASAP7_75t_L g14357 ( 
.A(n_14142),
.Y(n_14357)
);

NOR2xp67_ASAP7_75t_L g14358 ( 
.A(n_14149),
.B(n_14013),
.Y(n_14358)
);

INVx2_ASAP7_75t_L g14359 ( 
.A(n_14155),
.Y(n_14359)
);

NAND2xp5_ASAP7_75t_L g14360 ( 
.A(n_14125),
.B(n_14070),
.Y(n_14360)
);

INVx1_ASAP7_75t_L g14361 ( 
.A(n_14154),
.Y(n_14361)
);

AND2x2_ASAP7_75t_L g14362 ( 
.A(n_14140),
.B(n_14205),
.Y(n_14362)
);

NOR3xp33_ASAP7_75t_L g14363 ( 
.A(n_14201),
.B(n_14058),
.C(n_14055),
.Y(n_14363)
);

AND2x2_ASAP7_75t_L g14364 ( 
.A(n_14105),
.B(n_14037),
.Y(n_14364)
);

INVx2_ASAP7_75t_L g14365 ( 
.A(n_14239),
.Y(n_14365)
);

INVx1_ASAP7_75t_L g14366 ( 
.A(n_14102),
.Y(n_14366)
);

INVx1_ASAP7_75t_L g14367 ( 
.A(n_14234),
.Y(n_14367)
);

OAI21xp5_ASAP7_75t_L g14368 ( 
.A1(n_14174),
.A2(n_14065),
.B(n_14054),
.Y(n_14368)
);

INVx1_ASAP7_75t_L g14369 ( 
.A(n_14185),
.Y(n_14369)
);

OAI21xp33_ASAP7_75t_SL g14370 ( 
.A1(n_14148),
.A2(n_14093),
.B(n_13959),
.Y(n_14370)
);

NAND2xp5_ASAP7_75t_L g14371 ( 
.A(n_14109),
.B(n_14007),
.Y(n_14371)
);

OAI22xp5_ASAP7_75t_L g14372 ( 
.A1(n_14228),
.A2(n_14063),
.B1(n_13931),
.B2(n_14067),
.Y(n_14372)
);

AND2x2_ASAP7_75t_L g14373 ( 
.A(n_14120),
.B(n_8340),
.Y(n_14373)
);

INVx1_ASAP7_75t_L g14374 ( 
.A(n_14289),
.Y(n_14374)
);

AOI211xp5_ASAP7_75t_L g14375 ( 
.A1(n_14215),
.A2(n_5500),
.B(n_7481),
.C(n_7362),
.Y(n_14375)
);

INVx2_ASAP7_75t_L g14376 ( 
.A(n_14175),
.Y(n_14376)
);

INVx1_ASAP7_75t_L g14377 ( 
.A(n_14290),
.Y(n_14377)
);

AND2x2_ASAP7_75t_L g14378 ( 
.A(n_14196),
.B(n_8795),
.Y(n_14378)
);

NOR3xp33_ASAP7_75t_L g14379 ( 
.A(n_14233),
.B(n_6231),
.C(n_6230),
.Y(n_14379)
);

AOI211xp5_ASAP7_75t_SL g14380 ( 
.A1(n_14249),
.A2(n_6302),
.B(n_6449),
.C(n_6366),
.Y(n_14380)
);

INVx1_ASAP7_75t_L g14381 ( 
.A(n_14134),
.Y(n_14381)
);

OAI21xp33_ASAP7_75t_L g14382 ( 
.A1(n_14190),
.A2(n_7362),
.B(n_7225),
.Y(n_14382)
);

NAND2xp5_ASAP7_75t_L g14383 ( 
.A(n_14202),
.B(n_8192),
.Y(n_14383)
);

INVx2_ASAP7_75t_L g14384 ( 
.A(n_14334),
.Y(n_14384)
);

INVx1_ASAP7_75t_L g14385 ( 
.A(n_14291),
.Y(n_14385)
);

OAI21xp5_ASAP7_75t_L g14386 ( 
.A1(n_14195),
.A2(n_7386),
.B(n_7346),
.Y(n_14386)
);

AOI21xp5_ASAP7_75t_L g14387 ( 
.A1(n_14263),
.A2(n_8188),
.B(n_8183),
.Y(n_14387)
);

INVx1_ASAP7_75t_L g14388 ( 
.A(n_14221),
.Y(n_14388)
);

NOR3xp33_ASAP7_75t_L g14389 ( 
.A(n_14209),
.B(n_6231),
.C(n_6230),
.Y(n_14389)
);

AOI22xp5_ASAP7_75t_L g14390 ( 
.A1(n_14253),
.A2(n_7590),
.B1(n_7667),
.B2(n_7575),
.Y(n_14390)
);

AOI21xp33_ASAP7_75t_SL g14391 ( 
.A1(n_14236),
.A2(n_9371),
.B(n_9317),
.Y(n_14391)
);

NAND2xp5_ASAP7_75t_L g14392 ( 
.A(n_14211),
.B(n_8195),
.Y(n_14392)
);

OAI21xp33_ASAP7_75t_SL g14393 ( 
.A1(n_14107),
.A2(n_8188),
.B(n_8183),
.Y(n_14393)
);

INVx1_ASAP7_75t_L g14394 ( 
.A(n_14103),
.Y(n_14394)
);

NAND2xp5_ASAP7_75t_L g14395 ( 
.A(n_14212),
.B(n_8318),
.Y(n_14395)
);

NAND3xp33_ASAP7_75t_SL g14396 ( 
.A(n_14250),
.B(n_14265),
.C(n_14220),
.Y(n_14396)
);

AND2x2_ASAP7_75t_L g14397 ( 
.A(n_14261),
.B(n_8805),
.Y(n_14397)
);

OR2x2_ASAP7_75t_L g14398 ( 
.A(n_14183),
.B(n_8188),
.Y(n_14398)
);

OAI22xp5_ASAP7_75t_L g14399 ( 
.A1(n_14307),
.A2(n_8192),
.B1(n_8195),
.B2(n_8189),
.Y(n_14399)
);

OAI21xp5_ASAP7_75t_L g14400 ( 
.A1(n_14153),
.A2(n_7420),
.B(n_7386),
.Y(n_14400)
);

NAND2xp5_ASAP7_75t_L g14401 ( 
.A(n_14176),
.B(n_8244),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_14114),
.Y(n_14402)
);

INVx2_ASAP7_75t_L g14403 ( 
.A(n_14237),
.Y(n_14403)
);

OAI21xp5_ASAP7_75t_L g14404 ( 
.A1(n_14214),
.A2(n_7506),
.B(n_7420),
.Y(n_14404)
);

INVx1_ASAP7_75t_L g14405 ( 
.A(n_14113),
.Y(n_14405)
);

INVxp33_ASAP7_75t_L g14406 ( 
.A(n_14132),
.Y(n_14406)
);

AOI22xp5_ASAP7_75t_L g14407 ( 
.A1(n_14262),
.A2(n_7667),
.B1(n_7699),
.B2(n_7590),
.Y(n_14407)
);

NAND2xp5_ASAP7_75t_L g14408 ( 
.A(n_14280),
.B(n_8244),
.Y(n_14408)
);

NAND2xp5_ASAP7_75t_L g14409 ( 
.A(n_14282),
.B(n_8244),
.Y(n_14409)
);

INVx1_ASAP7_75t_L g14410 ( 
.A(n_14284),
.Y(n_14410)
);

OAI21xp5_ASAP7_75t_L g14411 ( 
.A1(n_14123),
.A2(n_7506),
.B(n_7420),
.Y(n_14411)
);

AOI22xp5_ASAP7_75t_L g14412 ( 
.A1(n_14322),
.A2(n_7667),
.B1(n_7699),
.B2(n_7590),
.Y(n_14412)
);

INVx1_ASAP7_75t_L g14413 ( 
.A(n_14172),
.Y(n_14413)
);

OAI22xp33_ASAP7_75t_SL g14414 ( 
.A1(n_14169),
.A2(n_6976),
.B1(n_6992),
.B2(n_6955),
.Y(n_14414)
);

NAND2x1p5_ASAP7_75t_L g14415 ( 
.A(n_14225),
.B(n_14188),
.Y(n_14415)
);

NOR2xp33_ASAP7_75t_L g14416 ( 
.A(n_14112),
.B(n_7699),
.Y(n_14416)
);

AOI222xp33_ASAP7_75t_L g14417 ( 
.A1(n_14254),
.A2(n_7481),
.B1(n_7362),
.B2(n_7510),
.C1(n_7370),
.C2(n_7225),
.Y(n_14417)
);

INVx1_ASAP7_75t_L g14418 ( 
.A(n_14108),
.Y(n_14418)
);

OAI21xp5_ASAP7_75t_L g14419 ( 
.A1(n_14124),
.A2(n_7522),
.B(n_7506),
.Y(n_14419)
);

NAND2xp5_ASAP7_75t_L g14420 ( 
.A(n_14227),
.B(n_8195),
.Y(n_14420)
);

AOI322xp5_ASAP7_75t_L g14421 ( 
.A1(n_14170),
.A2(n_6958),
.A3(n_6973),
.B1(n_7061),
.B2(n_7073),
.C1(n_7019),
.C2(n_7011),
.Y(n_14421)
);

AND2x2_ASAP7_75t_L g14422 ( 
.A(n_14259),
.B(n_8795),
.Y(n_14422)
);

INVxp67_ASAP7_75t_L g14423 ( 
.A(n_14118),
.Y(n_14423)
);

OAI22xp5_ASAP7_75t_L g14424 ( 
.A1(n_14273),
.A2(n_8192),
.B1(n_8201),
.B2(n_8189),
.Y(n_14424)
);

INVx1_ASAP7_75t_L g14425 ( 
.A(n_14242),
.Y(n_14425)
);

AOI221xp5_ASAP7_75t_L g14426 ( 
.A1(n_14297),
.A2(n_7362),
.B1(n_7481),
.B2(n_7370),
.C(n_7225),
.Y(n_14426)
);

INVx1_ASAP7_75t_SL g14427 ( 
.A(n_14131),
.Y(n_14427)
);

AOI221xp5_ASAP7_75t_L g14428 ( 
.A1(n_14145),
.A2(n_7362),
.B1(n_7481),
.B2(n_7370),
.C(n_7225),
.Y(n_14428)
);

NOR2xp33_ASAP7_75t_L g14429 ( 
.A(n_14338),
.B(n_7736),
.Y(n_14429)
);

AOI21xp33_ASAP7_75t_L g14430 ( 
.A1(n_14339),
.A2(n_7736),
.B(n_7703),
.Y(n_14430)
);

NAND2xp5_ASAP7_75t_L g14431 ( 
.A(n_14165),
.B(n_8208),
.Y(n_14431)
);

NAND2xp5_ASAP7_75t_L g14432 ( 
.A(n_14168),
.B(n_8208),
.Y(n_14432)
);

INVx2_ASAP7_75t_SL g14433 ( 
.A(n_14248),
.Y(n_14433)
);

NAND3xp33_ASAP7_75t_SL g14434 ( 
.A(n_14106),
.B(n_7061),
.C(n_6973),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_14235),
.Y(n_14435)
);

NAND2xp5_ASAP7_75t_L g14436 ( 
.A(n_14135),
.B(n_8189),
.Y(n_14436)
);

OAI211xp5_ASAP7_75t_L g14437 ( 
.A1(n_14324),
.A2(n_14177),
.B(n_14230),
.C(n_14162),
.Y(n_14437)
);

OR2x2_ASAP7_75t_L g14438 ( 
.A(n_14179),
.B(n_8201),
.Y(n_14438)
);

INVx1_ASAP7_75t_L g14439 ( 
.A(n_14189),
.Y(n_14439)
);

INVx2_ASAP7_75t_L g14440 ( 
.A(n_14321),
.Y(n_14440)
);

OAI21xp33_ASAP7_75t_L g14441 ( 
.A1(n_14308),
.A2(n_7370),
.B(n_7225),
.Y(n_14441)
);

OAI21xp33_ASAP7_75t_SL g14442 ( 
.A1(n_14119),
.A2(n_8208),
.B(n_8201),
.Y(n_14442)
);

INVx1_ASAP7_75t_SL g14443 ( 
.A(n_14139),
.Y(n_14443)
);

AOI22xp5_ASAP7_75t_L g14444 ( 
.A1(n_14305),
.A2(n_7736),
.B1(n_7754),
.B2(n_7703),
.Y(n_14444)
);

INVx1_ASAP7_75t_SL g14445 ( 
.A(n_14144),
.Y(n_14445)
);

OAI221xp5_ASAP7_75t_L g14446 ( 
.A1(n_14166),
.A2(n_6793),
.B1(n_6815),
.B2(n_6772),
.C(n_6760),
.Y(n_14446)
);

AOI22xp33_ASAP7_75t_L g14447 ( 
.A1(n_14182),
.A2(n_7754),
.B1(n_7791),
.B2(n_7703),
.Y(n_14447)
);

NAND3xp33_ASAP7_75t_L g14448 ( 
.A(n_14121),
.B(n_7481),
.C(n_7370),
.Y(n_14448)
);

NAND4xp25_ASAP7_75t_L g14449 ( 
.A(n_14110),
.B(n_6606),
.C(n_6667),
.D(n_6533),
.Y(n_14449)
);

INVx1_ASAP7_75t_L g14450 ( 
.A(n_14323),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_14294),
.Y(n_14451)
);

INVx1_ASAP7_75t_L g14452 ( 
.A(n_14295),
.Y(n_14452)
);

INVx1_ASAP7_75t_L g14453 ( 
.A(n_14271),
.Y(n_14453)
);

NAND2xp5_ASAP7_75t_L g14454 ( 
.A(n_14317),
.B(n_8232),
.Y(n_14454)
);

INVx2_ASAP7_75t_L g14455 ( 
.A(n_14191),
.Y(n_14455)
);

AOI32xp33_ASAP7_75t_L g14456 ( 
.A1(n_14127),
.A2(n_7073),
.A3(n_7133),
.B1(n_7096),
.B2(n_7011),
.Y(n_14456)
);

INVxp67_ASAP7_75t_SL g14457 ( 
.A(n_14260),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_14129),
.Y(n_14458)
);

INVxp33_ASAP7_75t_L g14459 ( 
.A(n_14141),
.Y(n_14459)
);

NAND4xp25_ASAP7_75t_L g14460 ( 
.A(n_14222),
.B(n_6606),
.C(n_6667),
.D(n_6533),
.Y(n_14460)
);

INVx1_ASAP7_75t_L g14461 ( 
.A(n_14157),
.Y(n_14461)
);

O2A1O1Ixp33_ASAP7_75t_L g14462 ( 
.A1(n_14146),
.A2(n_7522),
.B(n_7767),
.C(n_7650),
.Y(n_14462)
);

INVx1_ASAP7_75t_L g14463 ( 
.A(n_14226),
.Y(n_14463)
);

NAND2xp5_ASAP7_75t_L g14464 ( 
.A(n_14270),
.B(n_14268),
.Y(n_14464)
);

OAI21xp33_ASAP7_75t_L g14465 ( 
.A1(n_14300),
.A2(n_7481),
.B(n_7370),
.Y(n_14465)
);

NAND2xp5_ASAP7_75t_L g14466 ( 
.A(n_14243),
.B(n_8264),
.Y(n_14466)
);

NAND2xp5_ASAP7_75t_L g14467 ( 
.A(n_14187),
.B(n_14336),
.Y(n_14467)
);

AND2x2_ASAP7_75t_L g14468 ( 
.A(n_14283),
.B(n_8795),
.Y(n_14468)
);

AOI221xp5_ASAP7_75t_L g14469 ( 
.A1(n_14287),
.A2(n_7711),
.B1(n_7714),
.B2(n_7510),
.C(n_7096),
.Y(n_14469)
);

AND2x2_ASAP7_75t_L g14470 ( 
.A(n_14275),
.B(n_8798),
.Y(n_14470)
);

AND2x2_ASAP7_75t_L g14471 ( 
.A(n_14304),
.B(n_8798),
.Y(n_14471)
);

OAI22xp33_ASAP7_75t_L g14472 ( 
.A1(n_14104),
.A2(n_7711),
.B1(n_7714),
.B2(n_7510),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_14318),
.Y(n_14473)
);

OR2x2_ASAP7_75t_L g14474 ( 
.A(n_14264),
.B(n_8215),
.Y(n_14474)
);

INVx1_ASAP7_75t_L g14475 ( 
.A(n_14198),
.Y(n_14475)
);

OA211x2_ASAP7_75t_L g14476 ( 
.A1(n_14208),
.A2(n_6366),
.B(n_6362),
.C(n_7101),
.Y(n_14476)
);

NAND2xp5_ASAP7_75t_L g14477 ( 
.A(n_14187),
.B(n_8232),
.Y(n_14477)
);

OAI221xp5_ASAP7_75t_SL g14478 ( 
.A1(n_14223),
.A2(n_7331),
.B1(n_7196),
.B2(n_7239),
.C(n_7163),
.Y(n_14478)
);

AOI22xp33_ASAP7_75t_SL g14479 ( 
.A1(n_14277),
.A2(n_14218),
.B1(n_14301),
.B2(n_14206),
.Y(n_14479)
);

OR2x2_ASAP7_75t_L g14480 ( 
.A(n_14255),
.B(n_8215),
.Y(n_14480)
);

NAND2xp5_ASAP7_75t_L g14481 ( 
.A(n_14336),
.B(n_14256),
.Y(n_14481)
);

INVx2_ASAP7_75t_SL g14482 ( 
.A(n_14258),
.Y(n_14482)
);

INVx1_ASAP7_75t_L g14483 ( 
.A(n_14231),
.Y(n_14483)
);

INVx2_ASAP7_75t_SL g14484 ( 
.A(n_14204),
.Y(n_14484)
);

INVx1_ASAP7_75t_L g14485 ( 
.A(n_14319),
.Y(n_14485)
);

AOI221xp5_ASAP7_75t_L g14486 ( 
.A1(n_14171),
.A2(n_14126),
.B1(n_14246),
.B2(n_14116),
.C(n_14167),
.Y(n_14486)
);

AOI22xp5_ASAP7_75t_L g14487 ( 
.A1(n_14219),
.A2(n_7791),
.B1(n_7754),
.B2(n_7711),
.Y(n_14487)
);

OAI22xp5_ASAP7_75t_L g14488 ( 
.A1(n_14276),
.A2(n_8220),
.B1(n_8232),
.B2(n_8215),
.Y(n_14488)
);

INVxp67_ASAP7_75t_SL g14489 ( 
.A(n_14210),
.Y(n_14489)
);

NAND2xp5_ASAP7_75t_L g14490 ( 
.A(n_14296),
.B(n_8283),
.Y(n_14490)
);

INVx2_ASAP7_75t_L g14491 ( 
.A(n_14238),
.Y(n_14491)
);

INVx1_ASAP7_75t_L g14492 ( 
.A(n_14137),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_14143),
.Y(n_14493)
);

CKINVDCx16_ASAP7_75t_R g14494 ( 
.A(n_14293),
.Y(n_14494)
);

INVx1_ASAP7_75t_L g14495 ( 
.A(n_14203),
.Y(n_14495)
);

NAND2xp5_ASAP7_75t_L g14496 ( 
.A(n_14296),
.B(n_8283),
.Y(n_14496)
);

OR2x2_ASAP7_75t_L g14497 ( 
.A(n_14310),
.B(n_8220),
.Y(n_14497)
);

OAI211xp5_ASAP7_75t_L g14498 ( 
.A1(n_14298),
.A2(n_7711),
.B(n_7714),
.C(n_7510),
.Y(n_14498)
);

NOR2xp33_ASAP7_75t_L g14499 ( 
.A(n_14314),
.B(n_7791),
.Y(n_14499)
);

NAND2xp5_ASAP7_75t_L g14500 ( 
.A(n_14331),
.B(n_8259),
.Y(n_14500)
);

INVx2_ASAP7_75t_L g14501 ( 
.A(n_14326),
.Y(n_14501)
);

INVxp67_ASAP7_75t_L g14502 ( 
.A(n_14213),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_14224),
.Y(n_14503)
);

NOR2xp33_ASAP7_75t_L g14504 ( 
.A(n_14286),
.B(n_6772),
.Y(n_14504)
);

INVx1_ASAP7_75t_L g14505 ( 
.A(n_14192),
.Y(n_14505)
);

OAI22xp5_ASAP7_75t_L g14506 ( 
.A1(n_14269),
.A2(n_8234),
.B1(n_8251),
.B2(n_8220),
.Y(n_14506)
);

INVx1_ASAP7_75t_L g14507 ( 
.A(n_14278),
.Y(n_14507)
);

AOI211xp5_ASAP7_75t_L g14508 ( 
.A1(n_14266),
.A2(n_7714),
.B(n_7711),
.C(n_7510),
.Y(n_14508)
);

AND2x2_ASAP7_75t_L g14509 ( 
.A(n_14313),
.B(n_8810),
.Y(n_14509)
);

CKINVDCx16_ASAP7_75t_R g14510 ( 
.A(n_14312),
.Y(n_14510)
);

NOR2xp33_ASAP7_75t_L g14511 ( 
.A(n_14315),
.B(n_6772),
.Y(n_14511)
);

INVx1_ASAP7_75t_L g14512 ( 
.A(n_14285),
.Y(n_14512)
);

NAND2xp5_ASAP7_75t_L g14513 ( 
.A(n_14332),
.B(n_8291),
.Y(n_14513)
);

NAND2xp5_ASAP7_75t_L g14514 ( 
.A(n_14158),
.B(n_8291),
.Y(n_14514)
);

OAI211xp5_ASAP7_75t_L g14515 ( 
.A1(n_14333),
.A2(n_7711),
.B(n_7714),
.C(n_7510),
.Y(n_14515)
);

AOI221x1_ASAP7_75t_L g14516 ( 
.A1(n_14163),
.A2(n_8158),
.B1(n_8174),
.B2(n_8169),
.C(n_8152),
.Y(n_14516)
);

OAI22xp33_ASAP7_75t_L g14517 ( 
.A1(n_14292),
.A2(n_7714),
.B1(n_6815),
.B2(n_6819),
.Y(n_14517)
);

NOR2xp67_ASAP7_75t_L g14518 ( 
.A(n_14150),
.B(n_8234),
.Y(n_14518)
);

INVx1_ASAP7_75t_L g14519 ( 
.A(n_14267),
.Y(n_14519)
);

OR2x2_ASAP7_75t_L g14520 ( 
.A(n_14251),
.B(n_8234),
.Y(n_14520)
);

INVx2_ASAP7_75t_SL g14521 ( 
.A(n_14229),
.Y(n_14521)
);

INVx1_ASAP7_75t_L g14522 ( 
.A(n_14274),
.Y(n_14522)
);

AND2x2_ASAP7_75t_L g14523 ( 
.A(n_14180),
.B(n_8345),
.Y(n_14523)
);

AOI22xp33_ASAP7_75t_L g14524 ( 
.A1(n_14147),
.A2(n_6955),
.B1(n_6992),
.B2(n_6976),
.Y(n_14524)
);

NAND2xp5_ASAP7_75t_L g14525 ( 
.A(n_14244),
.B(n_8318),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_14245),
.Y(n_14526)
);

A2O1A1Ixp33_ASAP7_75t_L g14527 ( 
.A1(n_14247),
.A2(n_8254),
.B(n_8259),
.C(n_8251),
.Y(n_14527)
);

AOI221xp5_ASAP7_75t_L g14528 ( 
.A1(n_14152),
.A2(n_14281),
.B1(n_14328),
.B2(n_14337),
.C(n_14252),
.Y(n_14528)
);

A2O1A1Ixp33_ASAP7_75t_L g14529 ( 
.A1(n_14306),
.A2(n_8254),
.B(n_8259),
.C(n_8251),
.Y(n_14529)
);

INVx3_ASAP7_75t_L g14530 ( 
.A(n_14330),
.Y(n_14530)
);

INVx1_ASAP7_75t_L g14531 ( 
.A(n_14325),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_14303),
.B(n_8798),
.Y(n_14532)
);

O2A1O1Ixp5_ASAP7_75t_L g14533 ( 
.A1(n_14311),
.A2(n_8264),
.B(n_8270),
.C(n_8254),
.Y(n_14533)
);

AOI311xp33_ASAP7_75t_L g14534 ( 
.A1(n_14288),
.A2(n_14151),
.A3(n_14133),
.B(n_14161),
.C(n_14335),
.Y(n_14534)
);

NOR2xp33_ASAP7_75t_L g14535 ( 
.A(n_14232),
.B(n_6793),
.Y(n_14535)
);

AND2x4_ASAP7_75t_L g14536 ( 
.A(n_14329),
.B(n_8264),
.Y(n_14536)
);

AOI21xp33_ASAP7_75t_L g14537 ( 
.A1(n_14199),
.A2(n_14327),
.B(n_14159),
.Y(n_14537)
);

AOI32xp33_ASAP7_75t_L g14538 ( 
.A1(n_14217),
.A2(n_7163),
.A3(n_7239),
.B1(n_7196),
.B2(n_7133),
.Y(n_14538)
);

AOI22xp33_ASAP7_75t_SL g14539 ( 
.A1(n_14279),
.A2(n_6815),
.B1(n_6819),
.B2(n_6793),
.Y(n_14539)
);

AOI221xp5_ASAP7_75t_L g14540 ( 
.A1(n_14240),
.A2(n_8169),
.B1(n_8174),
.B2(n_8158),
.C(n_8152),
.Y(n_14540)
);

AND2x2_ASAP7_75t_L g14541 ( 
.A(n_14362),
.B(n_14164),
.Y(n_14541)
);

AND2x2_ASAP7_75t_L g14542 ( 
.A(n_14348),
.B(n_14197),
.Y(n_14542)
);

NAND2xp5_ASAP7_75t_L g14543 ( 
.A(n_14352),
.B(n_14257),
.Y(n_14543)
);

INVx1_ASAP7_75t_L g14544 ( 
.A(n_14344),
.Y(n_14544)
);

AOI22xp33_ASAP7_75t_L g14545 ( 
.A1(n_14396),
.A2(n_14181),
.B1(n_14216),
.B2(n_14320),
.Y(n_14545)
);

NAND2xp5_ASAP7_75t_L g14546 ( 
.A(n_14484),
.B(n_14200),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_14347),
.Y(n_14547)
);

AOI22xp33_ASAP7_75t_L g14548 ( 
.A1(n_14389),
.A2(n_14299),
.B1(n_14186),
.B2(n_14302),
.Y(n_14548)
);

INVx1_ASAP7_75t_L g14549 ( 
.A(n_14415),
.Y(n_14549)
);

INVx1_ASAP7_75t_L g14550 ( 
.A(n_14439),
.Y(n_14550)
);

NAND2xp5_ASAP7_75t_L g14551 ( 
.A(n_14367),
.B(n_14128),
.Y(n_14551)
);

AOI22xp33_ASAP7_75t_L g14552 ( 
.A1(n_14379),
.A2(n_14111),
.B1(n_14241),
.B2(n_14316),
.Y(n_14552)
);

NOR2xp33_ASAP7_75t_L g14553 ( 
.A(n_14443),
.B(n_14309),
.Y(n_14553)
);

INVx1_ASAP7_75t_L g14554 ( 
.A(n_14342),
.Y(n_14554)
);

NAND2xp5_ASAP7_75t_SL g14555 ( 
.A(n_14426),
.B(n_8270),
.Y(n_14555)
);

INVx1_ASAP7_75t_SL g14556 ( 
.A(n_14356),
.Y(n_14556)
);

INVx1_ASAP7_75t_SL g14557 ( 
.A(n_14364),
.Y(n_14557)
);

INVx1_ASAP7_75t_L g14558 ( 
.A(n_14345),
.Y(n_14558)
);

AND2x2_ASAP7_75t_L g14559 ( 
.A(n_14435),
.B(n_8345),
.Y(n_14559)
);

NAND2xp5_ASAP7_75t_L g14560 ( 
.A(n_14457),
.B(n_8270),
.Y(n_14560)
);

AND2x2_ASAP7_75t_L g14561 ( 
.A(n_14357),
.B(n_8350),
.Y(n_14561)
);

AND2x2_ASAP7_75t_L g14562 ( 
.A(n_14361),
.B(n_8350),
.Y(n_14562)
);

AND2x2_ASAP7_75t_L g14563 ( 
.A(n_14381),
.B(n_8351),
.Y(n_14563)
);

AND2x4_ASAP7_75t_L g14564 ( 
.A(n_14358),
.B(n_14403),
.Y(n_14564)
);

INVx1_ASAP7_75t_L g14565 ( 
.A(n_14467),
.Y(n_14565)
);

AND2x2_ASAP7_75t_L g14566 ( 
.A(n_14366),
.B(n_8351),
.Y(n_14566)
);

NOR2xp33_ASAP7_75t_L g14567 ( 
.A(n_14445),
.B(n_6793),
.Y(n_14567)
);

AND2x2_ASAP7_75t_L g14568 ( 
.A(n_14350),
.B(n_8351),
.Y(n_14568)
);

NAND2xp5_ASAP7_75t_SL g14569 ( 
.A(n_14494),
.B(n_8283),
.Y(n_14569)
);

INVxp33_ASAP7_75t_L g14570 ( 
.A(n_14504),
.Y(n_14570)
);

INVx1_ASAP7_75t_SL g14571 ( 
.A(n_14346),
.Y(n_14571)
);

INVxp67_ASAP7_75t_L g14572 ( 
.A(n_14511),
.Y(n_14572)
);

NAND2xp5_ASAP7_75t_L g14573 ( 
.A(n_14394),
.B(n_8286),
.Y(n_14573)
);

HB1xp67_ASAP7_75t_L g14574 ( 
.A(n_14374),
.Y(n_14574)
);

NOR3xp33_ASAP7_75t_SL g14575 ( 
.A(n_14437),
.B(n_6362),
.C(n_6409),
.Y(n_14575)
);

NAND2xp5_ASAP7_75t_L g14576 ( 
.A(n_14455),
.B(n_8286),
.Y(n_14576)
);

AND2x2_ASAP7_75t_L g14577 ( 
.A(n_14369),
.B(n_8360),
.Y(n_14577)
);

OAI321xp33_ASAP7_75t_L g14578 ( 
.A1(n_14341),
.A2(n_7767),
.A3(n_7522),
.B1(n_7650),
.B2(n_6482),
.C(n_7350),
.Y(n_14578)
);

NAND2xp5_ASAP7_75t_L g14579 ( 
.A(n_14375),
.B(n_8286),
.Y(n_14579)
);

NAND2xp5_ASAP7_75t_L g14580 ( 
.A(n_14385),
.B(n_8287),
.Y(n_14580)
);

NOR2xp33_ASAP7_75t_L g14581 ( 
.A(n_14427),
.B(n_6815),
.Y(n_14581)
);

AND2x2_ASAP7_75t_L g14582 ( 
.A(n_14451),
.B(n_8360),
.Y(n_14582)
);

OAI221xp5_ASAP7_75t_L g14583 ( 
.A1(n_14539),
.A2(n_6815),
.B1(n_6836),
.B2(n_6834),
.C(n_6819),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_14452),
.B(n_8360),
.Y(n_14584)
);

INVx1_ASAP7_75t_L g14585 ( 
.A(n_14481),
.Y(n_14585)
);

BUFx2_ASAP7_75t_L g14586 ( 
.A(n_14489),
.Y(n_14586)
);

INVx1_ASAP7_75t_SL g14587 ( 
.A(n_14355),
.Y(n_14587)
);

INVx2_ASAP7_75t_L g14588 ( 
.A(n_14377),
.Y(n_14588)
);

OR2x2_ASAP7_75t_L g14589 ( 
.A(n_14434),
.B(n_8287),
.Y(n_14589)
);

NAND2xp5_ASAP7_75t_SL g14590 ( 
.A(n_14510),
.B(n_8287),
.Y(n_14590)
);

AND2x2_ASAP7_75t_L g14591 ( 
.A(n_14453),
.B(n_8362),
.Y(n_14591)
);

NAND2xp5_ASAP7_75t_L g14592 ( 
.A(n_14351),
.B(n_14410),
.Y(n_14592)
);

INVx1_ASAP7_75t_L g14593 ( 
.A(n_14464),
.Y(n_14593)
);

INVxp67_ASAP7_75t_L g14594 ( 
.A(n_14429),
.Y(n_14594)
);

AOI22xp33_ASAP7_75t_L g14595 ( 
.A1(n_14363),
.A2(n_6976),
.B1(n_6992),
.B2(n_6955),
.Y(n_14595)
);

INVx2_ASAP7_75t_SL g14596 ( 
.A(n_14433),
.Y(n_14596)
);

OA21x2_ASAP7_75t_L g14597 ( 
.A1(n_14354),
.A2(n_8296),
.B(n_8291),
.Y(n_14597)
);

NOR2xp33_ASAP7_75t_L g14598 ( 
.A(n_14406),
.B(n_6819),
.Y(n_14598)
);

NOR2xp33_ASAP7_75t_L g14599 ( 
.A(n_14459),
.B(n_6819),
.Y(n_14599)
);

AND2x2_ASAP7_75t_L g14600 ( 
.A(n_14376),
.B(n_8362),
.Y(n_14600)
);

NOR2xp33_ASAP7_75t_L g14601 ( 
.A(n_14425),
.B(n_6834),
.Y(n_14601)
);

INVx1_ASAP7_75t_SL g14602 ( 
.A(n_14378),
.Y(n_14602)
);

AOI22xp33_ASAP7_75t_L g14603 ( 
.A1(n_14359),
.A2(n_6976),
.B1(n_6992),
.B2(n_6955),
.Y(n_14603)
);

OR2x2_ASAP7_75t_L g14604 ( 
.A(n_14449),
.B(n_8296),
.Y(n_14604)
);

OR2x2_ASAP7_75t_L g14605 ( 
.A(n_14461),
.B(n_8296),
.Y(n_14605)
);

OAI22xp5_ASAP7_75t_L g14606 ( 
.A1(n_14447),
.A2(n_14390),
.B1(n_14444),
.B2(n_14446),
.Y(n_14606)
);

INVxp67_ASAP7_75t_L g14607 ( 
.A(n_14499),
.Y(n_14607)
);

INVx1_ASAP7_75t_L g14608 ( 
.A(n_14371),
.Y(n_14608)
);

NOR2xp33_ASAP7_75t_L g14609 ( 
.A(n_14353),
.B(n_6834),
.Y(n_14609)
);

AOI22xp33_ASAP7_75t_L g14610 ( 
.A1(n_14365),
.A2(n_6976),
.B1(n_6992),
.B2(n_6955),
.Y(n_14610)
);

NAND2xp5_ASAP7_75t_L g14611 ( 
.A(n_14450),
.B(n_8299),
.Y(n_14611)
);

NOR2xp33_ASAP7_75t_L g14612 ( 
.A(n_14463),
.B(n_6834),
.Y(n_14612)
);

INVx1_ASAP7_75t_L g14613 ( 
.A(n_14388),
.Y(n_14613)
);

AND2x2_ASAP7_75t_L g14614 ( 
.A(n_14535),
.B(n_8362),
.Y(n_14614)
);

AND2x4_ASAP7_75t_L g14615 ( 
.A(n_14482),
.B(n_8299),
.Y(n_14615)
);

NAND2xp5_ASAP7_75t_L g14616 ( 
.A(n_14491),
.B(n_8299),
.Y(n_14616)
);

NAND2xp5_ASAP7_75t_SL g14617 ( 
.A(n_14414),
.B(n_8302),
.Y(n_14617)
);

INVxp67_ASAP7_75t_L g14618 ( 
.A(n_14349),
.Y(n_14618)
);

INVx2_ASAP7_75t_SL g14619 ( 
.A(n_14397),
.Y(n_14619)
);

NAND3xp33_ASAP7_75t_SL g14620 ( 
.A(n_14343),
.B(n_5981),
.C(n_7354),
.Y(n_14620)
);

OR2x2_ASAP7_75t_L g14621 ( 
.A(n_14340),
.B(n_8302),
.Y(n_14621)
);

AND2x4_ASAP7_75t_L g14622 ( 
.A(n_14368),
.B(n_14521),
.Y(n_14622)
);

NAND2xp5_ASAP7_75t_L g14623 ( 
.A(n_14405),
.B(n_8302),
.Y(n_14623)
);

INVx1_ASAP7_75t_L g14624 ( 
.A(n_14373),
.Y(n_14624)
);

NAND2xp5_ASAP7_75t_L g14625 ( 
.A(n_14485),
.B(n_8311),
.Y(n_14625)
);

AND2x2_ASAP7_75t_L g14626 ( 
.A(n_14473),
.B(n_8367),
.Y(n_14626)
);

NAND2xp5_ASAP7_75t_L g14627 ( 
.A(n_14468),
.B(n_8311),
.Y(n_14627)
);

INVx1_ASAP7_75t_L g14628 ( 
.A(n_14398),
.Y(n_14628)
);

AND2x2_ASAP7_75t_L g14629 ( 
.A(n_14440),
.B(n_8367),
.Y(n_14629)
);

NOR2xp33_ASAP7_75t_L g14630 ( 
.A(n_14460),
.B(n_6834),
.Y(n_14630)
);

AND2x2_ASAP7_75t_L g14631 ( 
.A(n_14416),
.B(n_8367),
.Y(n_14631)
);

INVx2_ASAP7_75t_L g14632 ( 
.A(n_14480),
.Y(n_14632)
);

NAND2x1_ASAP7_75t_L g14633 ( 
.A(n_14384),
.B(n_14475),
.Y(n_14633)
);

NAND2xp5_ASAP7_75t_L g14634 ( 
.A(n_14470),
.B(n_8311),
.Y(n_14634)
);

NOR2xp33_ASAP7_75t_L g14635 ( 
.A(n_14402),
.B(n_6836),
.Y(n_14635)
);

AND2x2_ASAP7_75t_L g14636 ( 
.A(n_14509),
.B(n_8396),
.Y(n_14636)
);

AOI22xp33_ASAP7_75t_L g14637 ( 
.A1(n_14465),
.A2(n_7090),
.B1(n_7127),
.B2(n_7059),
.Y(n_14637)
);

NAND2xp5_ASAP7_75t_L g14638 ( 
.A(n_14471),
.B(n_8316),
.Y(n_14638)
);

INVxp67_ASAP7_75t_SL g14639 ( 
.A(n_14431),
.Y(n_14639)
);

INVx4_ASAP7_75t_L g14640 ( 
.A(n_14530),
.Y(n_14640)
);

INVx1_ASAP7_75t_L g14641 ( 
.A(n_14438),
.Y(n_14641)
);

NOR2xp33_ASAP7_75t_L g14642 ( 
.A(n_14370),
.B(n_6836),
.Y(n_14642)
);

AND2x2_ASAP7_75t_L g14643 ( 
.A(n_14479),
.B(n_8396),
.Y(n_14643)
);

BUFx2_ASAP7_75t_L g14644 ( 
.A(n_14483),
.Y(n_14644)
);

AND2x2_ASAP7_75t_L g14645 ( 
.A(n_14422),
.B(n_8396),
.Y(n_14645)
);

AND2x2_ASAP7_75t_L g14646 ( 
.A(n_14430),
.B(n_8397),
.Y(n_14646)
);

AOI22xp33_ASAP7_75t_SL g14647 ( 
.A1(n_14448),
.A2(n_6903),
.B1(n_6838),
.B2(n_6854),
.Y(n_14647)
);

INVx1_ASAP7_75t_L g14648 ( 
.A(n_14474),
.Y(n_14648)
);

INVx1_ASAP7_75t_L g14649 ( 
.A(n_14432),
.Y(n_14649)
);

INVx1_ASAP7_75t_SL g14650 ( 
.A(n_14360),
.Y(n_14650)
);

AND2x2_ASAP7_75t_L g14651 ( 
.A(n_14458),
.B(n_8397),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_14408),
.Y(n_14652)
);

AND2x4_ASAP7_75t_L g14653 ( 
.A(n_14418),
.B(n_8316),
.Y(n_14653)
);

NAND2xp5_ASAP7_75t_L g14654 ( 
.A(n_14530),
.B(n_14493),
.Y(n_14654)
);

NAND2xp5_ASAP7_75t_L g14655 ( 
.A(n_14486),
.B(n_8316),
.Y(n_14655)
);

NAND2xp5_ASAP7_75t_L g14656 ( 
.A(n_14528),
.B(n_8318),
.Y(n_14656)
);

OR2x2_ASAP7_75t_L g14657 ( 
.A(n_14383),
.B(n_8322),
.Y(n_14657)
);

INVx3_ASAP7_75t_L g14658 ( 
.A(n_14501),
.Y(n_14658)
);

NAND2xp5_ASAP7_75t_L g14659 ( 
.A(n_14413),
.B(n_8322),
.Y(n_14659)
);

NAND2xp5_ASAP7_75t_L g14660 ( 
.A(n_14492),
.B(n_8322),
.Y(n_14660)
);

NAND2xp5_ASAP7_75t_L g14661 ( 
.A(n_14495),
.B(n_8185),
.Y(n_14661)
);

AOI22xp33_ASAP7_75t_L g14662 ( 
.A1(n_14441),
.A2(n_7090),
.B1(n_7127),
.B2(n_7059),
.Y(n_14662)
);

AND2x2_ASAP7_75t_L g14663 ( 
.A(n_14534),
.B(n_8397),
.Y(n_14663)
);

INVx1_ASAP7_75t_L g14664 ( 
.A(n_14409),
.Y(n_14664)
);

INVx1_ASAP7_75t_L g14665 ( 
.A(n_14392),
.Y(n_14665)
);

NAND2xp5_ASAP7_75t_L g14666 ( 
.A(n_14503),
.B(n_8185),
.Y(n_14666)
);

AOI22xp5_ASAP7_75t_L g14667 ( 
.A1(n_14407),
.A2(n_14412),
.B1(n_14487),
.B2(n_14372),
.Y(n_14667)
);

AND2x2_ASAP7_75t_L g14668 ( 
.A(n_14380),
.B(n_8402),
.Y(n_14668)
);

INVxp33_ASAP7_75t_L g14669 ( 
.A(n_14395),
.Y(n_14669)
);

AND2x2_ASAP7_75t_L g14670 ( 
.A(n_14423),
.B(n_14502),
.Y(n_14670)
);

INVxp67_ASAP7_75t_L g14671 ( 
.A(n_14401),
.Y(n_14671)
);

HB1xp67_ASAP7_75t_L g14672 ( 
.A(n_14514),
.Y(n_14672)
);

NAND2x1p5_ASAP7_75t_L g14673 ( 
.A(n_14507),
.B(n_6230),
.Y(n_14673)
);

NAND2xp5_ASAP7_75t_L g14674 ( 
.A(n_14512),
.B(n_8194),
.Y(n_14674)
);

INVx1_ASAP7_75t_L g14675 ( 
.A(n_14420),
.Y(n_14675)
);

AND2x2_ASAP7_75t_L g14676 ( 
.A(n_14531),
.B(n_8402),
.Y(n_14676)
);

OR2x2_ASAP7_75t_L g14677 ( 
.A(n_14500),
.B(n_14478),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_14436),
.Y(n_14678)
);

INVx2_ASAP7_75t_L g14679 ( 
.A(n_14520),
.Y(n_14679)
);

INVxp67_ASAP7_75t_L g14680 ( 
.A(n_14466),
.Y(n_14680)
);

INVx1_ASAP7_75t_L g14681 ( 
.A(n_14454),
.Y(n_14681)
);

NAND2xp5_ASAP7_75t_SL g14682 ( 
.A(n_14517),
.B(n_7650),
.Y(n_14682)
);

AOI22xp33_ASAP7_75t_L g14683 ( 
.A1(n_14428),
.A2(n_7090),
.B1(n_7127),
.B2(n_7059),
.Y(n_14683)
);

INVx1_ASAP7_75t_L g14684 ( 
.A(n_14513),
.Y(n_14684)
);

NAND2xp5_ASAP7_75t_L g14685 ( 
.A(n_14505),
.B(n_8194),
.Y(n_14685)
);

INVx1_ASAP7_75t_L g14686 ( 
.A(n_14519),
.Y(n_14686)
);

OR2x2_ASAP7_75t_L g14687 ( 
.A(n_14522),
.B(n_9317),
.Y(n_14687)
);

NAND2xp5_ASAP7_75t_SL g14688 ( 
.A(n_14417),
.B(n_7767),
.Y(n_14688)
);

INVxp67_ASAP7_75t_L g14689 ( 
.A(n_14526),
.Y(n_14689)
);

NOR2x1p5_ASAP7_75t_L g14690 ( 
.A(n_14525),
.B(n_7331),
.Y(n_14690)
);

AND2x2_ASAP7_75t_L g14691 ( 
.A(n_14404),
.B(n_8402),
.Y(n_14691)
);

INVx2_ASAP7_75t_L g14692 ( 
.A(n_14497),
.Y(n_14692)
);

AOI22xp5_ASAP7_75t_L g14693 ( 
.A1(n_14382),
.A2(n_7374),
.B1(n_7434),
.B2(n_7300),
.Y(n_14693)
);

NAND2xp5_ASAP7_75t_L g14694 ( 
.A(n_14537),
.B(n_8197),
.Y(n_14694)
);

NAND2xp33_ASAP7_75t_L g14695 ( 
.A(n_14523),
.B(n_8417),
.Y(n_14695)
);

INVx1_ASAP7_75t_L g14696 ( 
.A(n_14477),
.Y(n_14696)
);

NAND2xp5_ASAP7_75t_L g14697 ( 
.A(n_14419),
.B(n_8197),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_14490),
.Y(n_14698)
);

INVxp67_ASAP7_75t_L g14699 ( 
.A(n_14496),
.Y(n_14699)
);

NAND2xp5_ASAP7_75t_L g14700 ( 
.A(n_14387),
.B(n_8204),
.Y(n_14700)
);

INVx1_ASAP7_75t_L g14701 ( 
.A(n_14518),
.Y(n_14701)
);

NAND2xp33_ASAP7_75t_L g14702 ( 
.A(n_14456),
.B(n_8417),
.Y(n_14702)
);

NOR2xp33_ASAP7_75t_L g14703 ( 
.A(n_14442),
.B(n_6836),
.Y(n_14703)
);

NAND2xp5_ASAP7_75t_L g14704 ( 
.A(n_14469),
.B(n_14462),
.Y(n_14704)
);

INVx1_ASAP7_75t_L g14705 ( 
.A(n_14498),
.Y(n_14705)
);

OR2x2_ASAP7_75t_L g14706 ( 
.A(n_14411),
.B(n_9317),
.Y(n_14706)
);

NAND2xp5_ASAP7_75t_L g14707 ( 
.A(n_14532),
.B(n_8204),
.Y(n_14707)
);

NAND2xp5_ASAP7_75t_L g14708 ( 
.A(n_14536),
.B(n_8205),
.Y(n_14708)
);

INVx2_ASAP7_75t_L g14709 ( 
.A(n_14536),
.Y(n_14709)
);

OR2x2_ASAP7_75t_L g14710 ( 
.A(n_14515),
.B(n_9371),
.Y(n_14710)
);

AND2x2_ASAP7_75t_L g14711 ( 
.A(n_14524),
.B(n_8417),
.Y(n_14711)
);

NOR2xp33_ASAP7_75t_L g14712 ( 
.A(n_14472),
.B(n_6836),
.Y(n_14712)
);

OR2x2_ASAP7_75t_L g14713 ( 
.A(n_14400),
.B(n_9371),
.Y(n_14713)
);

INVx1_ASAP7_75t_SL g14714 ( 
.A(n_14386),
.Y(n_14714)
);

NAND2xp5_ASAP7_75t_L g14715 ( 
.A(n_14508),
.B(n_14421),
.Y(n_14715)
);

AND2x2_ASAP7_75t_L g14716 ( 
.A(n_14540),
.B(n_8425),
.Y(n_14716)
);

INVx2_ASAP7_75t_L g14717 ( 
.A(n_14476),
.Y(n_14717)
);

NAND2xp5_ASAP7_75t_L g14718 ( 
.A(n_14538),
.B(n_8205),
.Y(n_14718)
);

NAND2xp5_ASAP7_75t_SL g14719 ( 
.A(n_14393),
.B(n_7338),
.Y(n_14719)
);

AND2x2_ASAP7_75t_L g14720 ( 
.A(n_14527),
.B(n_8425),
.Y(n_14720)
);

NAND2xp5_ASAP7_75t_L g14721 ( 
.A(n_14516),
.B(n_8210),
.Y(n_14721)
);

INVx1_ASAP7_75t_SL g14722 ( 
.A(n_14424),
.Y(n_14722)
);

AOI22xp5_ASAP7_75t_L g14723 ( 
.A1(n_14609),
.A2(n_14399),
.B1(n_14488),
.B2(n_14506),
.Y(n_14723)
);

INVx2_ASAP7_75t_L g14724 ( 
.A(n_14564),
.Y(n_14724)
);

AO22x2_ASAP7_75t_L g14725 ( 
.A1(n_14556),
.A2(n_14391),
.B1(n_14533),
.B2(n_14529),
.Y(n_14725)
);

AOI22xp5_ASAP7_75t_L g14726 ( 
.A1(n_14642),
.A2(n_6838),
.B1(n_6903),
.B2(n_6854),
.Y(n_14726)
);

INVx1_ASAP7_75t_L g14727 ( 
.A(n_14574),
.Y(n_14727)
);

NAND4xp75_ASAP7_75t_L g14728 ( 
.A(n_14549),
.B(n_9467),
.C(n_9471),
.D(n_6057),
.Y(n_14728)
);

OAI322xp33_ASAP7_75t_L g14729 ( 
.A1(n_14633),
.A2(n_8440),
.A3(n_8429),
.B1(n_8452),
.B2(n_8467),
.C1(n_8435),
.C2(n_8425),
.Y(n_14729)
);

INVx1_ASAP7_75t_L g14730 ( 
.A(n_14586),
.Y(n_14730)
);

INVx1_ASAP7_75t_L g14731 ( 
.A(n_14644),
.Y(n_14731)
);

AOI22xp5_ASAP7_75t_L g14732 ( 
.A1(n_14571),
.A2(n_6838),
.B1(n_6903),
.B2(n_6854),
.Y(n_14732)
);

INVx1_ASAP7_75t_L g14733 ( 
.A(n_14564),
.Y(n_14733)
);

INVx1_ASAP7_75t_L g14734 ( 
.A(n_14544),
.Y(n_14734)
);

OA22x2_ASAP7_75t_L g14735 ( 
.A1(n_14667),
.A2(n_8213),
.B1(n_8217),
.B2(n_8210),
.Y(n_14735)
);

INVx1_ASAP7_75t_L g14736 ( 
.A(n_14547),
.Y(n_14736)
);

OA22x2_ASAP7_75t_L g14737 ( 
.A1(n_14557),
.A2(n_8217),
.B1(n_8225),
.B2(n_8213),
.Y(n_14737)
);

AND4x1_ASAP7_75t_L g14738 ( 
.A(n_14585),
.B(n_7081),
.C(n_5981),
.D(n_6057),
.Y(n_14738)
);

INVx1_ASAP7_75t_L g14739 ( 
.A(n_14672),
.Y(n_14739)
);

INVx1_ASAP7_75t_L g14740 ( 
.A(n_14554),
.Y(n_14740)
);

OAI22xp5_ASAP7_75t_L g14741 ( 
.A1(n_14595),
.A2(n_14610),
.B1(n_14603),
.B2(n_14545),
.Y(n_14741)
);

BUFx4_ASAP7_75t_R g14742 ( 
.A(n_14717),
.Y(n_14742)
);

OAI22xp5_ASAP7_75t_L g14743 ( 
.A1(n_14583),
.A2(n_8435),
.B1(n_8637),
.B2(n_8484),
.Y(n_14743)
);

AOI22xp5_ASAP7_75t_L g14744 ( 
.A1(n_14567),
.A2(n_6838),
.B1(n_6903),
.B2(n_6854),
.Y(n_14744)
);

INVx1_ASAP7_75t_L g14745 ( 
.A(n_14592),
.Y(n_14745)
);

AOI221xp5_ASAP7_75t_L g14746 ( 
.A1(n_14578),
.A2(n_8227),
.B1(n_8237),
.B2(n_8230),
.C(n_8225),
.Y(n_14746)
);

INVx1_ASAP7_75t_L g14747 ( 
.A(n_14622),
.Y(n_14747)
);

OA22x2_ASAP7_75t_L g14748 ( 
.A1(n_14596),
.A2(n_14619),
.B1(n_14714),
.B2(n_14722),
.Y(n_14748)
);

NAND4xp25_ASAP7_75t_L g14749 ( 
.A(n_14581),
.B(n_6667),
.C(n_6606),
.D(n_6230),
.Y(n_14749)
);

OA22x2_ASAP7_75t_SL g14750 ( 
.A1(n_14613),
.A2(n_8230),
.B1(n_8237),
.B2(n_8227),
.Y(n_14750)
);

INVx1_ASAP7_75t_L g14751 ( 
.A(n_14622),
.Y(n_14751)
);

OA22x2_ASAP7_75t_L g14752 ( 
.A1(n_14550),
.A2(n_8243),
.B1(n_8247),
.B2(n_8240),
.Y(n_14752)
);

INVx1_ASAP7_75t_L g14753 ( 
.A(n_14643),
.Y(n_14753)
);

INVx1_ASAP7_75t_L g14754 ( 
.A(n_14640),
.Y(n_14754)
);

INVx1_ASAP7_75t_L g14755 ( 
.A(n_14640),
.Y(n_14755)
);

INVx1_ASAP7_75t_L g14756 ( 
.A(n_14694),
.Y(n_14756)
);

HB1xp67_ASAP7_75t_L g14757 ( 
.A(n_14597),
.Y(n_14757)
);

AOI22xp5_ASAP7_75t_L g14758 ( 
.A1(n_14601),
.A2(n_6838),
.B1(n_6903),
.B2(n_6854),
.Y(n_14758)
);

INVx1_ASAP7_75t_L g14759 ( 
.A(n_14663),
.Y(n_14759)
);

INVx2_ASAP7_75t_L g14760 ( 
.A(n_14658),
.Y(n_14760)
);

NAND4xp75_ASAP7_75t_L g14761 ( 
.A(n_14541),
.B(n_9471),
.C(n_9467),
.D(n_8796),
.Y(n_14761)
);

AOI22xp5_ASAP7_75t_L g14762 ( 
.A1(n_14612),
.A2(n_6904),
.B1(n_9471),
.B2(n_9467),
.Y(n_14762)
);

AND4x1_ASAP7_75t_L g14763 ( 
.A(n_14553),
.B(n_7382),
.C(n_7377),
.D(n_7384),
.Y(n_14763)
);

INVx2_ASAP7_75t_L g14764 ( 
.A(n_14597),
.Y(n_14764)
);

OAI322xp33_ASAP7_75t_L g14765 ( 
.A1(n_14618),
.A2(n_8452),
.A3(n_8435),
.B1(n_8467),
.B2(n_8470),
.C1(n_8440),
.C2(n_8429),
.Y(n_14765)
);

AOI22xp5_ASAP7_75t_L g14766 ( 
.A1(n_14598),
.A2(n_6904),
.B1(n_9471),
.B2(n_7090),
.Y(n_14766)
);

AOI22xp5_ASAP7_75t_L g14767 ( 
.A1(n_14599),
.A2(n_6904),
.B1(n_7090),
.B2(n_7059),
.Y(n_14767)
);

INVx1_ASAP7_75t_SL g14768 ( 
.A(n_14587),
.Y(n_14768)
);

HB1xp67_ASAP7_75t_L g14769 ( 
.A(n_14673),
.Y(n_14769)
);

INVx1_ASAP7_75t_L g14770 ( 
.A(n_14588),
.Y(n_14770)
);

OAI31xp33_ASAP7_75t_L g14771 ( 
.A1(n_14690),
.A2(n_8308),
.A3(n_8332),
.B(n_8257),
.Y(n_14771)
);

NAND4xp25_ASAP7_75t_SL g14772 ( 
.A(n_14552),
.B(n_7396),
.C(n_8809),
.D(n_8243),
.Y(n_14772)
);

INVx1_ASAP7_75t_L g14773 ( 
.A(n_14656),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_14654),
.Y(n_14774)
);

INVx1_ASAP7_75t_L g14775 ( 
.A(n_14560),
.Y(n_14775)
);

AOI221xp5_ASAP7_75t_L g14776 ( 
.A1(n_14703),
.A2(n_8247),
.B1(n_8250),
.B2(n_8249),
.C(n_8240),
.Y(n_14776)
);

INVx1_ASAP7_75t_L g14777 ( 
.A(n_14561),
.Y(n_14777)
);

INVx1_ASAP7_75t_L g14778 ( 
.A(n_14562),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14563),
.Y(n_14779)
);

INVx1_ASAP7_75t_L g14780 ( 
.A(n_14655),
.Y(n_14780)
);

OAI22xp33_ASAP7_75t_SL g14781 ( 
.A1(n_14719),
.A2(n_6904),
.B1(n_7127),
.B2(n_7059),
.Y(n_14781)
);

AOI22xp5_ASAP7_75t_L g14782 ( 
.A1(n_14630),
.A2(n_6904),
.B1(n_7203),
.B2(n_7127),
.Y(n_14782)
);

INVx1_ASAP7_75t_L g14783 ( 
.A(n_14566),
.Y(n_14783)
);

AO22x2_ASAP7_75t_L g14784 ( 
.A1(n_14709),
.A2(n_8440),
.B1(n_8452),
.B2(n_8429),
.Y(n_14784)
);

NOR4xp25_ASAP7_75t_L g14785 ( 
.A(n_14546),
.B(n_8257),
.C(n_8258),
.D(n_8249),
.Y(n_14785)
);

INVx1_ASAP7_75t_L g14786 ( 
.A(n_14559),
.Y(n_14786)
);

INVx2_ASAP7_75t_L g14787 ( 
.A(n_14615),
.Y(n_14787)
);

OA22x2_ASAP7_75t_L g14788 ( 
.A1(n_14602),
.A2(n_8258),
.B1(n_8266),
.B2(n_8250),
.Y(n_14788)
);

INVx2_ASAP7_75t_SL g14789 ( 
.A(n_14615),
.Y(n_14789)
);

AOI31xp33_ASAP7_75t_L g14790 ( 
.A1(n_14570),
.A2(n_6482),
.A3(n_7439),
.B(n_7437),
.Y(n_14790)
);

OAI31xp33_ASAP7_75t_L g14791 ( 
.A1(n_14606),
.A2(n_8320),
.A3(n_8348),
.B(n_8277),
.Y(n_14791)
);

NAND4xp25_ASAP7_75t_SL g14792 ( 
.A(n_14548),
.B(n_8809),
.C(n_8267),
.D(n_8268),
.Y(n_14792)
);

OAI22xp5_ASAP7_75t_L g14793 ( 
.A1(n_14647),
.A2(n_8495),
.B1(n_8524),
.B2(n_8475),
.Y(n_14793)
);

AOI22x1_ASAP7_75t_L g14794 ( 
.A1(n_14650),
.A2(n_6403),
.B1(n_6407),
.B2(n_6231),
.Y(n_14794)
);

OAI322xp33_ASAP7_75t_L g14795 ( 
.A1(n_14677),
.A2(n_8475),
.A3(n_8470),
.B1(n_8481),
.B2(n_8484),
.C1(n_8472),
.C2(n_8467),
.Y(n_14795)
);

AOI22x1_ASAP7_75t_L g14796 ( 
.A1(n_14632),
.A2(n_6407),
.B1(n_6439),
.B2(n_6403),
.Y(n_14796)
);

OA22x2_ASAP7_75t_L g14797 ( 
.A1(n_14705),
.A2(n_8267),
.B1(n_8268),
.B2(n_8266),
.Y(n_14797)
);

OAI322xp33_ASAP7_75t_L g14798 ( 
.A1(n_14635),
.A2(n_8481),
.A3(n_8472),
.B1(n_8484),
.B2(n_8490),
.C1(n_8475),
.C2(n_8470),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_14582),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_14584),
.Y(n_14800)
);

NAND4xp75_ASAP7_75t_L g14801 ( 
.A(n_14542),
.B(n_8790),
.C(n_8793),
.D(n_8789),
.Y(n_14801)
);

INVx1_ASAP7_75t_L g14802 ( 
.A(n_14591),
.Y(n_14802)
);

INVx1_ASAP7_75t_L g14803 ( 
.A(n_14565),
.Y(n_14803)
);

NAND4xp75_ASAP7_75t_L g14804 ( 
.A(n_14551),
.B(n_8790),
.C(n_8793),
.D(n_8789),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_14624),
.Y(n_14805)
);

O2A1O1Ixp33_ASAP7_75t_L g14806 ( 
.A1(n_14543),
.A2(n_8305),
.B(n_8307),
.C(n_8277),
.Y(n_14806)
);

BUFx4_ASAP7_75t_R g14807 ( 
.A(n_14679),
.Y(n_14807)
);

OA22x2_ASAP7_75t_L g14808 ( 
.A1(n_14593),
.A2(n_8307),
.B1(n_8308),
.B2(n_8305),
.Y(n_14808)
);

INVx1_ASAP7_75t_L g14809 ( 
.A(n_14605),
.Y(n_14809)
);

AOI22xp5_ASAP7_75t_L g14810 ( 
.A1(n_14712),
.A2(n_7203),
.B1(n_7270),
.B2(n_7221),
.Y(n_14810)
);

AND4x1_ASAP7_75t_L g14811 ( 
.A(n_14608),
.B(n_6409),
.C(n_7360),
.D(n_7357),
.Y(n_14811)
);

OAI322xp33_ASAP7_75t_L g14812 ( 
.A1(n_14704),
.A2(n_8491),
.A3(n_8481),
.B1(n_8495),
.B2(n_8501),
.C1(n_8490),
.C2(n_8472),
.Y(n_14812)
);

INVx1_ASAP7_75t_L g14813 ( 
.A(n_14568),
.Y(n_14813)
);

INVx2_ASAP7_75t_L g14814 ( 
.A(n_14589),
.Y(n_14814)
);

INVx1_ASAP7_75t_L g14815 ( 
.A(n_14569),
.Y(n_14815)
);

INVx2_ASAP7_75t_L g14816 ( 
.A(n_14645),
.Y(n_14816)
);

NAND2x1_ASAP7_75t_SL g14817 ( 
.A(n_14628),
.B(n_8309),
.Y(n_14817)
);

INVx1_ASAP7_75t_L g14818 ( 
.A(n_14590),
.Y(n_14818)
);

OAI22xp5_ASAP7_75t_L g14819 ( 
.A1(n_14683),
.A2(n_8529),
.B1(n_8545),
.B2(n_8501),
.Y(n_14819)
);

INVx1_ASAP7_75t_L g14820 ( 
.A(n_14641),
.Y(n_14820)
);

OAI322xp33_ASAP7_75t_L g14821 ( 
.A1(n_14715),
.A2(n_8501),
.A3(n_8491),
.B1(n_8521),
.B2(n_8524),
.C1(n_8495),
.C2(n_8490),
.Y(n_14821)
);

AOI22xp5_ASAP7_75t_L g14822 ( 
.A1(n_14620),
.A2(n_7203),
.B1(n_7270),
.B2(n_7221),
.Y(n_14822)
);

OA22x2_ASAP7_75t_L g14823 ( 
.A1(n_14616),
.A2(n_8310),
.B1(n_8314),
.B2(n_8309),
.Y(n_14823)
);

AND4x1_ASAP7_75t_L g14824 ( 
.A(n_14558),
.B(n_7480),
.C(n_7457),
.D(n_6436),
.Y(n_14824)
);

AOI22xp5_ASAP7_75t_L g14825 ( 
.A1(n_14572),
.A2(n_7203),
.B1(n_7270),
.B2(n_7221),
.Y(n_14825)
);

OAI22xp5_ASAP7_75t_L g14826 ( 
.A1(n_14689),
.A2(n_8521),
.B1(n_8643),
.B2(n_8561),
.Y(n_14826)
);

BUFx3_ASAP7_75t_L g14827 ( 
.A(n_14670),
.Y(n_14827)
);

INVx1_ASAP7_75t_SL g14828 ( 
.A(n_14600),
.Y(n_14828)
);

INVx1_ASAP7_75t_L g14829 ( 
.A(n_14648),
.Y(n_14829)
);

INVx1_ASAP7_75t_L g14830 ( 
.A(n_14580),
.Y(n_14830)
);

INVx1_ASAP7_75t_L g14831 ( 
.A(n_14623),
.Y(n_14831)
);

INVx1_ASAP7_75t_L g14832 ( 
.A(n_14611),
.Y(n_14832)
);

OAI221xp5_ASAP7_75t_SL g14833 ( 
.A1(n_14604),
.A2(n_7733),
.B1(n_7748),
.B2(n_7692),
.C(n_7677),
.Y(n_14833)
);

INVx1_ASAP7_75t_SL g14834 ( 
.A(n_14629),
.Y(n_14834)
);

INVx1_ASAP7_75t_L g14835 ( 
.A(n_14573),
.Y(n_14835)
);

NAND4xp75_ASAP7_75t_L g14836 ( 
.A(n_14686),
.B(n_8803),
.C(n_8310),
.D(n_8319),
.Y(n_14836)
);

OAI22xp5_ASAP7_75t_L g14837 ( 
.A1(n_14637),
.A2(n_14662),
.B1(n_14575),
.B2(n_14607),
.Y(n_14837)
);

HB1xp67_ASAP7_75t_L g14838 ( 
.A(n_14701),
.Y(n_14838)
);

INVx1_ASAP7_75t_L g14839 ( 
.A(n_14626),
.Y(n_14839)
);

AOI221xp5_ASAP7_75t_L g14840 ( 
.A1(n_14702),
.A2(n_8319),
.B1(n_8326),
.B2(n_8320),
.C(n_8314),
.Y(n_14840)
);

INVx1_ASAP7_75t_L g14841 ( 
.A(n_14621),
.Y(n_14841)
);

INVx1_ASAP7_75t_L g14842 ( 
.A(n_14577),
.Y(n_14842)
);

OA22x2_ASAP7_75t_L g14843 ( 
.A1(n_14682),
.A2(n_8329),
.B1(n_8332),
.B2(n_8326),
.Y(n_14843)
);

INVx1_ASAP7_75t_L g14844 ( 
.A(n_14576),
.Y(n_14844)
);

AOI22xp5_ASAP7_75t_L g14845 ( 
.A1(n_14594),
.A2(n_7203),
.B1(n_7270),
.B2(n_7221),
.Y(n_14845)
);

HB1xp67_ASAP7_75t_L g14846 ( 
.A(n_14653),
.Y(n_14846)
);

AOI22xp5_ASAP7_75t_L g14847 ( 
.A1(n_14614),
.A2(n_7221),
.B1(n_7300),
.B2(n_7270),
.Y(n_14847)
);

AND4x1_ASAP7_75t_L g14848 ( 
.A(n_14665),
.B(n_6436),
.C(n_7296),
.D(n_7279),
.Y(n_14848)
);

INVx1_ASAP7_75t_L g14849 ( 
.A(n_14625),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_14659),
.Y(n_14850)
);

OAI322xp33_ASAP7_75t_L g14851 ( 
.A1(n_14699),
.A2(n_8529),
.A3(n_8521),
.B1(n_8532),
.B2(n_8543),
.C1(n_8524),
.C2(n_8491),
.Y(n_14851)
);

AOI22xp5_ASAP7_75t_L g14852 ( 
.A1(n_14631),
.A2(n_7300),
.B1(n_7365),
.B2(n_7319),
.Y(n_14852)
);

OAI322xp33_ASAP7_75t_L g14853 ( 
.A1(n_14671),
.A2(n_8545),
.A3(n_8532),
.B1(n_8554),
.B2(n_8561),
.C1(n_8543),
.C2(n_8529),
.Y(n_14853)
);

NAND4xp75_ASAP7_75t_L g14854 ( 
.A(n_14675),
.B(n_8803),
.C(n_8329),
.D(n_8335),
.Y(n_14854)
);

AOI22xp5_ASAP7_75t_L g14855 ( 
.A1(n_14646),
.A2(n_7300),
.B1(n_7365),
.B2(n_7319),
.Y(n_14855)
);

AND4x1_ASAP7_75t_L g14856 ( 
.A(n_14681),
.B(n_7315),
.C(n_7299),
.D(n_7314),
.Y(n_14856)
);

NAND4xp75_ASAP7_75t_L g14857 ( 
.A(n_14678),
.B(n_8774),
.C(n_8778),
.D(n_8773),
.Y(n_14857)
);

AND4x1_ASAP7_75t_L g14858 ( 
.A(n_14649),
.B(n_7311),
.C(n_7317),
.D(n_7409),
.Y(n_14858)
);

OAI322xp33_ASAP7_75t_L g14859 ( 
.A1(n_14680),
.A2(n_8554),
.A3(n_8543),
.B1(n_8561),
.B2(n_8563),
.C1(n_8545),
.C2(n_8532),
.Y(n_14859)
);

OAI22xp5_ASAP7_75t_L g14860 ( 
.A1(n_14693),
.A2(n_8608),
.B1(n_8657),
.B2(n_8589),
.Y(n_14860)
);

INVx1_ASAP7_75t_L g14861 ( 
.A(n_14660),
.Y(n_14861)
);

AOI22xp5_ASAP7_75t_L g14862 ( 
.A1(n_14711),
.A2(n_7300),
.B1(n_7365),
.B2(n_7319),
.Y(n_14862)
);

HB1xp67_ASAP7_75t_L g14863 ( 
.A(n_14653),
.Y(n_14863)
);

INVx1_ASAP7_75t_L g14864 ( 
.A(n_14661),
.Y(n_14864)
);

AOI22xp5_ASAP7_75t_L g14865 ( 
.A1(n_14668),
.A2(n_7319),
.B1(n_7373),
.B2(n_7365),
.Y(n_14865)
);

AO22x2_ASAP7_75t_L g14866 ( 
.A1(n_14652),
.A2(n_8563),
.B1(n_8565),
.B2(n_8554),
.Y(n_14866)
);

INVx1_ASAP7_75t_L g14867 ( 
.A(n_14666),
.Y(n_14867)
);

INVx1_ASAP7_75t_L g14868 ( 
.A(n_14674),
.Y(n_14868)
);

NAND4xp75_ASAP7_75t_L g14869 ( 
.A(n_14664),
.B(n_14684),
.C(n_14696),
.D(n_14698),
.Y(n_14869)
);

INVx2_ASAP7_75t_L g14870 ( 
.A(n_14657),
.Y(n_14870)
);

INVx1_ASAP7_75t_L g14871 ( 
.A(n_14685),
.Y(n_14871)
);

OAI22xp5_ASAP7_75t_L g14872 ( 
.A1(n_14718),
.A2(n_8662),
.B1(n_8763),
.B2(n_8563),
.Y(n_14872)
);

OAI22xp33_ASAP7_75t_L g14873 ( 
.A1(n_14669),
.A2(n_8581),
.B1(n_8589),
.B2(n_8565),
.Y(n_14873)
);

AOI221xp5_ASAP7_75t_L g14874 ( 
.A1(n_14579),
.A2(n_8799),
.B1(n_8796),
.B2(n_8335),
.C(n_8339),
.Y(n_14874)
);

AOI31xp33_ASAP7_75t_L g14875 ( 
.A1(n_14639),
.A2(n_6482),
.A3(n_6440),
.B(n_6423),
.Y(n_14875)
);

AOI221xp5_ASAP7_75t_L g14876 ( 
.A1(n_14617),
.A2(n_8337),
.B1(n_8348),
.B2(n_8339),
.C(n_8334),
.Y(n_14876)
);

INVx3_ASAP7_75t_L g14877 ( 
.A(n_14692),
.Y(n_14877)
);

AOI22xp5_ASAP7_75t_L g14878 ( 
.A1(n_14688),
.A2(n_7319),
.B1(n_7373),
.B2(n_7365),
.Y(n_14878)
);

NAND4xp25_ASAP7_75t_SL g14879 ( 
.A(n_14707),
.B(n_8774),
.C(n_8778),
.D(n_8773),
.Y(n_14879)
);

AOI22xp33_ASAP7_75t_L g14880 ( 
.A1(n_14636),
.A2(n_7374),
.B1(n_7434),
.B2(n_7373),
.Y(n_14880)
);

AOI22xp5_ASAP7_75t_L g14881 ( 
.A1(n_14695),
.A2(n_7373),
.B1(n_7434),
.B2(n_7374),
.Y(n_14881)
);

NAND4xp75_ASAP7_75t_L g14882 ( 
.A(n_14651),
.B(n_8785),
.C(n_8799),
.D(n_8781),
.Y(n_14882)
);

OAI22xp5_ASAP7_75t_L g14883 ( 
.A1(n_14713),
.A2(n_8608),
.B1(n_8657),
.B2(n_8589),
.Y(n_14883)
);

NOR4xp25_ASAP7_75t_L g14884 ( 
.A(n_14676),
.B(n_8337),
.C(n_8352),
.D(n_8334),
.Y(n_14884)
);

AOI22xp5_ASAP7_75t_L g14885 ( 
.A1(n_14555),
.A2(n_7373),
.B1(n_7434),
.B2(n_7374),
.Y(n_14885)
);

AND2x2_ASAP7_75t_L g14886 ( 
.A(n_14691),
.B(n_8565),
.Y(n_14886)
);

AOI22xp5_ASAP7_75t_L g14887 ( 
.A1(n_14716),
.A2(n_7374),
.B1(n_7456),
.B2(n_7434),
.Y(n_14887)
);

AOI22xp5_ASAP7_75t_L g14888 ( 
.A1(n_14720),
.A2(n_7456),
.B1(n_7512),
.B2(n_7484),
.Y(n_14888)
);

OA22x2_ASAP7_75t_L g14889 ( 
.A1(n_14638),
.A2(n_8354),
.B1(n_8358),
.B2(n_8352),
.Y(n_14889)
);

INVx1_ASAP7_75t_L g14890 ( 
.A(n_14721),
.Y(n_14890)
);

OAI322xp33_ASAP7_75t_L g14891 ( 
.A1(n_14687),
.A2(n_8608),
.A3(n_8598),
.B1(n_8618),
.B2(n_8623),
.C1(n_8601),
.C2(n_8581),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_14700),
.Y(n_14892)
);

HB1xp67_ASAP7_75t_L g14893 ( 
.A(n_14627),
.Y(n_14893)
);

AO22x2_ASAP7_75t_L g14894 ( 
.A1(n_14708),
.A2(n_14634),
.B1(n_14697),
.B2(n_14710),
.Y(n_14894)
);

AOI22xp33_ASAP7_75t_L g14895 ( 
.A1(n_14706),
.A2(n_7484),
.B1(n_7512),
.B2(n_7456),
.Y(n_14895)
);

INVx1_ASAP7_75t_L g14896 ( 
.A(n_14574),
.Y(n_14896)
);

AO22x2_ASAP7_75t_L g14897 ( 
.A1(n_14556),
.A2(n_8598),
.B1(n_8601),
.B2(n_8581),
.Y(n_14897)
);

NAND4xp25_ASAP7_75t_L g14898 ( 
.A(n_14642),
.B(n_6667),
.C(n_6606),
.D(n_6403),
.Y(n_14898)
);

AOI22xp5_ASAP7_75t_L g14899 ( 
.A1(n_14609),
.A2(n_7456),
.B1(n_7512),
.B2(n_7484),
.Y(n_14899)
);

INVx1_ASAP7_75t_L g14900 ( 
.A(n_14574),
.Y(n_14900)
);

OAI22xp5_ASAP7_75t_L g14901 ( 
.A1(n_14595),
.A2(n_8723),
.B1(n_8783),
.B2(n_8647),
.Y(n_14901)
);

NOR2x1_ASAP7_75t_L g14902 ( 
.A(n_14640),
.B(n_8354),
.Y(n_14902)
);

AO22x2_ASAP7_75t_L g14903 ( 
.A1(n_14556),
.A2(n_8601),
.B1(n_8623),
.B2(n_8618),
.Y(n_14903)
);

INVxp67_ASAP7_75t_L g14904 ( 
.A(n_14642),
.Y(n_14904)
);

INVx1_ASAP7_75t_L g14905 ( 
.A(n_14574),
.Y(n_14905)
);

NAND4xp75_ASAP7_75t_L g14906 ( 
.A(n_14549),
.B(n_8781),
.C(n_8785),
.D(n_8770),
.Y(n_14906)
);

NAND2xp5_ASAP7_75t_SL g14907 ( 
.A(n_14747),
.B(n_8598),
.Y(n_14907)
);

AOI21xp5_ASAP7_75t_L g14908 ( 
.A1(n_14751),
.A2(n_14731),
.B(n_14768),
.Y(n_14908)
);

AOI22xp5_ASAP7_75t_L g14909 ( 
.A1(n_14730),
.A2(n_7456),
.B1(n_7512),
.B2(n_7484),
.Y(n_14909)
);

NAND2xp5_ASAP7_75t_L g14910 ( 
.A(n_14733),
.B(n_8618),
.Y(n_14910)
);

AND2x2_ASAP7_75t_L g14911 ( 
.A(n_14724),
.B(n_8623),
.Y(n_14911)
);

INVx1_ASAP7_75t_L g14912 ( 
.A(n_14846),
.Y(n_14912)
);

AOI21xp33_ASAP7_75t_L g14913 ( 
.A1(n_14748),
.A2(n_6407),
.B(n_6403),
.Y(n_14913)
);

NAND2xp5_ASAP7_75t_L g14914 ( 
.A(n_14727),
.B(n_8625),
.Y(n_14914)
);

NOR3x1_ASAP7_75t_L g14915 ( 
.A(n_14869),
.B(n_5734),
.C(n_8358),
.Y(n_14915)
);

NOR3x1_ASAP7_75t_L g14916 ( 
.A(n_14898),
.B(n_8365),
.C(n_8364),
.Y(n_14916)
);

AOI211x1_ASAP7_75t_SL g14917 ( 
.A1(n_14741),
.A2(n_8787),
.B(n_8805),
.C(n_8784),
.Y(n_14917)
);

OAI21xp33_ASAP7_75t_L g14918 ( 
.A1(n_14732),
.A2(n_6098),
.B(n_8364),
.Y(n_14918)
);

NOR3xp33_ASAP7_75t_L g14919 ( 
.A(n_14877),
.B(n_6439),
.C(n_6403),
.Y(n_14919)
);

INVx1_ASAP7_75t_L g14920 ( 
.A(n_14863),
.Y(n_14920)
);

INVx2_ASAP7_75t_L g14921 ( 
.A(n_14817),
.Y(n_14921)
);

OAI31xp33_ASAP7_75t_L g14922 ( 
.A1(n_14896),
.A2(n_14900),
.A3(n_14905),
.B(n_14792),
.Y(n_14922)
);

OAI21xp5_ASAP7_75t_L g14923 ( 
.A1(n_14904),
.A2(n_8369),
.B(n_8365),
.Y(n_14923)
);

NOR3xp33_ASAP7_75t_L g14924 ( 
.A(n_14820),
.B(n_6439),
.C(n_6407),
.Y(n_14924)
);

AND2x2_ASAP7_75t_L g14925 ( 
.A(n_14760),
.B(n_8625),
.Y(n_14925)
);

NOR3xp33_ASAP7_75t_L g14926 ( 
.A(n_14829),
.B(n_6439),
.C(n_6407),
.Y(n_14926)
);

AOI21xp5_ASAP7_75t_L g14927 ( 
.A1(n_14754),
.A2(n_8637),
.B(n_8625),
.Y(n_14927)
);

AOI22xp5_ASAP7_75t_L g14928 ( 
.A1(n_14770),
.A2(n_7484),
.B1(n_7527),
.B2(n_7512),
.Y(n_14928)
);

A2O1A1Ixp33_ASAP7_75t_L g14929 ( 
.A1(n_14791),
.A2(n_8369),
.B(n_8373),
.C(n_8372),
.Y(n_14929)
);

NOR3xp33_ASAP7_75t_L g14930 ( 
.A(n_14803),
.B(n_6624),
.C(n_6439),
.Y(n_14930)
);

AO22x2_ASAP7_75t_L g14931 ( 
.A1(n_14789),
.A2(n_8643),
.B1(n_8645),
.B2(n_8637),
.Y(n_14931)
);

NOR2x1_ASAP7_75t_L g14932 ( 
.A(n_14764),
.B(n_8373),
.Y(n_14932)
);

NAND2xp5_ASAP7_75t_L g14933 ( 
.A(n_14740),
.B(n_8643),
.Y(n_14933)
);

NOR3xp33_ASAP7_75t_SL g14934 ( 
.A(n_14734),
.B(n_6387),
.C(n_6035),
.Y(n_14934)
);

NAND2xp5_ASAP7_75t_L g14935 ( 
.A(n_14755),
.B(n_8645),
.Y(n_14935)
);

INVx1_ASAP7_75t_L g14936 ( 
.A(n_14757),
.Y(n_14936)
);

NAND2xp5_ASAP7_75t_L g14937 ( 
.A(n_14736),
.B(n_8645),
.Y(n_14937)
);

AOI21xp5_ASAP7_75t_L g14938 ( 
.A1(n_14769),
.A2(n_8655),
.B(n_8647),
.Y(n_14938)
);

AOI211xp5_ASAP7_75t_L g14939 ( 
.A1(n_14837),
.A2(n_8372),
.B(n_8379),
.C(n_8378),
.Y(n_14939)
);

AOI211xp5_ASAP7_75t_L g14940 ( 
.A1(n_14759),
.A2(n_8378),
.B(n_8380),
.C(n_8379),
.Y(n_14940)
);

AOI22xp5_ASAP7_75t_L g14941 ( 
.A1(n_14774),
.A2(n_14805),
.B1(n_14726),
.B2(n_14745),
.Y(n_14941)
);

INVx1_ASAP7_75t_L g14942 ( 
.A(n_14902),
.Y(n_14942)
);

NAND2xp5_ASAP7_75t_L g14943 ( 
.A(n_14753),
.B(n_8647),
.Y(n_14943)
);

AND2x2_ASAP7_75t_L g14944 ( 
.A(n_14827),
.B(n_8655),
.Y(n_14944)
);

INVxp67_ASAP7_75t_SL g14945 ( 
.A(n_14787),
.Y(n_14945)
);

NAND2xp5_ASAP7_75t_L g14946 ( 
.A(n_14828),
.B(n_8655),
.Y(n_14946)
);

AOI22xp5_ASAP7_75t_L g14947 ( 
.A1(n_14772),
.A2(n_7527),
.B1(n_8385),
.B2(n_8380),
.Y(n_14947)
);

AOI22xp5_ASAP7_75t_L g14948 ( 
.A1(n_14749),
.A2(n_7527),
.B1(n_8386),
.B2(n_8385),
.Y(n_14948)
);

NAND2xp5_ASAP7_75t_L g14949 ( 
.A(n_14834),
.B(n_8657),
.Y(n_14949)
);

AOI211x1_ASAP7_75t_L g14950 ( 
.A1(n_14739),
.A2(n_8770),
.B(n_8766),
.C(n_8386),
.Y(n_14950)
);

NOR2xp67_ASAP7_75t_L g14951 ( 
.A(n_14809),
.B(n_8387),
.Y(n_14951)
);

AOI21xp5_ASAP7_75t_L g14952 ( 
.A1(n_14838),
.A2(n_8662),
.B(n_8661),
.Y(n_14952)
);

AOI211xp5_ASAP7_75t_L g14953 ( 
.A1(n_14780),
.A2(n_8387),
.B(n_8390),
.C(n_8389),
.Y(n_14953)
);

NOR2x1_ASAP7_75t_L g14954 ( 
.A(n_14815),
.B(n_8389),
.Y(n_14954)
);

INVx1_ASAP7_75t_L g14955 ( 
.A(n_14725),
.Y(n_14955)
);

INVx2_ASAP7_75t_L g14956 ( 
.A(n_14807),
.Y(n_14956)
);

INVx1_ASAP7_75t_L g14957 ( 
.A(n_14725),
.Y(n_14957)
);

NAND2xp5_ASAP7_75t_L g14958 ( 
.A(n_14777),
.B(n_8661),
.Y(n_14958)
);

NAND3xp33_ASAP7_75t_L g14959 ( 
.A(n_14818),
.B(n_14756),
.C(n_14773),
.Y(n_14959)
);

NAND2xp5_ASAP7_75t_L g14960 ( 
.A(n_14778),
.B(n_8661),
.Y(n_14960)
);

OAI22xp33_ASAP7_75t_L g14961 ( 
.A1(n_14744),
.A2(n_8666),
.B1(n_8668),
.B2(n_8662),
.Y(n_14961)
);

NOR2x1_ASAP7_75t_L g14962 ( 
.A(n_14779),
.B(n_8390),
.Y(n_14962)
);

AOI21xp5_ASAP7_75t_L g14963 ( 
.A1(n_14894),
.A2(n_8668),
.B(n_8666),
.Y(n_14963)
);

NAND2xp5_ASAP7_75t_SL g14964 ( 
.A(n_14781),
.B(n_8666),
.Y(n_14964)
);

INVx1_ASAP7_75t_L g14965 ( 
.A(n_14894),
.Y(n_14965)
);

OAI222xp33_ASAP7_75t_L g14966 ( 
.A1(n_14794),
.A2(n_8424),
.B1(n_8391),
.B2(n_8431),
.C1(n_8416),
.C2(n_8403),
.Y(n_14966)
);

AOI211xp5_ASAP7_75t_L g14967 ( 
.A1(n_14783),
.A2(n_8391),
.B(n_8416),
.C(n_8403),
.Y(n_14967)
);

OAI211xp5_ASAP7_75t_SL g14968 ( 
.A1(n_14723),
.A2(n_7336),
.B(n_7672),
.C(n_7417),
.Y(n_14968)
);

AOI21xp5_ASAP7_75t_L g14969 ( 
.A1(n_14814),
.A2(n_8672),
.B(n_8668),
.Y(n_14969)
);

NOR4xp25_ASAP7_75t_L g14970 ( 
.A(n_14890),
.B(n_8766),
.C(n_8761),
.D(n_8431),
.Y(n_14970)
);

AO22x2_ASAP7_75t_L g14971 ( 
.A1(n_14786),
.A2(n_8686),
.B1(n_8687),
.B2(n_8672),
.Y(n_14971)
);

NAND3xp33_ASAP7_75t_L g14972 ( 
.A(n_14799),
.B(n_14802),
.C(n_14800),
.Y(n_14972)
);

AOI21xp5_ASAP7_75t_L g14973 ( 
.A1(n_14841),
.A2(n_8686),
.B(n_8672),
.Y(n_14973)
);

NAND3xp33_ASAP7_75t_SL g14974 ( 
.A(n_14813),
.B(n_6624),
.C(n_6482),
.Y(n_14974)
);

HB1xp67_ASAP7_75t_L g14975 ( 
.A(n_14742),
.Y(n_14975)
);

OAI22xp33_ASAP7_75t_L g14976 ( 
.A1(n_14758),
.A2(n_8687),
.B1(n_8691),
.B2(n_8686),
.Y(n_14976)
);

INVx1_ASAP7_75t_L g14977 ( 
.A(n_14839),
.Y(n_14977)
);

AOI221xp5_ASAP7_75t_L g14978 ( 
.A1(n_14785),
.A2(n_8438),
.B1(n_8442),
.B2(n_8439),
.C(n_8424),
.Y(n_14978)
);

NOR3xp33_ASAP7_75t_L g14979 ( 
.A(n_14816),
.B(n_6624),
.C(n_5251),
.Y(n_14979)
);

OA21x2_ASAP7_75t_L g14980 ( 
.A1(n_14842),
.A2(n_8691),
.B(n_8687),
.Y(n_14980)
);

NAND2xp5_ASAP7_75t_L g14981 ( 
.A(n_14870),
.B(n_8691),
.Y(n_14981)
);

NOR3xp33_ASAP7_75t_L g14982 ( 
.A(n_14775),
.B(n_6624),
.C(n_6363),
.Y(n_14982)
);

NAND3xp33_ASAP7_75t_L g14983 ( 
.A(n_14893),
.B(n_14830),
.C(n_14892),
.Y(n_14983)
);

NOR2x1_ASAP7_75t_L g14984 ( 
.A(n_14831),
.B(n_8439),
.Y(n_14984)
);

AOI21xp33_ASAP7_75t_L g14985 ( 
.A1(n_14844),
.A2(n_14835),
.B(n_14849),
.Y(n_14985)
);

INVx1_ASAP7_75t_L g14986 ( 
.A(n_14797),
.Y(n_14986)
);

AOI21xp5_ASAP7_75t_L g14987 ( 
.A1(n_14832),
.A2(n_8711),
.B(n_8704),
.Y(n_14987)
);

OAI21xp5_ASAP7_75t_L g14988 ( 
.A1(n_14796),
.A2(n_8442),
.B(n_8438),
.Y(n_14988)
);

INVx1_ASAP7_75t_L g14989 ( 
.A(n_14735),
.Y(n_14989)
);

NAND2xp5_ASAP7_75t_L g14990 ( 
.A(n_14771),
.B(n_8704),
.Y(n_14990)
);

INVx1_ASAP7_75t_L g14991 ( 
.A(n_14843),
.Y(n_14991)
);

AOI21xp5_ASAP7_75t_L g14992 ( 
.A1(n_14850),
.A2(n_8711),
.B(n_8704),
.Y(n_14992)
);

OA22x2_ASAP7_75t_L g14993 ( 
.A1(n_14822),
.A2(n_8444),
.B1(n_8446),
.B2(n_8443),
.Y(n_14993)
);

XNOR2x1_ASAP7_75t_SL g14994 ( 
.A(n_14864),
.B(n_6423),
.Y(n_14994)
);

NAND2xp5_ASAP7_75t_SL g14995 ( 
.A(n_14782),
.B(n_8711),
.Y(n_14995)
);

AND2x2_ASAP7_75t_L g14996 ( 
.A(n_14861),
.B(n_8715),
.Y(n_14996)
);

INVx2_ASAP7_75t_L g14997 ( 
.A(n_14906),
.Y(n_14997)
);

OAI211xp5_ASAP7_75t_L g14998 ( 
.A1(n_14867),
.A2(n_8444),
.B(n_8446),
.C(n_8443),
.Y(n_14998)
);

NAND2xp5_ASAP7_75t_L g14999 ( 
.A(n_14868),
.B(n_8715),
.Y(n_14999)
);

NOR2xp33_ASAP7_75t_L g15000 ( 
.A(n_14871),
.B(n_14804),
.Y(n_15000)
);

NAND2xp5_ASAP7_75t_L g15001 ( 
.A(n_14886),
.B(n_8715),
.Y(n_15001)
);

INVx1_ASAP7_75t_L g15002 ( 
.A(n_14737),
.Y(n_15002)
);

HB1xp67_ASAP7_75t_L g15003 ( 
.A(n_14801),
.Y(n_15003)
);

NAND2xp5_ASAP7_75t_L g15004 ( 
.A(n_14776),
.B(n_8723),
.Y(n_15004)
);

NAND3xp33_ASAP7_75t_L g15005 ( 
.A(n_14845),
.B(n_8451),
.C(n_8449),
.Y(n_15005)
);

NAND4xp25_ASAP7_75t_L g15006 ( 
.A(n_14806),
.B(n_6624),
.C(n_6098),
.D(n_7548),
.Y(n_15006)
);

AO22x2_ASAP7_75t_L g15007 ( 
.A1(n_14836),
.A2(n_8724),
.B1(n_8732),
.B2(n_8723),
.Y(n_15007)
);

AOI22xp5_ASAP7_75t_L g15008 ( 
.A1(n_14825),
.A2(n_7527),
.B1(n_8451),
.B2(n_8449),
.Y(n_15008)
);

NOR3xp33_ASAP7_75t_L g15009 ( 
.A(n_14854),
.B(n_5608),
.C(n_5595),
.Y(n_15009)
);

INVxp67_ASAP7_75t_SL g15010 ( 
.A(n_14788),
.Y(n_15010)
);

INVx1_ASAP7_75t_L g15011 ( 
.A(n_14752),
.Y(n_15011)
);

NAND2xp5_ASAP7_75t_L g15012 ( 
.A(n_14878),
.B(n_8724),
.Y(n_15012)
);

NAND2xp5_ASAP7_75t_L g15013 ( 
.A(n_14857),
.B(n_8724),
.Y(n_15013)
);

AOI22xp5_ASAP7_75t_L g15014 ( 
.A1(n_14767),
.A2(n_7527),
.B1(n_8459),
.B2(n_8453),
.Y(n_15014)
);

OAI211xp5_ASAP7_75t_SL g15015 ( 
.A1(n_14895),
.A2(n_7579),
.B(n_7588),
.C(n_7578),
.Y(n_15015)
);

AOI22xp5_ASAP7_75t_L g15016 ( 
.A1(n_14865),
.A2(n_14899),
.B1(n_14810),
.B2(n_14887),
.Y(n_15016)
);

NAND2xp5_ASAP7_75t_L g15017 ( 
.A(n_14884),
.B(n_8732),
.Y(n_15017)
);

INVx1_ASAP7_75t_L g15018 ( 
.A(n_14823),
.Y(n_15018)
);

NAND2xp5_ASAP7_75t_L g15019 ( 
.A(n_14855),
.B(n_8732),
.Y(n_15019)
);

OAI222xp33_ASAP7_75t_L g15020 ( 
.A1(n_14808),
.A2(n_8461),
.B1(n_8459),
.B2(n_8463),
.C1(n_8460),
.C2(n_8453),
.Y(n_15020)
);

NOR2x1_ASAP7_75t_L g15021 ( 
.A(n_14879),
.B(n_8460),
.Y(n_15021)
);

INVx1_ASAP7_75t_L g15022 ( 
.A(n_14889),
.Y(n_15022)
);

OAI22xp5_ASAP7_75t_L g15023 ( 
.A1(n_14885),
.A2(n_8747),
.B1(n_8756),
.B2(n_8736),
.Y(n_15023)
);

NAND4xp75_ASAP7_75t_L g15024 ( 
.A(n_14888),
.B(n_8461),
.C(n_8464),
.D(n_8463),
.Y(n_15024)
);

AOI221xp5_ASAP7_75t_L g15025 ( 
.A1(n_14883),
.A2(n_8478),
.B1(n_8489),
.B2(n_8474),
.C(n_8464),
.Y(n_15025)
);

NAND3xp33_ASAP7_75t_L g15026 ( 
.A(n_14738),
.B(n_8478),
.C(n_8474),
.Y(n_15026)
);

NOR3x1_ASAP7_75t_L g15027 ( 
.A(n_14882),
.B(n_8494),
.C(n_8489),
.Y(n_15027)
);

AOI21xp5_ASAP7_75t_L g15028 ( 
.A1(n_14897),
.A2(n_8747),
.B(n_8736),
.Y(n_15028)
);

AO22x2_ASAP7_75t_SL g15029 ( 
.A1(n_14750),
.A2(n_8747),
.B1(n_8756),
.B2(n_8736),
.Y(n_15029)
);

NOR3xp33_ASAP7_75t_L g15030 ( 
.A(n_14833),
.B(n_5608),
.C(n_5595),
.Y(n_15030)
);

OAI21xp33_ASAP7_75t_L g15031 ( 
.A1(n_14862),
.A2(n_8504),
.B(n_8494),
.Y(n_15031)
);

NAND4xp25_ASAP7_75t_SL g15032 ( 
.A(n_14881),
.B(n_8505),
.C(n_8514),
.D(n_8504),
.Y(n_15032)
);

NAND2xp5_ASAP7_75t_SL g15033 ( 
.A(n_14852),
.B(n_8756),
.Y(n_15033)
);

INVx1_ASAP7_75t_L g15034 ( 
.A(n_14897),
.Y(n_15034)
);

INVx1_ASAP7_75t_L g15035 ( 
.A(n_14903),
.Y(n_15035)
);

AOI21xp5_ASAP7_75t_L g15036 ( 
.A1(n_14903),
.A2(n_8765),
.B(n_8763),
.Y(n_15036)
);

AOI221xp5_ASAP7_75t_L g15037 ( 
.A1(n_14873),
.A2(n_8515),
.B1(n_8518),
.B2(n_8514),
.C(n_8505),
.Y(n_15037)
);

OAI21xp5_ASAP7_75t_L g15038 ( 
.A1(n_14847),
.A2(n_8518),
.B(n_8515),
.Y(n_15038)
);

INVx1_ASAP7_75t_L g15039 ( 
.A(n_14784),
.Y(n_15039)
);

AOI31xp33_ASAP7_75t_L g15040 ( 
.A1(n_14880),
.A2(n_6440),
.A3(n_6423),
.B(n_6406),
.Y(n_15040)
);

AOI22xp5_ASAP7_75t_L g15041 ( 
.A1(n_14826),
.A2(n_8533),
.B1(n_8536),
.B2(n_8535),
.Y(n_15041)
);

NAND2xp5_ASAP7_75t_L g15042 ( 
.A(n_14811),
.B(n_8763),
.Y(n_15042)
);

NOR2x1_ASAP7_75t_L g15043 ( 
.A(n_14761),
.B(n_8533),
.Y(n_15043)
);

NAND2xp5_ASAP7_75t_L g15044 ( 
.A(n_14876),
.B(n_8765),
.Y(n_15044)
);

INVx2_ASAP7_75t_SL g15045 ( 
.A(n_14784),
.Y(n_15045)
);

AND2x2_ASAP7_75t_L g15046 ( 
.A(n_14848),
.B(n_8765),
.Y(n_15046)
);

OAI21xp33_ASAP7_75t_L g15047 ( 
.A1(n_14766),
.A2(n_8536),
.B(n_8535),
.Y(n_15047)
);

NOR3x1_ASAP7_75t_L g15048 ( 
.A(n_14728),
.B(n_8539),
.C(n_8538),
.Y(n_15048)
);

AOI21xp5_ASAP7_75t_L g15049 ( 
.A1(n_14872),
.A2(n_8769),
.B(n_8768),
.Y(n_15049)
);

NOR3x1_ASAP7_75t_L g15050 ( 
.A(n_14743),
.B(n_8539),
.C(n_8538),
.Y(n_15050)
);

AO22x2_ASAP7_75t_L g15051 ( 
.A1(n_14793),
.A2(n_8769),
.B1(n_8772),
.B2(n_8768),
.Y(n_15051)
);

OA22x2_ASAP7_75t_L g15052 ( 
.A1(n_14762),
.A2(n_8553),
.B1(n_8555),
.B2(n_8548),
.Y(n_15052)
);

NAND2xp5_ASAP7_75t_L g15053 ( 
.A(n_14840),
.B(n_8768),
.Y(n_15053)
);

AOI21xp5_ASAP7_75t_L g15054 ( 
.A1(n_14875),
.A2(n_8772),
.B(n_8769),
.Y(n_15054)
);

NAND2xp5_ASAP7_75t_SL g15055 ( 
.A(n_14746),
.B(n_8772),
.Y(n_15055)
);

INVx1_ASAP7_75t_L g15056 ( 
.A(n_14866),
.Y(n_15056)
);

AOI21xp5_ASAP7_75t_L g15057 ( 
.A1(n_14795),
.A2(n_8780),
.B(n_8776),
.Y(n_15057)
);

OAI21x1_ASAP7_75t_SL g15058 ( 
.A1(n_14874),
.A2(n_8787),
.B(n_8780),
.Y(n_15058)
);

INVx1_ASAP7_75t_L g15059 ( 
.A(n_14866),
.Y(n_15059)
);

AND2x2_ASAP7_75t_L g15060 ( 
.A(n_14763),
.B(n_8776),
.Y(n_15060)
);

AOI211x1_ASAP7_75t_L g15061 ( 
.A1(n_14856),
.A2(n_8548),
.B(n_8555),
.C(n_8553),
.Y(n_15061)
);

NOR3xp33_ASAP7_75t_L g15062 ( 
.A(n_14972),
.B(n_14821),
.C(n_14790),
.Y(n_15062)
);

INVx1_ASAP7_75t_L g15063 ( 
.A(n_14975),
.Y(n_15063)
);

NOR3xp33_ASAP7_75t_L g15064 ( 
.A(n_14912),
.B(n_14819),
.C(n_14901),
.Y(n_15064)
);

NAND3xp33_ASAP7_75t_SL g15065 ( 
.A(n_14922),
.B(n_14824),
.C(n_14858),
.Y(n_15065)
);

AOI21xp5_ASAP7_75t_L g15066 ( 
.A1(n_14908),
.A2(n_14860),
.B(n_14812),
.Y(n_15066)
);

AOI22xp5_ASAP7_75t_L g15067 ( 
.A1(n_14919),
.A2(n_14765),
.B1(n_14729),
.B2(n_14798),
.Y(n_15067)
);

NAND2xp5_ASAP7_75t_L g15068 ( 
.A(n_14920),
.B(n_14891),
.Y(n_15068)
);

INVx1_ASAP7_75t_L g15069 ( 
.A(n_14945),
.Y(n_15069)
);

NAND3xp33_ASAP7_75t_L g15070 ( 
.A(n_14955),
.B(n_14859),
.C(n_14853),
.Y(n_15070)
);

INVx1_ASAP7_75t_L g15071 ( 
.A(n_14956),
.Y(n_15071)
);

OAI22x1_ASAP7_75t_L g15072 ( 
.A1(n_14941),
.A2(n_14851),
.B1(n_8599),
.B2(n_8633),
.Y(n_15072)
);

NOR3xp33_ASAP7_75t_L g15073 ( 
.A(n_14959),
.B(n_5608),
.C(n_5595),
.Y(n_15073)
);

NAND2xp5_ASAP7_75t_L g15074 ( 
.A(n_14957),
.B(n_8776),
.Y(n_15074)
);

NOR2xp33_ASAP7_75t_L g15075 ( 
.A(n_14913),
.B(n_6642),
.Y(n_15075)
);

AOI22x1_ASAP7_75t_L g15076 ( 
.A1(n_14965),
.A2(n_8567),
.B1(n_8568),
.B2(n_8556),
.Y(n_15076)
);

NOR2xp33_ASAP7_75t_L g15077 ( 
.A(n_14977),
.B(n_6642),
.Y(n_15077)
);

XOR2xp5_ASAP7_75t_L g15078 ( 
.A(n_14983),
.B(n_7600),
.Y(n_15078)
);

AOI221xp5_ASAP7_75t_L g15079 ( 
.A1(n_14924),
.A2(n_8728),
.B1(n_8568),
.B2(n_8571),
.C(n_8567),
.Y(n_15079)
);

NOR3x1_ASAP7_75t_L g15080 ( 
.A(n_15010),
.B(n_8571),
.C(n_8556),
.Y(n_15080)
);

NOR2xp67_ASAP7_75t_L g15081 ( 
.A(n_14942),
.B(n_8572),
.Y(n_15081)
);

INVx1_ASAP7_75t_L g15082 ( 
.A(n_14936),
.Y(n_15082)
);

NAND2xp5_ASAP7_75t_L g15083 ( 
.A(n_14926),
.B(n_8780),
.Y(n_15083)
);

NOR2xp67_ASAP7_75t_L g15084 ( 
.A(n_14921),
.B(n_8572),
.Y(n_15084)
);

OAI211xp5_ASAP7_75t_L g15085 ( 
.A1(n_14985),
.A2(n_15003),
.B(n_14989),
.C(n_14986),
.Y(n_15085)
);

INVxp67_ASAP7_75t_L g15086 ( 
.A(n_15000),
.Y(n_15086)
);

AOI211xp5_ASAP7_75t_L g15087 ( 
.A1(n_14991),
.A2(n_15002),
.B(n_15011),
.C(n_15018),
.Y(n_15087)
);

NAND2xp5_ASAP7_75t_L g15088 ( 
.A(n_14930),
.B(n_8783),
.Y(n_15088)
);

NAND2xp5_ASAP7_75t_L g15089 ( 
.A(n_14944),
.B(n_8783),
.Y(n_15089)
);

AOI21xp33_ASAP7_75t_SL g15090 ( 
.A1(n_15022),
.A2(n_14997),
.B(n_15045),
.Y(n_15090)
);

INVxp67_ASAP7_75t_SL g15091 ( 
.A(n_14994),
.Y(n_15091)
);

NOR2xp33_ASAP7_75t_L g15092 ( 
.A(n_14910),
.B(n_6642),
.Y(n_15092)
);

AOI211x1_ASAP7_75t_L g15093 ( 
.A1(n_15055),
.A2(n_8573),
.B(n_8575),
.C(n_8574),
.Y(n_15093)
);

NOR4xp75_ASAP7_75t_L g15094 ( 
.A(n_14907),
.B(n_6044),
.C(n_6045),
.D(n_6026),
.Y(n_15094)
);

NAND4xp75_ASAP7_75t_L g15095 ( 
.A(n_15034),
.B(n_8573),
.C(n_8575),
.D(n_8574),
.Y(n_15095)
);

INVx1_ASAP7_75t_L g15096 ( 
.A(n_14911),
.Y(n_15096)
);

NAND4xp75_ASAP7_75t_L g15097 ( 
.A(n_15035),
.B(n_8578),
.C(n_8583),
.D(n_8582),
.Y(n_15097)
);

NOR2xp33_ASAP7_75t_L g15098 ( 
.A(n_14946),
.B(n_6642),
.Y(n_15098)
);

NOR3x1_ASAP7_75t_L g15099 ( 
.A(n_14914),
.B(n_8582),
.C(n_8578),
.Y(n_15099)
);

NOR3x1_ASAP7_75t_L g15100 ( 
.A(n_14933),
.B(n_8588),
.C(n_8583),
.Y(n_15100)
);

NAND3xp33_ASAP7_75t_L g15101 ( 
.A(n_15016),
.B(n_8590),
.C(n_8588),
.Y(n_15101)
);

NOR3xp33_ASAP7_75t_SL g15102 ( 
.A(n_15039),
.B(n_15059),
.C(n_15056),
.Y(n_15102)
);

INVx1_ASAP7_75t_L g15103 ( 
.A(n_14962),
.Y(n_15103)
);

NOR2x1_ASAP7_75t_L g15104 ( 
.A(n_14932),
.B(n_8590),
.Y(n_15104)
);

AOI21xp5_ASAP7_75t_L g15105 ( 
.A1(n_14937),
.A2(n_8787),
.B(n_8784),
.Y(n_15105)
);

INVx2_ASAP7_75t_L g15106 ( 
.A(n_14915),
.Y(n_15106)
);

NAND2xp5_ASAP7_75t_L g15107 ( 
.A(n_14925),
.B(n_8784),
.Y(n_15107)
);

NOR2xp67_ASAP7_75t_L g15108 ( 
.A(n_14949),
.B(n_8805),
.Y(n_15108)
);

AOI211xp5_ASAP7_75t_L g15109 ( 
.A1(n_14935),
.A2(n_8599),
.B(n_8605),
.C(n_8594),
.Y(n_15109)
);

INVx1_ASAP7_75t_L g15110 ( 
.A(n_14954),
.Y(n_15110)
);

AND4x1_ASAP7_75t_L g15111 ( 
.A(n_14917),
.B(n_7602),
.C(n_7657),
.D(n_7642),
.Y(n_15111)
);

AND5x1_ASAP7_75t_L g15112 ( 
.A(n_14939),
.B(n_15030),
.C(n_14963),
.D(n_15009),
.E(n_15014),
.Y(n_15112)
);

NOR2x1p5_ASAP7_75t_L g15113 ( 
.A(n_14943),
.B(n_6406),
.Y(n_15113)
);

AND3x1_ASAP7_75t_L g15114 ( 
.A(n_14918),
.B(n_8597),
.C(n_8594),
.Y(n_15114)
);

OA22x2_ASAP7_75t_L g15115 ( 
.A1(n_14964),
.A2(n_8810),
.B1(n_8605),
.B2(n_8611),
.Y(n_15115)
);

INVx1_ASAP7_75t_L g15116 ( 
.A(n_14984),
.Y(n_15116)
);

NAND2xp5_ASAP7_75t_L g15117 ( 
.A(n_15060),
.B(n_8810),
.Y(n_15117)
);

NAND3xp33_ASAP7_75t_SL g15118 ( 
.A(n_14981),
.B(n_14999),
.C(n_14960),
.Y(n_15118)
);

AND2x2_ASAP7_75t_L g15119 ( 
.A(n_15046),
.B(n_6614),
.Y(n_15119)
);

AND4x1_ASAP7_75t_L g15120 ( 
.A(n_15048),
.B(n_7789),
.C(n_7770),
.D(n_7665),
.Y(n_15120)
);

INVx1_ASAP7_75t_SL g15121 ( 
.A(n_14958),
.Y(n_15121)
);

NOR2x1_ASAP7_75t_L g15122 ( 
.A(n_15043),
.B(n_8597),
.Y(n_15122)
);

NOR2xp33_ASAP7_75t_L g15123 ( 
.A(n_15042),
.B(n_6642),
.Y(n_15123)
);

NOR2x1_ASAP7_75t_L g15124 ( 
.A(n_14951),
.B(n_8611),
.Y(n_15124)
);

NAND2xp5_ASAP7_75t_L g15125 ( 
.A(n_14996),
.B(n_8613),
.Y(n_15125)
);

NAND2xp5_ASAP7_75t_L g15126 ( 
.A(n_15061),
.B(n_8613),
.Y(n_15126)
);

INVx1_ASAP7_75t_L g15127 ( 
.A(n_15027),
.Y(n_15127)
);

OAI322xp33_ASAP7_75t_L g15128 ( 
.A1(n_15013),
.A2(n_8632),
.A3(n_8622),
.B1(n_8633),
.B2(n_8635),
.C1(n_8630),
.C2(n_8620),
.Y(n_15128)
);

NOR2x1_ASAP7_75t_SL g15129 ( 
.A(n_14974),
.B(n_8620),
.Y(n_15129)
);

NAND3xp33_ASAP7_75t_L g15130 ( 
.A(n_14995),
.B(n_8630),
.C(n_8622),
.Y(n_15130)
);

NAND3xp33_ASAP7_75t_SL g15131 ( 
.A(n_15012),
.B(n_8738),
.C(n_8728),
.Y(n_15131)
);

NOR2x1_ASAP7_75t_L g15132 ( 
.A(n_15021),
.B(n_8632),
.Y(n_15132)
);

NAND3xp33_ASAP7_75t_L g15133 ( 
.A(n_15019),
.B(n_8636),
.C(n_8635),
.Y(n_15133)
);

NOR3xp33_ASAP7_75t_L g15134 ( 
.A(n_14990),
.B(n_5608),
.C(n_5595),
.Y(n_15134)
);

AOI211x1_ASAP7_75t_L g15135 ( 
.A1(n_14923),
.A2(n_8636),
.B(n_8641),
.C(n_8639),
.Y(n_15135)
);

NAND3xp33_ASAP7_75t_L g15136 ( 
.A(n_15033),
.B(n_8641),
.C(n_8639),
.Y(n_15136)
);

NAND3xp33_ASAP7_75t_L g15137 ( 
.A(n_14982),
.B(n_8644),
.C(n_8642),
.Y(n_15137)
);

OAI21xp5_ASAP7_75t_L g15138 ( 
.A1(n_14909),
.A2(n_8644),
.B(n_8642),
.Y(n_15138)
);

AOI211xp5_ASAP7_75t_L g15139 ( 
.A1(n_15032),
.A2(n_8664),
.B(n_8665),
.C(n_8649),
.Y(n_15139)
);

INVx1_ASAP7_75t_L g15140 ( 
.A(n_14916),
.Y(n_15140)
);

AND5x1_ASAP7_75t_L g15141 ( 
.A(n_14952),
.B(n_14938),
.C(n_14979),
.D(n_15008),
.E(n_14969),
.Y(n_15141)
);

AOI211xp5_ASAP7_75t_SL g15142 ( 
.A1(n_14961),
.A2(n_8654),
.B(n_8664),
.C(n_8649),
.Y(n_15142)
);

NOR2x1_ASAP7_75t_L g15143 ( 
.A(n_15017),
.B(n_8654),
.Y(n_15143)
);

OAI211xp5_ASAP7_75t_SL g15144 ( 
.A1(n_15004),
.A2(n_7772),
.B(n_7668),
.C(n_7774),
.Y(n_15144)
);

NAND2xp5_ASAP7_75t_L g15145 ( 
.A(n_15050),
.B(n_8665),
.Y(n_15145)
);

AND3x4_ASAP7_75t_L g15146 ( 
.A(n_14934),
.B(n_6535),
.C(n_6530),
.Y(n_15146)
);

NOR2xp33_ASAP7_75t_L g15147 ( 
.A(n_15044),
.B(n_8667),
.Y(n_15147)
);

NOR3xp33_ASAP7_75t_L g15148 ( 
.A(n_15006),
.B(n_5608),
.C(n_5595),
.Y(n_15148)
);

INVx1_ASAP7_75t_L g15149 ( 
.A(n_15029),
.Y(n_15149)
);

NAND2xp5_ASAP7_75t_L g15150 ( 
.A(n_14950),
.B(n_8667),
.Y(n_15150)
);

INVxp67_ASAP7_75t_SL g15151 ( 
.A(n_15053),
.Y(n_15151)
);

INVx2_ASAP7_75t_L g15152 ( 
.A(n_15007),
.Y(n_15152)
);

AOI22xp5_ASAP7_75t_L g15153 ( 
.A1(n_14928),
.A2(n_8682),
.B1(n_8683),
.B2(n_8670),
.Y(n_15153)
);

INVxp33_ASAP7_75t_L g15154 ( 
.A(n_15001),
.Y(n_15154)
);

AOI22xp5_ASAP7_75t_L g15155 ( 
.A1(n_14993),
.A2(n_8682),
.B1(n_8683),
.B2(n_8670),
.Y(n_15155)
);

NOR3xp33_ASAP7_75t_L g15156 ( 
.A(n_15024),
.B(n_5700),
.C(n_5677),
.Y(n_15156)
);

OA22x2_ASAP7_75t_L g15157 ( 
.A1(n_14988),
.A2(n_14948),
.B1(n_14947),
.B2(n_15038),
.Y(n_15157)
);

NOR2x1p5_ASAP7_75t_L g15158 ( 
.A(n_15026),
.B(n_6021),
.Y(n_15158)
);

AND4x1_ASAP7_75t_L g15159 ( 
.A(n_14970),
.B(n_6393),
.C(n_6437),
.D(n_6293),
.Y(n_15159)
);

INVx1_ASAP7_75t_L g15160 ( 
.A(n_15052),
.Y(n_15160)
);

NAND5xp2_ASAP7_75t_L g15161 ( 
.A(n_14940),
.B(n_5900),
.C(n_5943),
.D(n_5884),
.E(n_5861),
.Y(n_15161)
);

NOR3x1_ASAP7_75t_L g15162 ( 
.A(n_15005),
.B(n_8689),
.C(n_8684),
.Y(n_15162)
);

NAND2xp5_ASAP7_75t_L g15163 ( 
.A(n_15031),
.B(n_8684),
.Y(n_15163)
);

NOR3xp33_ASAP7_75t_L g15164 ( 
.A(n_14966),
.B(n_5700),
.C(n_5677),
.Y(n_15164)
);

NAND3xp33_ASAP7_75t_L g15165 ( 
.A(n_14927),
.B(n_8692),
.C(n_8689),
.Y(n_15165)
);

CKINVDCx6p67_ASAP7_75t_R g15166 ( 
.A(n_15040),
.Y(n_15166)
);

INVxp67_ASAP7_75t_L g15167 ( 
.A(n_15007),
.Y(n_15167)
);

INVx1_ASAP7_75t_L g15168 ( 
.A(n_15051),
.Y(n_15168)
);

NOR3xp33_ASAP7_75t_L g15169 ( 
.A(n_14976),
.B(n_14968),
.C(n_15047),
.Y(n_15169)
);

NOR2xp33_ASAP7_75t_L g15170 ( 
.A(n_14998),
.B(n_8692),
.Y(n_15170)
);

NOR3x1_ASAP7_75t_L g15171 ( 
.A(n_15023),
.B(n_8700),
.C(n_8695),
.Y(n_15171)
);

INVx2_ASAP7_75t_L g15172 ( 
.A(n_15051),
.Y(n_15172)
);

INVx1_ASAP7_75t_L g15173 ( 
.A(n_14980),
.Y(n_15173)
);

NOR2xp33_ASAP7_75t_L g15174 ( 
.A(n_15020),
.B(n_8695),
.Y(n_15174)
);

NOR3xp33_ASAP7_75t_L g15175 ( 
.A(n_14953),
.B(n_5700),
.C(n_5677),
.Y(n_15175)
);

AND3x2_ASAP7_75t_L g15176 ( 
.A(n_14967),
.B(n_6220),
.C(n_8700),
.Y(n_15176)
);

NAND2xp5_ASAP7_75t_SL g15177 ( 
.A(n_14973),
.B(n_8703),
.Y(n_15177)
);

XNOR2x1_ASAP7_75t_SL g15178 ( 
.A(n_14931),
.B(n_6423),
.Y(n_15178)
);

NOR2x1_ASAP7_75t_L g15179 ( 
.A(n_14980),
.B(n_8703),
.Y(n_15179)
);

OAI211xp5_ASAP7_75t_L g15180 ( 
.A1(n_14987),
.A2(n_8716),
.B(n_8717),
.C(n_8709),
.Y(n_15180)
);

OAI222xp33_ASAP7_75t_R g15181 ( 
.A1(n_15057),
.A2(n_5869),
.B1(n_5820),
.B2(n_5937),
.C1(n_5842),
.C2(n_5791),
.Y(n_15181)
);

NAND4xp25_ASAP7_75t_SL g15182 ( 
.A(n_14992),
.B(n_8709),
.C(n_8717),
.D(n_8716),
.Y(n_15182)
);

INVx1_ASAP7_75t_L g15183 ( 
.A(n_15058),
.Y(n_15183)
);

NOR3xp33_ASAP7_75t_L g15184 ( 
.A(n_15015),
.B(n_5700),
.C(n_5677),
.Y(n_15184)
);

NAND3xp33_ASAP7_75t_L g15185 ( 
.A(n_14929),
.B(n_8738),
.C(n_8720),
.Y(n_15185)
);

INVxp67_ASAP7_75t_SL g15186 ( 
.A(n_15028),
.Y(n_15186)
);

NAND5xp2_ASAP7_75t_L g15187 ( 
.A(n_15054),
.B(n_15049),
.C(n_15036),
.D(n_14978),
.E(n_15041),
.Y(n_15187)
);

OAI322xp33_ASAP7_75t_L g15188 ( 
.A1(n_14931),
.A2(n_8744),
.A3(n_8739),
.B1(n_8750),
.B2(n_8759),
.C1(n_8740),
.C2(n_8720),
.Y(n_15188)
);

AOI22xp5_ASAP7_75t_L g15189 ( 
.A1(n_14971),
.A2(n_8740),
.B1(n_8744),
.B2(n_8739),
.Y(n_15189)
);

INVx2_ASAP7_75t_L g15190 ( 
.A(n_14971),
.Y(n_15190)
);

AND4x1_ASAP7_75t_L g15191 ( 
.A(n_15037),
.B(n_6393),
.C(n_6437),
.D(n_6293),
.Y(n_15191)
);

NOR2x1_ASAP7_75t_L g15192 ( 
.A(n_15025),
.B(n_8750),
.Y(n_15192)
);

BUFx6f_ASAP7_75t_L g15193 ( 
.A(n_15069),
.Y(n_15193)
);

NAND3xp33_ASAP7_75t_L g15194 ( 
.A(n_15087),
.B(n_8761),
.C(n_8759),
.Y(n_15194)
);

NAND2xp5_ASAP7_75t_L g15195 ( 
.A(n_15063),
.B(n_7418),
.Y(n_15195)
);

NOR3x1_ASAP7_75t_L g15196 ( 
.A(n_15085),
.B(n_15070),
.C(n_15065),
.Y(n_15196)
);

OAI22xp5_ASAP7_75t_L g15197 ( 
.A1(n_15071),
.A2(n_7232),
.B1(n_7241),
.B2(n_7224),
.Y(n_15197)
);

AOI211xp5_ASAP7_75t_SL g15198 ( 
.A1(n_15086),
.A2(n_15082),
.B(n_15066),
.C(n_15068),
.Y(n_15198)
);

NAND2xp5_ASAP7_75t_L g15199 ( 
.A(n_15077),
.B(n_15091),
.Y(n_15199)
);

OAI211xp5_ASAP7_75t_SL g15200 ( 
.A1(n_15102),
.A2(n_6044),
.B(n_6063),
.C(n_6045),
.Y(n_15200)
);

NAND4xp25_ASAP7_75t_L g15201 ( 
.A(n_15062),
.B(n_5813),
.C(n_5799),
.D(n_6063),
.Y(n_15201)
);

NOR2x1_ASAP7_75t_L g15202 ( 
.A(n_15110),
.B(n_6530),
.Y(n_15202)
);

AOI22xp33_ASAP7_75t_L g15203 ( 
.A1(n_15148),
.A2(n_7769),
.B1(n_7338),
.B2(n_7570),
.Y(n_15203)
);

INVx1_ASAP7_75t_L g15204 ( 
.A(n_15078),
.Y(n_15204)
);

OR2x2_ASAP7_75t_L g15205 ( 
.A(n_15096),
.B(n_6021),
.Y(n_15205)
);

NOR3x1_ASAP7_75t_L g15206 ( 
.A(n_15140),
.B(n_6075),
.C(n_5983),
.Y(n_15206)
);

NAND4xp25_ASAP7_75t_L g15207 ( 
.A(n_15080),
.B(n_6075),
.C(n_5855),
.D(n_5856),
.Y(n_15207)
);

NOR3xp33_ASAP7_75t_L g15208 ( 
.A(n_15090),
.B(n_5700),
.C(n_5677),
.Y(n_15208)
);

NOR4xp25_ASAP7_75t_L g15209 ( 
.A(n_15149),
.B(n_7744),
.C(n_7746),
.D(n_7737),
.Y(n_15209)
);

INVxp33_ASAP7_75t_L g15210 ( 
.A(n_15064),
.Y(n_15210)
);

AND2x2_ASAP7_75t_L g15211 ( 
.A(n_15119),
.B(n_6614),
.Y(n_15211)
);

NOR4xp25_ASAP7_75t_L g15212 ( 
.A(n_15118),
.B(n_7746),
.C(n_7753),
.D(n_7744),
.Y(n_15212)
);

NOR2x1_ASAP7_75t_L g15213 ( 
.A(n_15103),
.B(n_6530),
.Y(n_15213)
);

NOR2x1_ASAP7_75t_L g15214 ( 
.A(n_15173),
.B(n_6530),
.Y(n_15214)
);

NAND2xp5_ASAP7_75t_SL g15215 ( 
.A(n_15106),
.B(n_7338),
.Y(n_15215)
);

NOR3xp33_ASAP7_75t_L g15216 ( 
.A(n_15127),
.B(n_5707),
.C(n_5700),
.Y(n_15216)
);

INVx1_ASAP7_75t_L g15217 ( 
.A(n_15074),
.Y(n_15217)
);

NAND3xp33_ASAP7_75t_L g15218 ( 
.A(n_15160),
.B(n_6390),
.C(n_6334),
.Y(n_15218)
);

NOR3xp33_ASAP7_75t_L g15219 ( 
.A(n_15151),
.B(n_5735),
.C(n_5707),
.Y(n_15219)
);

NOR2x1_ASAP7_75t_L g15220 ( 
.A(n_15116),
.B(n_15190),
.Y(n_15220)
);

NAND2xp5_ASAP7_75t_L g15221 ( 
.A(n_15123),
.B(n_15075),
.Y(n_15221)
);

AND4x1_ASAP7_75t_L g15222 ( 
.A(n_15183),
.B(n_6168),
.C(n_6173),
.D(n_5815),
.Y(n_15222)
);

INVx1_ASAP7_75t_L g15223 ( 
.A(n_15081),
.Y(n_15223)
);

NOR3x1_ASAP7_75t_L g15224 ( 
.A(n_15186),
.B(n_5983),
.C(n_5976),
.Y(n_15224)
);

NAND3xp33_ASAP7_75t_L g15225 ( 
.A(n_15167),
.B(n_6390),
.C(n_6334),
.Y(n_15225)
);

NAND2xp5_ASAP7_75t_L g15226 ( 
.A(n_15098),
.B(n_7418),
.Y(n_15226)
);

NAND2xp5_ASAP7_75t_SL g15227 ( 
.A(n_15067),
.B(n_7338),
.Y(n_15227)
);

NOR3x1_ASAP7_75t_L g15228 ( 
.A(n_15168),
.B(n_5976),
.C(n_5942),
.Y(n_15228)
);

NAND3xp33_ASAP7_75t_SL g15229 ( 
.A(n_15121),
.B(n_5964),
.C(n_5150),
.Y(n_15229)
);

XOR2x1_ASAP7_75t_L g15230 ( 
.A(n_15152),
.B(n_6440),
.Y(n_15230)
);

NOR3xp33_ASAP7_75t_L g15231 ( 
.A(n_15187),
.B(n_5735),
.C(n_5707),
.Y(n_15231)
);

NAND3xp33_ASAP7_75t_L g15232 ( 
.A(n_15169),
.B(n_6429),
.C(n_6395),
.Y(n_15232)
);

NOR2x1_ASAP7_75t_L g15233 ( 
.A(n_15172),
.B(n_15084),
.Y(n_15233)
);

NAND2xp5_ASAP7_75t_L g15234 ( 
.A(n_15176),
.B(n_7418),
.Y(n_15234)
);

NOR3xp33_ASAP7_75t_L g15235 ( 
.A(n_15092),
.B(n_5735),
.C(n_5707),
.Y(n_15235)
);

AND2x4_ASAP7_75t_L g15236 ( 
.A(n_15112),
.B(n_7141),
.Y(n_15236)
);

AND4x1_ASAP7_75t_L g15237 ( 
.A(n_15122),
.B(n_6173),
.C(n_5815),
.D(n_5827),
.Y(n_15237)
);

NOR3xp33_ASAP7_75t_L g15238 ( 
.A(n_15154),
.B(n_5735),
.C(n_5707),
.Y(n_15238)
);

NOR2x1_ASAP7_75t_L g15239 ( 
.A(n_15104),
.B(n_6530),
.Y(n_15239)
);

AOI22xp5_ASAP7_75t_L g15240 ( 
.A1(n_15166),
.A2(n_6535),
.B1(n_6568),
.B2(n_6549),
.Y(n_15240)
);

NAND3xp33_ASAP7_75t_SL g15241 ( 
.A(n_15117),
.B(n_5964),
.C(n_5150),
.Y(n_15241)
);

NOR3xp33_ASAP7_75t_L g15242 ( 
.A(n_15083),
.B(n_5735),
.C(n_5707),
.Y(n_15242)
);

NOR4xp25_ASAP7_75t_L g15243 ( 
.A(n_15145),
.B(n_7753),
.C(n_7763),
.D(n_7755),
.Y(n_15243)
);

NOR3xp33_ASAP7_75t_L g15244 ( 
.A(n_15088),
.B(n_5739),
.C(n_5735),
.Y(n_15244)
);

AND2x2_ASAP7_75t_L g15245 ( 
.A(n_15113),
.B(n_6614),
.Y(n_15245)
);

NOR3xp33_ASAP7_75t_L g15246 ( 
.A(n_15147),
.B(n_15134),
.C(n_15073),
.Y(n_15246)
);

NOR2x1_ASAP7_75t_L g15247 ( 
.A(n_15124),
.B(n_6535),
.Y(n_15247)
);

NOR3xp33_ASAP7_75t_L g15248 ( 
.A(n_15126),
.B(n_5739),
.C(n_5100),
.Y(n_15248)
);

AND4x1_ASAP7_75t_L g15249 ( 
.A(n_15143),
.B(n_5827),
.C(n_5855),
.D(n_5851),
.Y(n_15249)
);

OAI21xp33_ASAP7_75t_L g15250 ( 
.A1(n_15157),
.A2(n_6549),
.B(n_6535),
.Y(n_15250)
);

NOR3xp33_ASAP7_75t_L g15251 ( 
.A(n_15150),
.B(n_5739),
.C(n_5851),
.Y(n_15251)
);

NAND2xp5_ASAP7_75t_L g15252 ( 
.A(n_15174),
.B(n_7465),
.Y(n_15252)
);

NOR2x1_ASAP7_75t_L g15253 ( 
.A(n_15132),
.B(n_6535),
.Y(n_15253)
);

AOI221x1_ASAP7_75t_L g15254 ( 
.A1(n_15072),
.A2(n_7224),
.B1(n_7255),
.B2(n_7241),
.C(n_7232),
.Y(n_15254)
);

NAND4xp25_ASAP7_75t_L g15255 ( 
.A(n_15162),
.B(n_5856),
.C(n_5871),
.D(n_5864),
.Y(n_15255)
);

NAND4xp25_ASAP7_75t_L g15256 ( 
.A(n_15093),
.B(n_15175),
.C(n_15171),
.D(n_15101),
.Y(n_15256)
);

INVx1_ASAP7_75t_L g15257 ( 
.A(n_15178),
.Y(n_15257)
);

NOR3xp33_ASAP7_75t_SL g15258 ( 
.A(n_15170),
.B(n_5871),
.C(n_5864),
.Y(n_15258)
);

NOR2x1_ASAP7_75t_L g15259 ( 
.A(n_15179),
.B(n_6549),
.Y(n_15259)
);

NAND4xp75_ASAP7_75t_L g15260 ( 
.A(n_15114),
.B(n_6317),
.C(n_5546),
.D(n_5942),
.Y(n_15260)
);

AND3x2_ASAP7_75t_L g15261 ( 
.A(n_15164),
.B(n_6220),
.C(n_6395),
.Y(n_15261)
);

OA22x2_ASAP7_75t_SL g15262 ( 
.A1(n_15181),
.A2(n_7255),
.B1(n_7261),
.B2(n_7241),
.Y(n_15262)
);

INVx2_ASAP7_75t_SL g15263 ( 
.A(n_15115),
.Y(n_15263)
);

NOR2x1p5_ASAP7_75t_L g15264 ( 
.A(n_15163),
.B(n_6417),
.Y(n_15264)
);

NOR3x1_ASAP7_75t_L g15265 ( 
.A(n_15125),
.B(n_5944),
.C(n_5928),
.Y(n_15265)
);

NOR2x1_ASAP7_75t_L g15266 ( 
.A(n_15108),
.B(n_6549),
.Y(n_15266)
);

NOR3xp33_ASAP7_75t_L g15267 ( 
.A(n_15141),
.B(n_5739),
.C(n_5876),
.Y(n_15267)
);

INVx2_ASAP7_75t_L g15268 ( 
.A(n_15095),
.Y(n_15268)
);

NOR4xp25_ASAP7_75t_L g15269 ( 
.A(n_15177),
.B(n_7755),
.C(n_7766),
.D(n_7763),
.Y(n_15269)
);

NOR2xp33_ASAP7_75t_SL g15270 ( 
.A(n_15108),
.B(n_7343),
.Y(n_15270)
);

INVx1_ASAP7_75t_L g15271 ( 
.A(n_15129),
.Y(n_15271)
);

INVx1_ASAP7_75t_L g15272 ( 
.A(n_15192),
.Y(n_15272)
);

AND2x2_ASAP7_75t_L g15273 ( 
.A(n_15158),
.B(n_6614),
.Y(n_15273)
);

NOR3xp33_ASAP7_75t_L g15274 ( 
.A(n_15107),
.B(n_5739),
.C(n_5876),
.Y(n_15274)
);

NOR2x1_ASAP7_75t_L g15275 ( 
.A(n_15097),
.B(n_6549),
.Y(n_15275)
);

NOR3x1_ASAP7_75t_L g15276 ( 
.A(n_15089),
.B(n_5944),
.C(n_5928),
.Y(n_15276)
);

NOR3xp33_ASAP7_75t_L g15277 ( 
.A(n_15131),
.B(n_5739),
.C(n_5950),
.Y(n_15277)
);

NOR2xp33_ASAP7_75t_L g15278 ( 
.A(n_15146),
.B(n_7343),
.Y(n_15278)
);

NAND3xp33_ASAP7_75t_L g15279 ( 
.A(n_15156),
.B(n_6441),
.C(n_6429),
.Y(n_15279)
);

AOI21xp5_ASAP7_75t_L g15280 ( 
.A1(n_15182),
.A2(n_7782),
.B(n_6413),
.Y(n_15280)
);

AND5x1_ASAP7_75t_L g15281 ( 
.A(n_15184),
.B(n_6413),
.C(n_6426),
.D(n_6422),
.E(n_6415),
.Y(n_15281)
);

INVx1_ASAP7_75t_L g15282 ( 
.A(n_15099),
.Y(n_15282)
);

NAND2xp5_ASAP7_75t_L g15283 ( 
.A(n_15100),
.B(n_7418),
.Y(n_15283)
);

NOR2x1_ASAP7_75t_L g15284 ( 
.A(n_15136),
.B(n_6568),
.Y(n_15284)
);

NAND4xp25_ASAP7_75t_L g15285 ( 
.A(n_15142),
.B(n_15135),
.C(n_15153),
.D(n_15137),
.Y(n_15285)
);

NAND4xp75_ASAP7_75t_L g15286 ( 
.A(n_15138),
.B(n_6317),
.C(n_5546),
.D(n_5950),
.Y(n_15286)
);

NOR2xp33_ASAP7_75t_L g15287 ( 
.A(n_15120),
.B(n_7343),
.Y(n_15287)
);

NAND2xp5_ASAP7_75t_L g15288 ( 
.A(n_15076),
.B(n_7465),
.Y(n_15288)
);

NOR2xp67_ASAP7_75t_L g15289 ( 
.A(n_15130),
.B(n_15133),
.Y(n_15289)
);

AND2x2_ASAP7_75t_L g15290 ( 
.A(n_15111),
.B(n_6614),
.Y(n_15290)
);

AND3x1_ASAP7_75t_L g15291 ( 
.A(n_15161),
.B(n_6417),
.C(n_5820),
.Y(n_15291)
);

NAND3xp33_ASAP7_75t_L g15292 ( 
.A(n_15109),
.B(n_6555),
.C(n_6441),
.Y(n_15292)
);

INVx1_ASAP7_75t_L g15293 ( 
.A(n_15185),
.Y(n_15293)
);

NOR4xp75_ASAP7_75t_SL g15294 ( 
.A(n_15128),
.B(n_5914),
.C(n_5926),
.D(n_5916),
.Y(n_15294)
);

OAI21xp33_ASAP7_75t_L g15295 ( 
.A1(n_15144),
.A2(n_6568),
.B(n_7465),
.Y(n_15295)
);

OAI211xp5_ASAP7_75t_L g15296 ( 
.A1(n_15105),
.A2(n_6588),
.B(n_6555),
.C(n_5823),
.Y(n_15296)
);

INVx1_ASAP7_75t_L g15297 ( 
.A(n_15165),
.Y(n_15297)
);

NOR2x1_ASAP7_75t_L g15298 ( 
.A(n_15188),
.B(n_15180),
.Y(n_15298)
);

NAND4xp25_ASAP7_75t_L g15299 ( 
.A(n_15139),
.B(n_6385),
.C(n_6386),
.D(n_6379),
.Y(n_15299)
);

INVx1_ASAP7_75t_L g15300 ( 
.A(n_15094),
.Y(n_15300)
);

AND4x2_ASAP7_75t_L g15301 ( 
.A(n_15079),
.B(n_7570),
.C(n_7663),
.D(n_7343),
.Y(n_15301)
);

INVx4_ASAP7_75t_L g15302 ( 
.A(n_15193),
.Y(n_15302)
);

AOI211xp5_ASAP7_75t_L g15303 ( 
.A1(n_15210),
.A2(n_15155),
.B(n_15189),
.C(n_15159),
.Y(n_15303)
);

NOR3xp33_ASAP7_75t_L g15304 ( 
.A(n_15199),
.B(n_15191),
.C(n_5916),
.Y(n_15304)
);

OAI211xp5_ASAP7_75t_L g15305 ( 
.A1(n_15220),
.A2(n_6588),
.B(n_7773),
.C(n_7766),
.Y(n_15305)
);

AOI321xp33_ASAP7_75t_L g15306 ( 
.A1(n_15227),
.A2(n_6499),
.A3(n_6523),
.B1(n_6465),
.B2(n_6166),
.C(n_6370),
.Y(n_15306)
);

AOI221xp5_ASAP7_75t_L g15307 ( 
.A1(n_15236),
.A2(n_6568),
.B1(n_7776),
.B2(n_7779),
.C(n_7773),
.Y(n_15307)
);

AOI22xp5_ASAP7_75t_L g15308 ( 
.A1(n_15236),
.A2(n_6568),
.B1(n_7663),
.B2(n_7570),
.Y(n_15308)
);

AOI221xp5_ASAP7_75t_L g15309 ( 
.A1(n_15257),
.A2(n_7785),
.B1(n_7790),
.B2(n_7779),
.C(n_7776),
.Y(n_15309)
);

AOI22xp33_ASAP7_75t_L g15310 ( 
.A1(n_15193),
.A2(n_7570),
.B1(n_7728),
.B2(n_7663),
.Y(n_15310)
);

OAI211xp5_ASAP7_75t_L g15311 ( 
.A1(n_15198),
.A2(n_7790),
.B(n_7792),
.C(n_7785),
.Y(n_15311)
);

NAND2xp5_ASAP7_75t_L g15312 ( 
.A(n_15287),
.B(n_7465),
.Y(n_15312)
);

AOI211x1_ASAP7_75t_SL g15313 ( 
.A1(n_15215),
.A2(n_7261),
.B(n_7292),
.C(n_7255),
.Y(n_15313)
);

INVx1_ASAP7_75t_L g15314 ( 
.A(n_15214),
.Y(n_15314)
);

O2A1O1Ixp33_ASAP7_75t_L g15315 ( 
.A1(n_15271),
.A2(n_5820),
.B(n_5842),
.C(n_5791),
.Y(n_15315)
);

CKINVDCx20_ASAP7_75t_R g15316 ( 
.A(n_15204),
.Y(n_15316)
);

AOI22xp5_ASAP7_75t_L g15317 ( 
.A1(n_15231),
.A2(n_7663),
.B1(n_7769),
.B2(n_7728),
.Y(n_15317)
);

XOR2x2_ASAP7_75t_L g15318 ( 
.A(n_15298),
.B(n_5150),
.Y(n_15318)
);

INVxp67_ASAP7_75t_SL g15319 ( 
.A(n_15233),
.Y(n_15319)
);

AOI22xp5_ASAP7_75t_L g15320 ( 
.A1(n_15195),
.A2(n_7769),
.B1(n_7728),
.B2(n_7329),
.Y(n_15320)
);

AOI211xp5_ASAP7_75t_L g15321 ( 
.A1(n_15289),
.A2(n_6317),
.B(n_6119),
.C(n_5853),
.Y(n_15321)
);

AOI221xp5_ASAP7_75t_L g15322 ( 
.A1(n_15194),
.A2(n_7792),
.B1(n_5866),
.B2(n_5880),
.C(n_5853),
.Y(n_15322)
);

OAI21xp5_ASAP7_75t_SL g15323 ( 
.A1(n_15202),
.A2(n_6066),
.B(n_6440),
.Y(n_15323)
);

AOI221xp5_ASAP7_75t_L g15324 ( 
.A1(n_15208),
.A2(n_5866),
.B1(n_5880),
.B2(n_5853),
.C(n_5830),
.Y(n_15324)
);

NAND2xp5_ASAP7_75t_L g15325 ( 
.A(n_15247),
.B(n_6748),
.Y(n_15325)
);

AOI21xp5_ASAP7_75t_L g15326 ( 
.A1(n_15223),
.A2(n_7782),
.B(n_6851),
.Y(n_15326)
);

INVxp33_ASAP7_75t_SL g15327 ( 
.A(n_15196),
.Y(n_15327)
);

BUFx2_ASAP7_75t_L g15328 ( 
.A(n_15213),
.Y(n_15328)
);

AOI22xp5_ASAP7_75t_L g15329 ( 
.A1(n_15278),
.A2(n_7728),
.B1(n_7769),
.B2(n_7329),
.Y(n_15329)
);

NAND2xp5_ASAP7_75t_SL g15330 ( 
.A(n_15193),
.B(n_7329),
.Y(n_15330)
);

OAI221xp5_ASAP7_75t_SL g15331 ( 
.A1(n_15250),
.A2(n_6851),
.B1(n_6119),
.B2(n_6605),
.C(n_7261),
.Y(n_15331)
);

AND4x1_ASAP7_75t_L g15332 ( 
.A(n_15217),
.B(n_6325),
.C(n_5926),
.D(n_5914),
.Y(n_15332)
);

NOR4xp75_ASAP7_75t_L g15333 ( 
.A(n_15221),
.B(n_6325),
.C(n_6376),
.D(n_6505),
.Y(n_15333)
);

AOI211xp5_ASAP7_75t_L g15334 ( 
.A1(n_15293),
.A2(n_5853),
.B(n_5866),
.C(n_5830),
.Y(n_15334)
);

AOI221xp5_ASAP7_75t_L g15335 ( 
.A1(n_15232),
.A2(n_5866),
.B1(n_5880),
.B2(n_5853),
.C(n_5830),
.Y(n_15335)
);

AOI322xp5_ASAP7_75t_L g15336 ( 
.A1(n_15267),
.A2(n_5842),
.A3(n_5869),
.B1(n_5958),
.B2(n_5977),
.C1(n_5937),
.C2(n_5791),
.Y(n_15336)
);

NAND2xp5_ASAP7_75t_L g15337 ( 
.A(n_15290),
.B(n_6748),
.Y(n_15337)
);

AOI222xp33_ASAP7_75t_L g15338 ( 
.A1(n_15218),
.A2(n_5880),
.B1(n_5853),
.B2(n_5993),
.C1(n_5933),
.C2(n_5866),
.Y(n_15338)
);

NAND5xp2_ASAP7_75t_L g15339 ( 
.A(n_15246),
.B(n_5121),
.C(n_5884),
.D(n_5900),
.E(n_5861),
.Y(n_15339)
);

NAND4xp75_ASAP7_75t_L g15340 ( 
.A(n_15282),
.B(n_5546),
.C(n_6361),
.D(n_6357),
.Y(n_15340)
);

BUFx6f_ASAP7_75t_L g15341 ( 
.A(n_15272),
.Y(n_15341)
);

OAI22xp5_ASAP7_75t_L g15342 ( 
.A1(n_15234),
.A2(n_7308),
.B1(n_7318),
.B2(n_7292),
.Y(n_15342)
);

NOR2x1_ASAP7_75t_L g15343 ( 
.A(n_15268),
.B(n_5501),
.Y(n_15343)
);

AOI22xp5_ASAP7_75t_L g15344 ( 
.A1(n_15270),
.A2(n_7329),
.B1(n_6871),
.B2(n_6962),
.Y(n_15344)
);

OAI22x1_ASAP7_75t_L g15345 ( 
.A1(n_15263),
.A2(n_15297),
.B1(n_15300),
.B2(n_15264),
.Y(n_15345)
);

AOI211xp5_ASAP7_75t_L g15346 ( 
.A1(n_15285),
.A2(n_5853),
.B(n_5866),
.C(n_5830),
.Y(n_15346)
);

AND2x2_ASAP7_75t_L g15347 ( 
.A(n_15273),
.B(n_15245),
.Y(n_15347)
);

AOI221xp5_ASAP7_75t_L g15348 ( 
.A1(n_15256),
.A2(n_5830),
.B1(n_5880),
.B2(n_5866),
.C(n_5853),
.Y(n_15348)
);

OAI21xp33_ASAP7_75t_SL g15349 ( 
.A1(n_15259),
.A2(n_6125),
.B(n_5937),
.Y(n_15349)
);

CKINVDCx20_ASAP7_75t_R g15350 ( 
.A(n_15252),
.Y(n_15350)
);

NAND4xp25_ASAP7_75t_L g15351 ( 
.A(n_15201),
.B(n_6605),
.C(n_6577),
.D(n_6523),
.Y(n_15351)
);

AOI221x1_ASAP7_75t_L g15352 ( 
.A1(n_15216),
.A2(n_7318),
.B1(n_7308),
.B2(n_7292),
.C(n_5880),
.Y(n_15352)
);

AOI322xp5_ASAP7_75t_L g15353 ( 
.A1(n_15275),
.A2(n_5869),
.A3(n_5977),
.B1(n_6060),
.B2(n_6085),
.C1(n_6022),
.C2(n_5958),
.Y(n_15353)
);

AOI22xp33_ASAP7_75t_L g15354 ( 
.A1(n_15248),
.A2(n_7329),
.B1(n_5866),
.B2(n_5880),
.Y(n_15354)
);

AOI22xp5_ASAP7_75t_L g15355 ( 
.A1(n_15225),
.A2(n_7329),
.B1(n_6871),
.B2(n_6962),
.Y(n_15355)
);

INVxp67_ASAP7_75t_L g15356 ( 
.A(n_15230),
.Y(n_15356)
);

AOI221xp5_ASAP7_75t_SL g15357 ( 
.A1(n_15288),
.A2(n_5933),
.B1(n_5993),
.B2(n_5880),
.C(n_5830),
.Y(n_15357)
);

INVx1_ASAP7_75t_L g15358 ( 
.A(n_15205),
.Y(n_15358)
);

AOI22xp5_ASAP7_75t_L g15359 ( 
.A1(n_15235),
.A2(n_7329),
.B1(n_6871),
.B2(n_6962),
.Y(n_15359)
);

INVx1_ASAP7_75t_L g15360 ( 
.A(n_15266),
.Y(n_15360)
);

HB1xp67_ASAP7_75t_L g15361 ( 
.A(n_15253),
.Y(n_15361)
);

NOR3xp33_ASAP7_75t_L g15362 ( 
.A(n_15283),
.B(n_5977),
.C(n_5958),
.Y(n_15362)
);

OAI211xp5_ASAP7_75t_L g15363 ( 
.A1(n_15239),
.A2(n_5823),
.B(n_5836),
.C(n_5795),
.Y(n_15363)
);

OAI221xp5_ASAP7_75t_SL g15364 ( 
.A1(n_15219),
.A2(n_6851),
.B1(n_7318),
.B2(n_7308),
.C(n_6264),
.Y(n_15364)
);

NAND4xp25_ASAP7_75t_L g15365 ( 
.A(n_15279),
.B(n_6577),
.C(n_6523),
.D(n_6499),
.Y(n_15365)
);

INVxp67_ASAP7_75t_L g15366 ( 
.A(n_15284),
.Y(n_15366)
);

O2A1O1Ixp33_ASAP7_75t_L g15367 ( 
.A1(n_15277),
.A2(n_6060),
.B(n_6085),
.C(n_6022),
.Y(n_15367)
);

OAI22xp5_ASAP7_75t_L g15368 ( 
.A1(n_15292),
.A2(n_6625),
.B1(n_6615),
.B2(n_5836),
.Y(n_15368)
);

OAI221xp5_ASAP7_75t_L g15369 ( 
.A1(n_15242),
.A2(n_6851),
.B1(n_6085),
.B2(n_6092),
.C(n_6060),
.Y(n_15369)
);

AOI22xp33_ASAP7_75t_L g15370 ( 
.A1(n_15238),
.A2(n_7329),
.B1(n_5830),
.B2(n_5993),
.Y(n_15370)
);

A2O1A1Ixp33_ASAP7_75t_L g15371 ( 
.A1(n_15244),
.A2(n_6625),
.B(n_6615),
.C(n_6092),
.Y(n_15371)
);

INVx1_ASAP7_75t_L g15372 ( 
.A(n_15261),
.Y(n_15372)
);

INVx1_ASAP7_75t_L g15373 ( 
.A(n_15226),
.Y(n_15373)
);

AOI211xp5_ASAP7_75t_SL g15374 ( 
.A1(n_15296),
.A2(n_15251),
.B(n_15200),
.C(n_15274),
.Y(n_15374)
);

NAND2xp5_ASAP7_75t_SL g15375 ( 
.A(n_15294),
.B(n_15291),
.Y(n_15375)
);

AND3x4_ASAP7_75t_L g15376 ( 
.A(n_15258),
.B(n_6166),
.C(n_6100),
.Y(n_15376)
);

AOI222xp33_ASAP7_75t_L g15377 ( 
.A1(n_15229),
.A2(n_5994),
.B1(n_5933),
.B2(n_6007),
.C1(n_5993),
.C2(n_5830),
.Y(n_15377)
);

AOI221x1_ASAP7_75t_L g15378 ( 
.A1(n_15255),
.A2(n_5994),
.B1(n_6007),
.B2(n_5993),
.C(n_5933),
.Y(n_15378)
);

NOR3x1_ASAP7_75t_L g15379 ( 
.A(n_15207),
.B(n_6092),
.C(n_6022),
.Y(n_15379)
);

NOR3xp33_ASAP7_75t_L g15380 ( 
.A(n_15241),
.B(n_6158),
.C(n_6130),
.Y(n_15380)
);

O2A1O1Ixp33_ASAP7_75t_L g15381 ( 
.A1(n_15209),
.A2(n_6158),
.B(n_6171),
.C(n_6130),
.Y(n_15381)
);

OAI211xp5_ASAP7_75t_L g15382 ( 
.A1(n_15254),
.A2(n_5925),
.B(n_5961),
.C(n_5795),
.Y(n_15382)
);

NAND2xp5_ASAP7_75t_L g15383 ( 
.A(n_15228),
.B(n_6748),
.Y(n_15383)
);

OAI22xp5_ASAP7_75t_L g15384 ( 
.A1(n_15240),
.A2(n_5961),
.B1(n_5979),
.B2(n_5925),
.Y(n_15384)
);

XNOR2xp5_ASAP7_75t_L g15385 ( 
.A(n_15222),
.B(n_5816),
.Y(n_15385)
);

AOI211xp5_ASAP7_75t_SL g15386 ( 
.A1(n_15295),
.A2(n_5979),
.B(n_6267),
.C(n_6259),
.Y(n_15386)
);

NAND2x1_ASAP7_75t_L g15387 ( 
.A(n_15211),
.B(n_6004),
.Y(n_15387)
);

NOR3xp33_ASAP7_75t_L g15388 ( 
.A(n_15280),
.B(n_6158),
.C(n_6130),
.Y(n_15388)
);

NAND4xp25_ASAP7_75t_L g15389 ( 
.A(n_15206),
.B(n_6523),
.C(n_6499),
.D(n_6166),
.Y(n_15389)
);

NAND2xp5_ASAP7_75t_L g15390 ( 
.A(n_15224),
.B(n_6748),
.Y(n_15390)
);

AOI22xp5_ASAP7_75t_L g15391 ( 
.A1(n_15203),
.A2(n_7329),
.B1(n_6962),
.B2(n_6871),
.Y(n_15391)
);

AOI211xp5_ASAP7_75t_L g15392 ( 
.A1(n_15243),
.A2(n_5993),
.B(n_5994),
.C(n_5933),
.Y(n_15392)
);

OAI211xp5_ASAP7_75t_SL g15393 ( 
.A1(n_15262),
.A2(n_6139),
.B(n_6422),
.C(n_6415),
.Y(n_15393)
);

NAND4xp25_ASAP7_75t_L g15394 ( 
.A(n_15276),
.B(n_6523),
.C(n_6499),
.D(n_6166),
.Y(n_15394)
);

AOI211xp5_ASAP7_75t_SL g15395 ( 
.A1(n_15197),
.A2(n_15301),
.B(n_15237),
.C(n_15281),
.Y(n_15395)
);

OAI311xp33_ASAP7_75t_L g15396 ( 
.A1(n_15299),
.A2(n_6078),
.A3(n_6376),
.B1(n_6622),
.C1(n_6608),
.Y(n_15396)
);

INVxp67_ASAP7_75t_L g15397 ( 
.A(n_15260),
.Y(n_15397)
);

OR2x2_ASAP7_75t_L g15398 ( 
.A(n_15212),
.B(n_6239),
.Y(n_15398)
);

OAI211xp5_ASAP7_75t_SL g15399 ( 
.A1(n_15265),
.A2(n_15249),
.B(n_15269),
.C(n_15286),
.Y(n_15399)
);

INVx1_ASAP7_75t_L g15400 ( 
.A(n_15214),
.Y(n_15400)
);

NOR2xp33_ASAP7_75t_L g15401 ( 
.A(n_15236),
.B(n_7782),
.Y(n_15401)
);

INVxp67_ASAP7_75t_L g15402 ( 
.A(n_15328),
.Y(n_15402)
);

INVx1_ASAP7_75t_L g15403 ( 
.A(n_15361),
.Y(n_15403)
);

AOI22xp5_ASAP7_75t_L g15404 ( 
.A1(n_15327),
.A2(n_7329),
.B1(n_6195),
.B2(n_6226),
.Y(n_15404)
);

INVxp67_ASAP7_75t_L g15405 ( 
.A(n_15319),
.Y(n_15405)
);

INVx1_ASAP7_75t_L g15406 ( 
.A(n_15302),
.Y(n_15406)
);

INVx2_ASAP7_75t_L g15407 ( 
.A(n_15302),
.Y(n_15407)
);

INVx1_ASAP7_75t_L g15408 ( 
.A(n_15314),
.Y(n_15408)
);

INVx3_ASAP7_75t_L g15409 ( 
.A(n_15400),
.Y(n_15409)
);

INVx2_ASAP7_75t_L g15410 ( 
.A(n_15341),
.Y(n_15410)
);

NAND2xp5_ASAP7_75t_SL g15411 ( 
.A(n_15341),
.B(n_5933),
.Y(n_15411)
);

AOI22xp5_ASAP7_75t_L g15412 ( 
.A1(n_15401),
.A2(n_6195),
.B1(n_6226),
.B2(n_6171),
.Y(n_15412)
);

AOI22xp33_ASAP7_75t_SL g15413 ( 
.A1(n_15341),
.A2(n_5933),
.B1(n_5994),
.B2(n_5993),
.Y(n_15413)
);

INVx1_ASAP7_75t_L g15414 ( 
.A(n_15318),
.Y(n_15414)
);

AOI22xp5_ASAP7_75t_L g15415 ( 
.A1(n_15316),
.A2(n_6195),
.B1(n_6226),
.B2(n_6171),
.Y(n_15415)
);

INVx1_ASAP7_75t_L g15416 ( 
.A(n_15347),
.Y(n_15416)
);

INVx1_ASAP7_75t_L g15417 ( 
.A(n_15360),
.Y(n_15417)
);

NOR2xp33_ASAP7_75t_L g15418 ( 
.A(n_15366),
.B(n_7782),
.Y(n_15418)
);

NOR2x1_ASAP7_75t_L g15419 ( 
.A(n_15372),
.B(n_5501),
.Y(n_15419)
);

AOI22xp5_ASAP7_75t_L g15420 ( 
.A1(n_15350),
.A2(n_6236),
.B1(n_6227),
.B2(n_5993),
.Y(n_15420)
);

INVx1_ASAP7_75t_L g15421 ( 
.A(n_15375),
.Y(n_15421)
);

INVx1_ASAP7_75t_L g15422 ( 
.A(n_15358),
.Y(n_15422)
);

HB1xp67_ASAP7_75t_L g15423 ( 
.A(n_15356),
.Y(n_15423)
);

INVx1_ASAP7_75t_L g15424 ( 
.A(n_15345),
.Y(n_15424)
);

INVx1_ASAP7_75t_L g15425 ( 
.A(n_15373),
.Y(n_15425)
);

INVx1_ASAP7_75t_L g15426 ( 
.A(n_15304),
.Y(n_15426)
);

INVx2_ASAP7_75t_L g15427 ( 
.A(n_15343),
.Y(n_15427)
);

AOI22xp5_ASAP7_75t_L g15428 ( 
.A1(n_15346),
.A2(n_6236),
.B1(n_6227),
.B2(n_5994),
.Y(n_15428)
);

INVx2_ASAP7_75t_L g15429 ( 
.A(n_15337),
.Y(n_15429)
);

INVx1_ASAP7_75t_L g15430 ( 
.A(n_15303),
.Y(n_15430)
);

INVx2_ASAP7_75t_L g15431 ( 
.A(n_15312),
.Y(n_15431)
);

OR2x2_ASAP7_75t_L g15432 ( 
.A(n_15325),
.B(n_6227),
.Y(n_15432)
);

INVx1_ASAP7_75t_L g15433 ( 
.A(n_15399),
.Y(n_15433)
);

NAND2xp5_ASAP7_75t_L g15434 ( 
.A(n_15362),
.B(n_6623),
.Y(n_15434)
);

INVx1_ASAP7_75t_L g15435 ( 
.A(n_15397),
.Y(n_15435)
);

CKINVDCx20_ASAP7_75t_R g15436 ( 
.A(n_15385),
.Y(n_15436)
);

HB1xp67_ASAP7_75t_L g15437 ( 
.A(n_15395),
.Y(n_15437)
);

INVx1_ASAP7_75t_L g15438 ( 
.A(n_15388),
.Y(n_15438)
);

INVx1_ASAP7_75t_L g15439 ( 
.A(n_15383),
.Y(n_15439)
);

INVx1_ASAP7_75t_L g15440 ( 
.A(n_15390),
.Y(n_15440)
);

HB1xp67_ASAP7_75t_L g15441 ( 
.A(n_15349),
.Y(n_15441)
);

INVx2_ASAP7_75t_SL g15442 ( 
.A(n_15376),
.Y(n_15442)
);

BUFx2_ASAP7_75t_L g15443 ( 
.A(n_15398),
.Y(n_15443)
);

INVx1_ASAP7_75t_L g15444 ( 
.A(n_15379),
.Y(n_15444)
);

NOR3xp33_ASAP7_75t_L g15445 ( 
.A(n_15363),
.B(n_15368),
.C(n_15380),
.Y(n_15445)
);

NAND2xp5_ASAP7_75t_SL g15446 ( 
.A(n_15308),
.B(n_5933),
.Y(n_15446)
);

AOI22xp5_ASAP7_75t_L g15447 ( 
.A1(n_15357),
.A2(n_6236),
.B1(n_6007),
.B2(n_6024),
.Y(n_15447)
);

NOR2x2_ASAP7_75t_L g15448 ( 
.A(n_15340),
.B(n_6851),
.Y(n_15448)
);

INVxp67_ASAP7_75t_L g15449 ( 
.A(n_15374),
.Y(n_15449)
);

INVxp67_ASAP7_75t_L g15450 ( 
.A(n_15311),
.Y(n_15450)
);

AOI22xp33_ASAP7_75t_L g15451 ( 
.A1(n_15330),
.A2(n_6007),
.B1(n_6024),
.B2(n_5994),
.Y(n_15451)
);

NOR2xp67_ASAP7_75t_L g15452 ( 
.A(n_15382),
.B(n_6047),
.Y(n_15452)
);

AOI22xp5_ASAP7_75t_L g15453 ( 
.A1(n_15323),
.A2(n_6007),
.B1(n_6024),
.B2(n_5994),
.Y(n_15453)
);

INVx1_ASAP7_75t_L g15454 ( 
.A(n_15305),
.Y(n_15454)
);

NOR2xp67_ASAP7_75t_L g15455 ( 
.A(n_15365),
.B(n_6047),
.Y(n_15455)
);

AND3x2_ASAP7_75t_L g15456 ( 
.A(n_15392),
.B(n_6581),
.C(n_6381),
.Y(n_15456)
);

INVx1_ASAP7_75t_L g15457 ( 
.A(n_15367),
.Y(n_15457)
);

AOI22xp5_ASAP7_75t_L g15458 ( 
.A1(n_15384),
.A2(n_6007),
.B1(n_6024),
.B2(n_5994),
.Y(n_15458)
);

INVx2_ASAP7_75t_L g15459 ( 
.A(n_15387),
.Y(n_15459)
);

NOR3xp33_ASAP7_75t_L g15460 ( 
.A(n_15331),
.B(n_5357),
.C(n_5315),
.Y(n_15460)
);

INVx1_ASAP7_75t_L g15461 ( 
.A(n_15313),
.Y(n_15461)
);

INVx1_ASAP7_75t_L g15462 ( 
.A(n_15371),
.Y(n_15462)
);

INVx1_ASAP7_75t_L g15463 ( 
.A(n_15315),
.Y(n_15463)
);

INVx2_ASAP7_75t_L g15464 ( 
.A(n_15369),
.Y(n_15464)
);

AOI22xp5_ASAP7_75t_L g15465 ( 
.A1(n_15307),
.A2(n_6024),
.B1(n_6062),
.B2(n_6007),
.Y(n_15465)
);

INVx1_ASAP7_75t_L g15466 ( 
.A(n_15378),
.Y(n_15466)
);

NOR2x1_ASAP7_75t_L g15467 ( 
.A(n_15389),
.B(n_5501),
.Y(n_15467)
);

NOR2xp67_ASAP7_75t_L g15468 ( 
.A(n_15326),
.B(n_6047),
.Y(n_15468)
);

AOI22xp5_ASAP7_75t_L g15469 ( 
.A1(n_15351),
.A2(n_6024),
.B1(n_6062),
.B2(n_6007),
.Y(n_15469)
);

NAND2xp5_ASAP7_75t_L g15470 ( 
.A(n_15386),
.B(n_6623),
.Y(n_15470)
);

INVx1_ASAP7_75t_L g15471 ( 
.A(n_15333),
.Y(n_15471)
);

AOI22xp5_ASAP7_75t_L g15472 ( 
.A1(n_15329),
.A2(n_6062),
.B1(n_6155),
.B2(n_6024),
.Y(n_15472)
);

INVx1_ASAP7_75t_L g15473 ( 
.A(n_15394),
.Y(n_15473)
);

NAND2xp5_ASAP7_75t_SL g15474 ( 
.A(n_15336),
.B(n_6024),
.Y(n_15474)
);

AOI22xp5_ASAP7_75t_L g15475 ( 
.A1(n_15310),
.A2(n_6155),
.B1(n_6203),
.B2(n_6062),
.Y(n_15475)
);

INVx1_ASAP7_75t_L g15476 ( 
.A(n_15352),
.Y(n_15476)
);

BUFx3_ASAP7_75t_L g15477 ( 
.A(n_15359),
.Y(n_15477)
);

NOR2x1_ASAP7_75t_L g15478 ( 
.A(n_15381),
.B(n_5582),
.Y(n_15478)
);

INVx1_ASAP7_75t_L g15479 ( 
.A(n_15334),
.Y(n_15479)
);

AOI22xp5_ASAP7_75t_L g15480 ( 
.A1(n_15354),
.A2(n_6155),
.B1(n_6203),
.B2(n_6062),
.Y(n_15480)
);

INVx1_ASAP7_75t_L g15481 ( 
.A(n_15364),
.Y(n_15481)
);

INVx1_ASAP7_75t_L g15482 ( 
.A(n_15321),
.Y(n_15482)
);

INVx1_ASAP7_75t_L g15483 ( 
.A(n_15306),
.Y(n_15483)
);

INVx1_ASAP7_75t_L g15484 ( 
.A(n_15416),
.Y(n_15484)
);

INVx1_ASAP7_75t_L g15485 ( 
.A(n_15418),
.Y(n_15485)
);

NAND2xp5_ASAP7_75t_L g15486 ( 
.A(n_15409),
.B(n_15353),
.Y(n_15486)
);

OA211x2_ASAP7_75t_L g15487 ( 
.A1(n_15405),
.A2(n_15322),
.B(n_15370),
.C(n_15348),
.Y(n_15487)
);

NOR2x1_ASAP7_75t_L g15488 ( 
.A(n_15409),
.B(n_15410),
.Y(n_15488)
);

AND2x4_ASAP7_75t_L g15489 ( 
.A(n_15403),
.B(n_15344),
.Y(n_15489)
);

NOR3xp33_ASAP7_75t_L g15490 ( 
.A(n_15402),
.B(n_15424),
.C(n_15408),
.Y(n_15490)
);

NAND4xp75_ASAP7_75t_L g15491 ( 
.A(n_15421),
.B(n_15320),
.C(n_15317),
.D(n_15391),
.Y(n_15491)
);

NOR4xp25_ASAP7_75t_L g15492 ( 
.A(n_15433),
.B(n_15396),
.C(n_15393),
.D(n_15342),
.Y(n_15492)
);

INVx1_ASAP7_75t_L g15493 ( 
.A(n_15423),
.Y(n_15493)
);

INVx1_ASAP7_75t_L g15494 ( 
.A(n_15441),
.Y(n_15494)
);

NAND2xp5_ASAP7_75t_L g15495 ( 
.A(n_15417),
.B(n_15452),
.Y(n_15495)
);

NOR2x1_ASAP7_75t_L g15496 ( 
.A(n_15406),
.B(n_15339),
.Y(n_15496)
);

OR2x2_ASAP7_75t_L g15497 ( 
.A(n_15470),
.B(n_15355),
.Y(n_15497)
);

AND2x4_ASAP7_75t_L g15498 ( 
.A(n_15422),
.B(n_15332),
.Y(n_15498)
);

NOR3xp33_ASAP7_75t_L g15499 ( 
.A(n_15449),
.B(n_15324),
.C(n_15309),
.Y(n_15499)
);

INVx1_ASAP7_75t_SL g15500 ( 
.A(n_15436),
.Y(n_15500)
);

NAND3xp33_ASAP7_75t_L g15501 ( 
.A(n_15437),
.B(n_15377),
.C(n_15335),
.Y(n_15501)
);

NOR2xp33_ASAP7_75t_L g15502 ( 
.A(n_15407),
.B(n_15338),
.Y(n_15502)
);

HB1xp67_ASAP7_75t_L g15503 ( 
.A(n_15476),
.Y(n_15503)
);

AND3x4_ASAP7_75t_L g15504 ( 
.A(n_15429),
.B(n_5821),
.C(n_5816),
.Y(n_15504)
);

NOR2x1_ASAP7_75t_L g15505 ( 
.A(n_15443),
.B(n_5582),
.Y(n_15505)
);

NOR2x1_ASAP7_75t_L g15506 ( 
.A(n_15425),
.B(n_15427),
.Y(n_15506)
);

AO221x1_ASAP7_75t_L g15507 ( 
.A1(n_15450),
.A2(n_6203),
.B1(n_6271),
.B2(n_6155),
.C(n_6062),
.Y(n_15507)
);

NOR2x1_ASAP7_75t_L g15508 ( 
.A(n_15435),
.B(n_5582),
.Y(n_15508)
);

NAND3x1_ASAP7_75t_L g15509 ( 
.A(n_15439),
.B(n_6241),
.C(n_6259),
.Y(n_15509)
);

AND2x2_ASAP7_75t_L g15510 ( 
.A(n_15483),
.B(n_6623),
.Y(n_15510)
);

AOI22xp5_ASAP7_75t_L g15511 ( 
.A1(n_15430),
.A2(n_15442),
.B1(n_15473),
.B2(n_15440),
.Y(n_15511)
);

BUFx2_ASAP7_75t_SL g15512 ( 
.A(n_15431),
.Y(n_15512)
);

AND3x4_ASAP7_75t_L g15513 ( 
.A(n_15477),
.B(n_5821),
.C(n_5816),
.Y(n_15513)
);

INVx2_ASAP7_75t_L g15514 ( 
.A(n_15419),
.Y(n_15514)
);

NAND2xp33_ASAP7_75t_L g15515 ( 
.A(n_15444),
.B(n_5411),
.Y(n_15515)
);

O2A1O1Ixp33_ASAP7_75t_L g15516 ( 
.A1(n_15414),
.A2(n_6286),
.B(n_6315),
.C(n_6277),
.Y(n_15516)
);

OR2x2_ASAP7_75t_L g15517 ( 
.A(n_15432),
.B(n_6239),
.Y(n_15517)
);

NOR2x1_ASAP7_75t_L g15518 ( 
.A(n_15426),
.B(n_5411),
.Y(n_15518)
);

INVxp67_ASAP7_75t_SL g15519 ( 
.A(n_15466),
.Y(n_15519)
);

NOR2xp67_ASAP7_75t_SL g15520 ( 
.A(n_15481),
.B(n_5411),
.Y(n_15520)
);

AOI22xp33_ASAP7_75t_L g15521 ( 
.A1(n_15445),
.A2(n_6155),
.B1(n_6203),
.B2(n_6062),
.Y(n_15521)
);

AOI211xp5_ASAP7_75t_L g15522 ( 
.A1(n_15454),
.A2(n_5417),
.B(n_5451),
.C(n_5420),
.Y(n_15522)
);

NOR2x1_ASAP7_75t_L g15523 ( 
.A(n_15459),
.B(n_5417),
.Y(n_15523)
);

NAND2xp5_ASAP7_75t_L g15524 ( 
.A(n_15455),
.B(n_6623),
.Y(n_15524)
);

AOI21xp5_ASAP7_75t_L g15525 ( 
.A1(n_15457),
.A2(n_7782),
.B(n_6851),
.Y(n_15525)
);

INVx1_ASAP7_75t_L g15526 ( 
.A(n_15411),
.Y(n_15526)
);

NAND2x1p5_ASAP7_75t_L g15527 ( 
.A(n_15464),
.B(n_5417),
.Y(n_15527)
);

XNOR2xp5_ASAP7_75t_L g15528 ( 
.A(n_15471),
.B(n_6066),
.Y(n_15528)
);

OAI222xp33_ASAP7_75t_L g15529 ( 
.A1(n_15461),
.A2(n_6257),
.B1(n_6258),
.B2(n_6047),
.C1(n_6286),
.C2(n_6277),
.Y(n_15529)
);

HB1xp67_ASAP7_75t_L g15530 ( 
.A(n_15463),
.Y(n_15530)
);

NAND3x1_ASAP7_75t_SL g15531 ( 
.A(n_15478),
.B(n_6656),
.C(n_6361),
.Y(n_15531)
);

CKINVDCx5p33_ASAP7_75t_R g15532 ( 
.A(n_15438),
.Y(n_15532)
);

NOR2x1_ASAP7_75t_L g15533 ( 
.A(n_15479),
.B(n_5417),
.Y(n_15533)
);

NAND4xp75_ASAP7_75t_L g15534 ( 
.A(n_15482),
.B(n_6361),
.C(n_6357),
.D(n_6336),
.Y(n_15534)
);

NAND4xp25_ASAP7_75t_L g15535 ( 
.A(n_15462),
.B(n_5266),
.C(n_5286),
.D(n_5243),
.Y(n_15535)
);

INVx2_ASAP7_75t_L g15536 ( 
.A(n_15448),
.Y(n_15536)
);

OAI22xp5_ASAP7_75t_L g15537 ( 
.A1(n_15468),
.A2(n_6062),
.B1(n_6203),
.B2(n_6155),
.Y(n_15537)
);

AOI22xp5_ASAP7_75t_L g15538 ( 
.A1(n_15460),
.A2(n_6203),
.B1(n_6271),
.B2(n_6155),
.Y(n_15538)
);

NOR3xp33_ASAP7_75t_L g15539 ( 
.A(n_15467),
.B(n_5357),
.C(n_5315),
.Y(n_15539)
);

INVx1_ASAP7_75t_L g15540 ( 
.A(n_15456),
.Y(n_15540)
);

XNOR2x1_ASAP7_75t_L g15541 ( 
.A(n_15434),
.B(n_5417),
.Y(n_15541)
);

NAND2xp5_ASAP7_75t_L g15542 ( 
.A(n_15474),
.B(n_15446),
.Y(n_15542)
);

NAND4xp25_ASAP7_75t_L g15543 ( 
.A(n_15415),
.B(n_5266),
.C(n_5286),
.D(n_5243),
.Y(n_15543)
);

NOR3xp33_ASAP7_75t_L g15544 ( 
.A(n_15420),
.B(n_5357),
.C(n_5315),
.Y(n_15544)
);

OR2x2_ASAP7_75t_L g15545 ( 
.A(n_15412),
.B(n_6239),
.Y(n_15545)
);

AND2x2_ASAP7_75t_SL g15546 ( 
.A(n_15469),
.B(n_5457),
.Y(n_15546)
);

AND2x2_ASAP7_75t_L g15547 ( 
.A(n_15404),
.B(n_6623),
.Y(n_15547)
);

INVx1_ASAP7_75t_L g15548 ( 
.A(n_15413),
.Y(n_15548)
);

O2A1O1Ixp33_ASAP7_75t_L g15549 ( 
.A1(n_15451),
.A2(n_6286),
.B(n_6315),
.C(n_6277),
.Y(n_15549)
);

INVx1_ASAP7_75t_L g15550 ( 
.A(n_15447),
.Y(n_15550)
);

BUFx6f_ASAP7_75t_L g15551 ( 
.A(n_15453),
.Y(n_15551)
);

NOR2xp67_ASAP7_75t_L g15552 ( 
.A(n_15428),
.B(n_6047),
.Y(n_15552)
);

INVx5_ASAP7_75t_L g15553 ( 
.A(n_15475),
.Y(n_15553)
);

NAND4xp75_ASAP7_75t_L g15554 ( 
.A(n_15488),
.B(n_15465),
.C(n_15472),
.D(n_15480),
.Y(n_15554)
);

NOR2x1_ASAP7_75t_L g15555 ( 
.A(n_15506),
.B(n_15458),
.Y(n_15555)
);

AOI21xp5_ASAP7_75t_L g15556 ( 
.A1(n_15519),
.A2(n_7782),
.B(n_6139),
.Y(n_15556)
);

AND2x2_ASAP7_75t_L g15557 ( 
.A(n_15510),
.B(n_6633),
.Y(n_15557)
);

INVx1_ASAP7_75t_L g15558 ( 
.A(n_15503),
.Y(n_15558)
);

NOR2x1_ASAP7_75t_L g15559 ( 
.A(n_15493),
.B(n_5420),
.Y(n_15559)
);

HB1xp67_ASAP7_75t_L g15560 ( 
.A(n_15484),
.Y(n_15560)
);

NAND2xp5_ASAP7_75t_L g15561 ( 
.A(n_15490),
.B(n_6672),
.Y(n_15561)
);

AOI222xp33_ASAP7_75t_L g15562 ( 
.A1(n_15515),
.A2(n_6271),
.B1(n_6155),
.B2(n_6282),
.C1(n_6280),
.C2(n_6203),
.Y(n_15562)
);

AOI221x1_ASAP7_75t_L g15563 ( 
.A1(n_15494),
.A2(n_6203),
.B1(n_6282),
.B2(n_6280),
.C(n_6271),
.Y(n_15563)
);

AND2x2_ASAP7_75t_L g15564 ( 
.A(n_15512),
.B(n_6633),
.Y(n_15564)
);

A2O1A1Ixp33_ASAP7_75t_L g15565 ( 
.A1(n_15502),
.A2(n_6125),
.B(n_6066),
.C(n_6315),
.Y(n_15565)
);

AOI322xp5_ASAP7_75t_L g15566 ( 
.A1(n_15500),
.A2(n_6434),
.A3(n_6355),
.B1(n_6460),
.B2(n_6466),
.C1(n_6392),
.C2(n_6339),
.Y(n_15566)
);

BUFx6f_ASAP7_75t_L g15567 ( 
.A(n_15495),
.Y(n_15567)
);

NAND4xp75_ASAP7_75t_L g15568 ( 
.A(n_15511),
.B(n_6357),
.C(n_6336),
.D(n_6340),
.Y(n_15568)
);

AOI32xp33_ASAP7_75t_L g15569 ( 
.A1(n_15496),
.A2(n_6066),
.A3(n_6211),
.B1(n_6264),
.B2(n_6177),
.Y(n_15569)
);

A2O1A1Ixp33_ASAP7_75t_L g15570 ( 
.A1(n_15540),
.A2(n_6355),
.B(n_6392),
.C(n_6339),
.Y(n_15570)
);

AO22x2_ASAP7_75t_L g15571 ( 
.A1(n_15536),
.A2(n_5514),
.B1(n_5540),
.B2(n_5455),
.Y(n_15571)
);

AOI21xp5_ASAP7_75t_L g15572 ( 
.A1(n_15486),
.A2(n_6426),
.B(n_6078),
.Y(n_15572)
);

INVx1_ASAP7_75t_L g15573 ( 
.A(n_15527),
.Y(n_15573)
);

NOR3xp33_ASAP7_75t_SL g15574 ( 
.A(n_15532),
.B(n_6267),
.C(n_6410),
.Y(n_15574)
);

AOI21xp33_ASAP7_75t_SL g15575 ( 
.A1(n_15501),
.A2(n_5121),
.B(n_5861),
.Y(n_15575)
);

NAND4xp75_ASAP7_75t_L g15576 ( 
.A(n_15487),
.B(n_6336),
.C(n_6340),
.D(n_6329),
.Y(n_15576)
);

OAI22xp5_ASAP7_75t_L g15577 ( 
.A1(n_15528),
.A2(n_6280),
.B1(n_6282),
.B2(n_6271),
.Y(n_15577)
);

OR2x2_ASAP7_75t_L g15578 ( 
.A(n_15524),
.B(n_6271),
.Y(n_15578)
);

NOR2x1p5_ASAP7_75t_L g15579 ( 
.A(n_15491),
.B(n_5420),
.Y(n_15579)
);

NOR4xp75_ASAP7_75t_L g15580 ( 
.A(n_15542),
.B(n_6241),
.C(n_6179),
.D(n_6184),
.Y(n_15580)
);

AND2x4_ASAP7_75t_L g15581 ( 
.A(n_15489),
.B(n_6639),
.Y(n_15581)
);

AOI322xp5_ASAP7_75t_L g15582 ( 
.A1(n_15530),
.A2(n_6434),
.A3(n_6355),
.B1(n_6460),
.B2(n_6466),
.C1(n_6392),
.C2(n_6339),
.Y(n_15582)
);

NOR2x1_ASAP7_75t_L g15583 ( 
.A(n_15526),
.B(n_5420),
.Y(n_15583)
);

OR2x2_ASAP7_75t_L g15584 ( 
.A(n_15492),
.B(n_6271),
.Y(n_15584)
);

AOI22x1_ASAP7_75t_L g15585 ( 
.A1(n_15514),
.A2(n_5420),
.B1(n_5457),
.B2(n_5451),
.Y(n_15585)
);

NOR2x1p5_ASAP7_75t_L g15586 ( 
.A(n_15497),
.B(n_15485),
.Y(n_15586)
);

AND2x4_ASAP7_75t_L g15587 ( 
.A(n_15498),
.B(n_6633),
.Y(n_15587)
);

NOR2x1_ASAP7_75t_L g15588 ( 
.A(n_15548),
.B(n_5420),
.Y(n_15588)
);

INVx1_ASAP7_75t_L g15589 ( 
.A(n_15520),
.Y(n_15589)
);

NOR3xp33_ASAP7_75t_L g15590 ( 
.A(n_15499),
.B(n_5357),
.C(n_5315),
.Y(n_15590)
);

NAND3xp33_ASAP7_75t_L g15591 ( 
.A(n_15553),
.B(n_5370),
.C(n_5321),
.Y(n_15591)
);

OAI211xp5_ASAP7_75t_SL g15592 ( 
.A1(n_15550),
.A2(n_6485),
.B(n_6211),
.C(n_6337),
.Y(n_15592)
);

INVx1_ASAP7_75t_SL g15593 ( 
.A(n_15553),
.Y(n_15593)
);

NAND2xp33_ASAP7_75t_SL g15594 ( 
.A(n_15551),
.B(n_5420),
.Y(n_15594)
);

NOR3xp33_ASAP7_75t_SL g15595 ( 
.A(n_15543),
.B(n_6410),
.C(n_6444),
.Y(n_15595)
);

INVx1_ASAP7_75t_L g15596 ( 
.A(n_15533),
.Y(n_15596)
);

OAI321xp33_ASAP7_75t_L g15597 ( 
.A1(n_15551),
.A2(n_6282),
.A3(n_6271),
.B1(n_6311),
.B2(n_6303),
.C(n_6280),
.Y(n_15597)
);

AND3x1_ASAP7_75t_L g15598 ( 
.A(n_15539),
.B(n_6460),
.C(n_6434),
.Y(n_15598)
);

AND2x4_ASAP7_75t_L g15599 ( 
.A(n_15523),
.B(n_6633),
.Y(n_15599)
);

AND2x4_ASAP7_75t_L g15600 ( 
.A(n_15547),
.B(n_6633),
.Y(n_15600)
);

NAND4xp75_ASAP7_75t_L g15601 ( 
.A(n_15518),
.B(n_15505),
.C(n_15552),
.D(n_15508),
.Y(n_15601)
);

OAI211xp5_ASAP7_75t_L g15602 ( 
.A1(n_15553),
.A2(n_5451),
.B(n_5457),
.C(n_5420),
.Y(n_15602)
);

AND2x2_ASAP7_75t_L g15603 ( 
.A(n_15541),
.B(n_6639),
.Y(n_15603)
);

NOR2x1_ASAP7_75t_L g15604 ( 
.A(n_15513),
.B(n_5451),
.Y(n_15604)
);

OR3x2_ASAP7_75t_L g15605 ( 
.A(n_15531),
.B(n_15535),
.C(n_15517),
.Y(n_15605)
);

NAND2xp5_ASAP7_75t_SL g15606 ( 
.A(n_15546),
.B(n_15522),
.Y(n_15606)
);

XNOR2x1_ASAP7_75t_L g15607 ( 
.A(n_15504),
.B(n_5451),
.Y(n_15607)
);

AOI221xp5_ASAP7_75t_L g15608 ( 
.A1(n_15525),
.A2(n_6282),
.B1(n_6311),
.B2(n_6303),
.C(n_6280),
.Y(n_15608)
);

INVx1_ASAP7_75t_L g15609 ( 
.A(n_15584),
.Y(n_15609)
);

NAND4xp75_ASAP7_75t_L g15610 ( 
.A(n_15555),
.B(n_15538),
.C(n_15507),
.D(n_15544),
.Y(n_15610)
);

NAND2xp5_ASAP7_75t_L g15611 ( 
.A(n_15593),
.B(n_15549),
.Y(n_15611)
);

NAND2xp5_ASAP7_75t_L g15612 ( 
.A(n_15558),
.B(n_15545),
.Y(n_15612)
);

INVx2_ASAP7_75t_L g15613 ( 
.A(n_15579),
.Y(n_15613)
);

INVx1_ASAP7_75t_L g15614 ( 
.A(n_15560),
.Y(n_15614)
);

OAI211xp5_ASAP7_75t_SL g15615 ( 
.A1(n_15589),
.A2(n_15516),
.B(n_15521),
.C(n_15537),
.Y(n_15615)
);

INVx4_ASAP7_75t_L g15616 ( 
.A(n_15567),
.Y(n_15616)
);

INVx2_ASAP7_75t_SL g15617 ( 
.A(n_15586),
.Y(n_15617)
);

HB1xp67_ASAP7_75t_L g15618 ( 
.A(n_15573),
.Y(n_15618)
);

XOR2xp5_ASAP7_75t_L g15619 ( 
.A(n_15605),
.B(n_15534),
.Y(n_15619)
);

INVx1_ASAP7_75t_L g15620 ( 
.A(n_15561),
.Y(n_15620)
);

XNOR2xp5_ASAP7_75t_L g15621 ( 
.A(n_15554),
.B(n_15509),
.Y(n_15621)
);

NAND2x1p5_ASAP7_75t_L g15622 ( 
.A(n_15567),
.B(n_15529),
.Y(n_15622)
);

INVx2_ASAP7_75t_L g15623 ( 
.A(n_15559),
.Y(n_15623)
);

AO22x1_ASAP7_75t_L g15624 ( 
.A1(n_15596),
.A2(n_5370),
.B1(n_5653),
.B2(n_5321),
.Y(n_15624)
);

XNOR2xp5_ASAP7_75t_L g15625 ( 
.A(n_15564),
.B(n_5121),
.Y(n_15625)
);

XNOR2x1_ASAP7_75t_L g15626 ( 
.A(n_15601),
.B(n_5516),
.Y(n_15626)
);

CKINVDCx5p33_ASAP7_75t_R g15627 ( 
.A(n_15606),
.Y(n_15627)
);

AND2x2_ASAP7_75t_L g15628 ( 
.A(n_15581),
.B(n_6639),
.Y(n_15628)
);

INVx2_ASAP7_75t_L g15629 ( 
.A(n_15583),
.Y(n_15629)
);

INVx2_ASAP7_75t_L g15630 ( 
.A(n_15588),
.Y(n_15630)
);

INVx3_ASAP7_75t_L g15631 ( 
.A(n_15587),
.Y(n_15631)
);

INVx1_ASAP7_75t_L g15632 ( 
.A(n_15594),
.Y(n_15632)
);

NAND2xp5_ASAP7_75t_L g15633 ( 
.A(n_15607),
.B(n_6639),
.Y(n_15633)
);

BUFx6f_ASAP7_75t_L g15634 ( 
.A(n_15578),
.Y(n_15634)
);

NOR2x1_ASAP7_75t_L g15635 ( 
.A(n_15604),
.B(n_5451),
.Y(n_15635)
);

INVx6_ASAP7_75t_L g15636 ( 
.A(n_15603),
.Y(n_15636)
);

HB1xp67_ASAP7_75t_L g15637 ( 
.A(n_15598),
.Y(n_15637)
);

INVx1_ASAP7_75t_L g15638 ( 
.A(n_15591),
.Y(n_15638)
);

AOI22xp5_ASAP7_75t_L g15639 ( 
.A1(n_15576),
.A2(n_15590),
.B1(n_15600),
.B2(n_15599),
.Y(n_15639)
);

INVxp33_ASAP7_75t_SL g15640 ( 
.A(n_15557),
.Y(n_15640)
);

AOI21xp5_ASAP7_75t_L g15641 ( 
.A1(n_15572),
.A2(n_6499),
.B(n_6381),
.Y(n_15641)
);

AND2x4_ASAP7_75t_L g15642 ( 
.A(n_15595),
.B(n_15563),
.Y(n_15642)
);

NOR3xp33_ASAP7_75t_L g15643 ( 
.A(n_15592),
.B(n_5357),
.C(n_5315),
.Y(n_15643)
);

CKINVDCx20_ASAP7_75t_R g15644 ( 
.A(n_15574),
.Y(n_15644)
);

OAI22xp5_ASAP7_75t_SL g15645 ( 
.A1(n_15577),
.A2(n_5451),
.B1(n_5458),
.B2(n_5457),
.Y(n_15645)
);

INVx1_ASAP7_75t_L g15646 ( 
.A(n_15571),
.Y(n_15646)
);

INVx1_ASAP7_75t_L g15647 ( 
.A(n_15571),
.Y(n_15647)
);

HB1xp67_ASAP7_75t_L g15648 ( 
.A(n_15580),
.Y(n_15648)
);

XOR2xp5_ASAP7_75t_L g15649 ( 
.A(n_15568),
.B(n_5451),
.Y(n_15649)
);

XNOR2xp5_ASAP7_75t_L g15650 ( 
.A(n_15556),
.B(n_5121),
.Y(n_15650)
);

INVx2_ASAP7_75t_L g15651 ( 
.A(n_15585),
.Y(n_15651)
);

INVx1_ASAP7_75t_L g15652 ( 
.A(n_15602),
.Y(n_15652)
);

NAND2xp33_ASAP7_75t_L g15653 ( 
.A(n_15569),
.B(n_5451),
.Y(n_15653)
);

AND3x4_ASAP7_75t_L g15654 ( 
.A(n_15575),
.B(n_5821),
.C(n_5816),
.Y(n_15654)
);

NAND2xp5_ASAP7_75t_L g15655 ( 
.A(n_15570),
.B(n_6639),
.Y(n_15655)
);

NAND2x1p5_ASAP7_75t_L g15656 ( 
.A(n_15597),
.B(n_5451),
.Y(n_15656)
);

NAND3xp33_ASAP7_75t_SL g15657 ( 
.A(n_15565),
.B(n_5884),
.C(n_5861),
.Y(n_15657)
);

NAND2xp5_ASAP7_75t_SL g15658 ( 
.A(n_15608),
.B(n_6280),
.Y(n_15658)
);

AOI22x1_ASAP7_75t_L g15659 ( 
.A1(n_15619),
.A2(n_15562),
.B1(n_15566),
.B2(n_15582),
.Y(n_15659)
);

NOR3xp33_ASAP7_75t_SL g15660 ( 
.A(n_15627),
.B(n_6443),
.C(n_6444),
.Y(n_15660)
);

OAI21xp5_ASAP7_75t_L g15661 ( 
.A1(n_15614),
.A2(n_15618),
.B(n_15617),
.Y(n_15661)
);

AO21x2_ASAP7_75t_L g15662 ( 
.A1(n_15609),
.A2(n_6239),
.B(n_6179),
.Y(n_15662)
);

INVx1_ASAP7_75t_L g15663 ( 
.A(n_15621),
.Y(n_15663)
);

XNOR2x1_ASAP7_75t_L g15664 ( 
.A(n_15622),
.B(n_5457),
.Y(n_15664)
);

OAI22x1_ASAP7_75t_L g15665 ( 
.A1(n_15616),
.A2(n_6257),
.B1(n_6258),
.B2(n_6047),
.Y(n_15665)
);

AOI22xp5_ASAP7_75t_L g15666 ( 
.A1(n_15640),
.A2(n_6311),
.B1(n_6328),
.B2(n_6282),
.Y(n_15666)
);

OAI22xp5_ASAP7_75t_L g15667 ( 
.A1(n_15626),
.A2(n_6282),
.B1(n_6303),
.B2(n_6280),
.Y(n_15667)
);

OAI22xp5_ASAP7_75t_L g15668 ( 
.A1(n_15639),
.A2(n_6282),
.B1(n_6303),
.B2(n_6280),
.Y(n_15668)
);

INVx2_ASAP7_75t_L g15669 ( 
.A(n_15631),
.Y(n_15669)
);

AOI22xp5_ASAP7_75t_L g15670 ( 
.A1(n_15636),
.A2(n_6303),
.B1(n_6328),
.B2(n_6311),
.Y(n_15670)
);

CKINVDCx20_ASAP7_75t_R g15671 ( 
.A(n_15644),
.Y(n_15671)
);

INVx2_ASAP7_75t_L g15672 ( 
.A(n_15634),
.Y(n_15672)
);

INVx2_ASAP7_75t_L g15673 ( 
.A(n_15634),
.Y(n_15673)
);

HB1xp67_ASAP7_75t_L g15674 ( 
.A(n_15637),
.Y(n_15674)
);

INVx1_ASAP7_75t_L g15675 ( 
.A(n_15613),
.Y(n_15675)
);

INVx1_ASAP7_75t_L g15676 ( 
.A(n_15648),
.Y(n_15676)
);

INVx2_ASAP7_75t_L g15677 ( 
.A(n_15636),
.Y(n_15677)
);

NAND2xp5_ASAP7_75t_L g15678 ( 
.A(n_15642),
.B(n_5816),
.Y(n_15678)
);

NAND3xp33_ASAP7_75t_L g15679 ( 
.A(n_15611),
.B(n_5370),
.C(n_5321),
.Y(n_15679)
);

AOI22xp5_ASAP7_75t_L g15680 ( 
.A1(n_15620),
.A2(n_6303),
.B1(n_6328),
.B2(n_6311),
.Y(n_15680)
);

NAND3xp33_ASAP7_75t_L g15681 ( 
.A(n_15612),
.B(n_5370),
.C(n_5321),
.Y(n_15681)
);

OA22x2_ASAP7_75t_L g15682 ( 
.A1(n_15638),
.A2(n_6479),
.B1(n_6512),
.B2(n_6466),
.Y(n_15682)
);

AO21x2_ASAP7_75t_L g15683 ( 
.A1(n_15630),
.A2(n_6239),
.B(n_6184),
.Y(n_15683)
);

OAI22x1_ASAP7_75t_L g15684 ( 
.A1(n_15652),
.A2(n_6257),
.B1(n_6258),
.B2(n_6047),
.Y(n_15684)
);

AOI22x1_ASAP7_75t_L g15685 ( 
.A1(n_15623),
.A2(n_5457),
.B1(n_5475),
.B2(n_5459),
.Y(n_15685)
);

INVx1_ASAP7_75t_L g15686 ( 
.A(n_15646),
.Y(n_15686)
);

XNOR2x1_ASAP7_75t_L g15687 ( 
.A(n_15610),
.B(n_5457),
.Y(n_15687)
);

INVx2_ASAP7_75t_L g15688 ( 
.A(n_15651),
.Y(n_15688)
);

INVx1_ASAP7_75t_L g15689 ( 
.A(n_15647),
.Y(n_15689)
);

INVx1_ASAP7_75t_L g15690 ( 
.A(n_15629),
.Y(n_15690)
);

AOI21xp5_ASAP7_75t_L g15691 ( 
.A1(n_15632),
.A2(n_6364),
.B(n_6455),
.Y(n_15691)
);

BUFx2_ASAP7_75t_L g15692 ( 
.A(n_15635),
.Y(n_15692)
);

INVx1_ASAP7_75t_L g15693 ( 
.A(n_15615),
.Y(n_15693)
);

OAI22xp5_ASAP7_75t_SL g15694 ( 
.A1(n_15649),
.A2(n_5457),
.B1(n_5459),
.B2(n_5458),
.Y(n_15694)
);

INVx1_ASAP7_75t_L g15695 ( 
.A(n_15653),
.Y(n_15695)
);

XOR2x2_ASAP7_75t_L g15696 ( 
.A(n_15633),
.B(n_5121),
.Y(n_15696)
);

OAI22xp5_ASAP7_75t_L g15697 ( 
.A1(n_15669),
.A2(n_15687),
.B1(n_15677),
.B2(n_15671),
.Y(n_15697)
);

OAI22xp5_ASAP7_75t_L g15698 ( 
.A1(n_15690),
.A2(n_15656),
.B1(n_15650),
.B2(n_15654),
.Y(n_15698)
);

AO22x1_ASAP7_75t_L g15699 ( 
.A1(n_15661),
.A2(n_15643),
.B1(n_15628),
.B2(n_15655),
.Y(n_15699)
);

AOI22xp5_ASAP7_75t_L g15700 ( 
.A1(n_15676),
.A2(n_15693),
.B1(n_15674),
.B2(n_15663),
.Y(n_15700)
);

INVx2_ASAP7_75t_L g15701 ( 
.A(n_15664),
.Y(n_15701)
);

INVx1_ASAP7_75t_L g15702 ( 
.A(n_15686),
.Y(n_15702)
);

INVx1_ASAP7_75t_L g15703 ( 
.A(n_15689),
.Y(n_15703)
);

OAI22x1_ASAP7_75t_L g15704 ( 
.A1(n_15672),
.A2(n_15625),
.B1(n_15658),
.B2(n_15657),
.Y(n_15704)
);

AOI22xp33_ASAP7_75t_SL g15705 ( 
.A1(n_15659),
.A2(n_15645),
.B1(n_15641),
.B2(n_15624),
.Y(n_15705)
);

OAI22xp5_ASAP7_75t_SL g15706 ( 
.A1(n_15675),
.A2(n_5458),
.B1(n_5459),
.B2(n_5457),
.Y(n_15706)
);

INVx1_ASAP7_75t_L g15707 ( 
.A(n_15692),
.Y(n_15707)
);

INVx1_ASAP7_75t_L g15708 ( 
.A(n_15673),
.Y(n_15708)
);

INVx1_ASAP7_75t_L g15709 ( 
.A(n_15688),
.Y(n_15709)
);

AOI22xp5_ASAP7_75t_L g15710 ( 
.A1(n_15678),
.A2(n_6303),
.B1(n_6328),
.B2(n_6311),
.Y(n_15710)
);

INVx1_ASAP7_75t_L g15711 ( 
.A(n_15695),
.Y(n_15711)
);

AND2x4_ASAP7_75t_L g15712 ( 
.A(n_15679),
.B(n_5821),
.Y(n_15712)
);

INVx1_ASAP7_75t_L g15713 ( 
.A(n_15696),
.Y(n_15713)
);

OAI22xp5_ASAP7_75t_L g15714 ( 
.A1(n_15681),
.A2(n_6311),
.B1(n_6328),
.B2(n_6303),
.Y(n_15714)
);

INVx1_ASAP7_75t_L g15715 ( 
.A(n_15694),
.Y(n_15715)
);

INVx1_ASAP7_75t_L g15716 ( 
.A(n_15691),
.Y(n_15716)
);

OAI22xp5_ASAP7_75t_SL g15717 ( 
.A1(n_15668),
.A2(n_5458),
.B1(n_5459),
.B2(n_5457),
.Y(n_15717)
);

AOI22xp33_ASAP7_75t_L g15718 ( 
.A1(n_15685),
.A2(n_6328),
.B1(n_6311),
.B2(n_5459),
.Y(n_15718)
);

INVx1_ASAP7_75t_L g15719 ( 
.A(n_15682),
.Y(n_15719)
);

AOI22xp5_ASAP7_75t_L g15720 ( 
.A1(n_15670),
.A2(n_6328),
.B1(n_6331),
.B2(n_6177),
.Y(n_15720)
);

AOI22xp5_ASAP7_75t_L g15721 ( 
.A1(n_15666),
.A2(n_6328),
.B1(n_6333),
.B2(n_6331),
.Y(n_15721)
);

OAI22x1_ASAP7_75t_L g15722 ( 
.A1(n_15680),
.A2(n_6257),
.B1(n_6258),
.B2(n_6047),
.Y(n_15722)
);

INVx1_ASAP7_75t_L g15723 ( 
.A(n_15660),
.Y(n_15723)
);

AOI22xp5_ASAP7_75t_L g15724 ( 
.A1(n_15667),
.A2(n_15684),
.B1(n_15665),
.B2(n_15662),
.Y(n_15724)
);

OAI22xp5_ASAP7_75t_L g15725 ( 
.A1(n_15683),
.A2(n_6258),
.B1(n_6257),
.B2(n_5458),
.Y(n_15725)
);

BUFx2_ASAP7_75t_L g15726 ( 
.A(n_15661),
.Y(n_15726)
);

AO22x2_ASAP7_75t_L g15727 ( 
.A1(n_15669),
.A2(n_5514),
.B1(n_5540),
.B2(n_5455),
.Y(n_15727)
);

OAI22x1_ASAP7_75t_L g15728 ( 
.A1(n_15669),
.A2(n_6258),
.B1(n_6257),
.B2(n_5878),
.Y(n_15728)
);

INVx1_ASAP7_75t_SL g15729 ( 
.A(n_15674),
.Y(n_15729)
);

OAI22xp5_ASAP7_75t_L g15730 ( 
.A1(n_15669),
.A2(n_6258),
.B1(n_6257),
.B2(n_5458),
.Y(n_15730)
);

AOI22xp5_ASAP7_75t_L g15731 ( 
.A1(n_15671),
.A2(n_6337),
.B1(n_6333),
.B2(n_5458),
.Y(n_15731)
);

AOI211xp5_ASAP7_75t_SL g15732 ( 
.A1(n_15674),
.A2(n_6364),
.B(n_6186),
.C(n_6189),
.Y(n_15732)
);

NOR4xp25_ASAP7_75t_SL g15733 ( 
.A(n_15726),
.B(n_6221),
.C(n_6265),
.D(n_6200),
.Y(n_15733)
);

NOR2x1_ASAP7_75t_L g15734 ( 
.A(n_15702),
.B(n_5458),
.Y(n_15734)
);

NAND2xp5_ASAP7_75t_L g15735 ( 
.A(n_15729),
.B(n_5821),
.Y(n_15735)
);

INVx1_ASAP7_75t_L g15736 ( 
.A(n_15703),
.Y(n_15736)
);

NOR2xp67_ASAP7_75t_L g15737 ( 
.A(n_15700),
.B(n_5458),
.Y(n_15737)
);

XNOR2xp5_ASAP7_75t_SL g15738 ( 
.A(n_15697),
.B(n_5959),
.Y(n_15738)
);

NOR3xp33_ASAP7_75t_L g15739 ( 
.A(n_15707),
.B(n_15708),
.C(n_15709),
.Y(n_15739)
);

NAND2xp5_ASAP7_75t_L g15740 ( 
.A(n_15711),
.B(n_15699),
.Y(n_15740)
);

INVx1_ASAP7_75t_L g15741 ( 
.A(n_15698),
.Y(n_15741)
);

INVx2_ASAP7_75t_L g15742 ( 
.A(n_15701),
.Y(n_15742)
);

AOI221xp5_ASAP7_75t_L g15743 ( 
.A1(n_15704),
.A2(n_5459),
.B1(n_5479),
.B2(n_5475),
.C(n_5458),
.Y(n_15743)
);

OAI322xp33_ASAP7_75t_L g15744 ( 
.A1(n_15719),
.A2(n_6359),
.A3(n_6347),
.B1(n_5479),
.B2(n_5487),
.C1(n_5459),
.C2(n_5492),
.Y(n_15744)
);

INVx2_ASAP7_75t_L g15745 ( 
.A(n_15723),
.Y(n_15745)
);

INVx1_ASAP7_75t_L g15746 ( 
.A(n_15724),
.Y(n_15746)
);

NAND4xp25_ASAP7_75t_L g15747 ( 
.A(n_15705),
.B(n_5266),
.C(n_5286),
.D(n_5243),
.Y(n_15747)
);

AND2x2_ASAP7_75t_SL g15748 ( 
.A(n_15713),
.B(n_5459),
.Y(n_15748)
);

NAND2xp5_ASAP7_75t_L g15749 ( 
.A(n_15716),
.B(n_5878),
.Y(n_15749)
);

NOR2x1_ASAP7_75t_L g15750 ( 
.A(n_15715),
.B(n_5459),
.Y(n_15750)
);

OAI22xp5_ASAP7_75t_L g15751 ( 
.A1(n_15731),
.A2(n_5459),
.B1(n_5479),
.B2(n_5475),
.Y(n_15751)
);

NAND4xp25_ASAP7_75t_L g15752 ( 
.A(n_15712),
.B(n_5266),
.C(n_5286),
.D(n_5243),
.Y(n_15752)
);

NOR4xp25_ASAP7_75t_L g15753 ( 
.A(n_15725),
.B(n_6462),
.C(n_6468),
.D(n_6467),
.Y(n_15753)
);

XNOR2xp5_ASAP7_75t_L g15754 ( 
.A(n_15721),
.B(n_6424),
.Y(n_15754)
);

NAND3xp33_ASAP7_75t_L g15755 ( 
.A(n_15720),
.B(n_5370),
.C(n_5321),
.Y(n_15755)
);

AOI22xp33_ASAP7_75t_L g15756 ( 
.A1(n_15706),
.A2(n_5479),
.B1(n_5487),
.B2(n_5475),
.Y(n_15756)
);

AND2x4_ASAP7_75t_L g15757 ( 
.A(n_15735),
.B(n_15710),
.Y(n_15757)
);

INVx1_ASAP7_75t_L g15758 ( 
.A(n_15740),
.Y(n_15758)
);

XNOR2xp5_ASAP7_75t_L g15759 ( 
.A(n_15741),
.B(n_15717),
.Y(n_15759)
);

INVx2_ASAP7_75t_L g15760 ( 
.A(n_15742),
.Y(n_15760)
);

AND2x4_ASAP7_75t_L g15761 ( 
.A(n_15739),
.B(n_15718),
.Y(n_15761)
);

NOR2x2_ASAP7_75t_L g15762 ( 
.A(n_15745),
.B(n_15732),
.Y(n_15762)
);

AOI22xp5_ASAP7_75t_L g15763 ( 
.A1(n_15746),
.A2(n_15714),
.B1(n_15730),
.B2(n_15727),
.Y(n_15763)
);

NAND3xp33_ASAP7_75t_SL g15764 ( 
.A(n_15736),
.B(n_15722),
.C(n_15727),
.Y(n_15764)
);

OR2x2_ASAP7_75t_L g15765 ( 
.A(n_15749),
.B(n_15728),
.Y(n_15765)
);

NOR3xp33_ASAP7_75t_L g15766 ( 
.A(n_15737),
.B(n_5357),
.C(n_5315),
.Y(n_15766)
);

INVx2_ASAP7_75t_L g15767 ( 
.A(n_15750),
.Y(n_15767)
);

XNOR2xp5_ASAP7_75t_L g15768 ( 
.A(n_15738),
.B(n_6424),
.Y(n_15768)
);

INVx1_ASAP7_75t_L g15769 ( 
.A(n_15734),
.Y(n_15769)
);

OAI221xp5_ASAP7_75t_SL g15770 ( 
.A1(n_15747),
.A2(n_6359),
.B1(n_6347),
.B2(n_6176),
.C(n_6154),
.Y(n_15770)
);

OAI22xp5_ASAP7_75t_L g15771 ( 
.A1(n_15760),
.A2(n_15748),
.B1(n_15755),
.B2(n_15754),
.Y(n_15771)
);

XOR2xp5_ASAP7_75t_L g15772 ( 
.A(n_15758),
.B(n_15759),
.Y(n_15772)
);

AOI21xp5_ASAP7_75t_L g15773 ( 
.A1(n_15761),
.A2(n_15752),
.B(n_15753),
.Y(n_15773)
);

OAI22x1_ASAP7_75t_SL g15774 ( 
.A1(n_15769),
.A2(n_15733),
.B1(n_15743),
.B2(n_15751),
.Y(n_15774)
);

BUFx6f_ASAP7_75t_L g15775 ( 
.A(n_15767),
.Y(n_15775)
);

OAI22xp5_ASAP7_75t_L g15776 ( 
.A1(n_15765),
.A2(n_15756),
.B1(n_15744),
.B2(n_5475),
.Y(n_15776)
);

AOI22x1_ASAP7_75t_L g15777 ( 
.A1(n_15757),
.A2(n_5479),
.B1(n_5489),
.B2(n_5487),
.Y(n_15777)
);

XOR2xp5_ASAP7_75t_L g15778 ( 
.A(n_15763),
.B(n_5475),
.Y(n_15778)
);

AOI21x1_ASAP7_75t_L g15779 ( 
.A1(n_15762),
.A2(n_5453),
.B(n_5878),
.Y(n_15779)
);

AOI21xp33_ASAP7_75t_L g15780 ( 
.A1(n_15764),
.A2(n_5370),
.B(n_5321),
.Y(n_15780)
);

AOI22xp5_ASAP7_75t_L g15781 ( 
.A1(n_15768),
.A2(n_5636),
.B1(n_5774),
.B2(n_5475),
.Y(n_15781)
);

OAI31xp33_ASAP7_75t_SL g15782 ( 
.A1(n_15766),
.A2(n_6166),
.A3(n_6370),
.B(n_6100),
.Y(n_15782)
);

OAI22xp5_ASAP7_75t_L g15783 ( 
.A1(n_15778),
.A2(n_15770),
.B1(n_5475),
.B2(n_5487),
.Y(n_15783)
);

NAND3xp33_ASAP7_75t_L g15784 ( 
.A(n_15775),
.B(n_5370),
.C(n_5321),
.Y(n_15784)
);

AOI21xp5_ASAP7_75t_L g15785 ( 
.A1(n_15772),
.A2(n_5453),
.B(n_5475),
.Y(n_15785)
);

INVxp67_ASAP7_75t_L g15786 ( 
.A(n_15775),
.Y(n_15786)
);

OAI22xp33_ASAP7_75t_SL g15787 ( 
.A1(n_15771),
.A2(n_6389),
.B1(n_6312),
.B2(n_6290),
.Y(n_15787)
);

INVx1_ASAP7_75t_SL g15788 ( 
.A(n_15773),
.Y(n_15788)
);

OAI22xp5_ASAP7_75t_L g15789 ( 
.A1(n_15776),
.A2(n_15780),
.B1(n_15781),
.B2(n_15774),
.Y(n_15789)
);

AOI22xp33_ASAP7_75t_L g15790 ( 
.A1(n_15777),
.A2(n_5479),
.B1(n_5487),
.B2(n_5475),
.Y(n_15790)
);

INVx2_ASAP7_75t_L g15791 ( 
.A(n_15779),
.Y(n_15791)
);

NAND2xp5_ASAP7_75t_L g15792 ( 
.A(n_15786),
.B(n_15782),
.Y(n_15792)
);

NAND2xp5_ASAP7_75t_L g15793 ( 
.A(n_15788),
.B(n_5479),
.Y(n_15793)
);

O2A1O1Ixp33_ASAP7_75t_L g15794 ( 
.A1(n_15789),
.A2(n_5900),
.B(n_5943),
.C(n_5884),
.Y(n_15794)
);

OAI21x1_ASAP7_75t_L g15795 ( 
.A1(n_15792),
.A2(n_15791),
.B(n_15785),
.Y(n_15795)
);

XNOR2x1_ASAP7_75t_L g15796 ( 
.A(n_15793),
.B(n_15784),
.Y(n_15796)
);

NAND3xp33_ASAP7_75t_L g15797 ( 
.A(n_15796),
.B(n_15783),
.C(n_15790),
.Y(n_15797)
);

NAND2xp5_ASAP7_75t_L g15798 ( 
.A(n_15795),
.B(n_15794),
.Y(n_15798)
);

AOI22xp5_ASAP7_75t_L g15799 ( 
.A1(n_15797),
.A2(n_15787),
.B1(n_5479),
.B2(n_5489),
.Y(n_15799)
);

AOI22xp33_ASAP7_75t_L g15800 ( 
.A1(n_15798),
.A2(n_5487),
.B1(n_5489),
.B2(n_5479),
.Y(n_15800)
);

OAI21xp5_ASAP7_75t_L g15801 ( 
.A1(n_15799),
.A2(n_15800),
.B(n_5453),
.Y(n_15801)
);

OAI221xp5_ASAP7_75t_R g15802 ( 
.A1(n_15801),
.A2(n_5798),
.B1(n_6097),
.B2(n_6656),
.C(n_5653),
.Y(n_15802)
);

AOI22xp33_ASAP7_75t_L g15803 ( 
.A1(n_15802),
.A2(n_5487),
.B1(n_5489),
.B2(n_5479),
.Y(n_15803)
);

AOI211xp5_ASAP7_75t_L g15804 ( 
.A1(n_15803),
.A2(n_5487),
.B(n_5492),
.C(n_5489),
.Y(n_15804)
);


endmodule