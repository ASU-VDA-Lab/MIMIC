module fake_jpeg_5627_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_38),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_39),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g47 ( 
.A(n_29),
.B(n_2),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_23),
.CI(n_31),
.CON(n_78),
.SN(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_57),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_32),
.B1(n_19),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_68),
.B1(n_70),
.B2(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_58),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_72),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_26),
.B1(n_16),
.B2(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_78),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_28),
.B1(n_31),
.B2(n_21),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_24),
.B(n_14),
.C(n_23),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_103),
.B(n_67),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_31),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_100),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_24),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_22),
.B(n_24),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_78),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_111),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_56),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_116),
.B(n_119),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_52),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_79),
.B1(n_53),
.B2(n_71),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_91),
.B1(n_102),
.B2(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_14),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_79),
.B1(n_71),
.B2(n_64),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_125),
.B1(n_80),
.B2(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_76),
.B1(n_24),
.B2(n_14),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_128),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_115),
.B1(n_108),
.B2(n_122),
.Y(n_152)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_96),
.A3(n_80),
.B1(n_97),
.B2(n_103),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_137),
.B1(n_109),
.B2(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_80),
.B1(n_84),
.B2(n_76),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_107),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_113),
.B1(n_80),
.B2(n_124),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_143),
.B(n_123),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_108),
.C(n_95),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_90),
.B1(n_14),
.B2(n_93),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_105),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_134),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_109),
.B(n_117),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_150),
.B(n_82),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_137),
.B1(n_128),
.B2(n_140),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_142),
.C(n_135),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_112),
.B(n_105),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_134),
.B(n_129),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_160),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_166),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_135),
.C(n_126),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_133),
.B(n_143),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_151),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_93),
.C(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_152),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_93),
.B(n_22),
.C(n_5),
.D(n_6),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_149),
.C(n_148),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_170),
.B(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_173),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_159),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_164),
.B(n_165),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_178),
.B(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_110),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_147),
.B(n_167),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_151),
.B(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_173),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_182),
.C(n_13),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_107),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_8),
.C(n_9),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_175),
.A3(n_172),
.B1(n_158),
.B2(n_154),
.C1(n_144),
.C2(n_12),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_186),
.C(n_13),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);


endmodule