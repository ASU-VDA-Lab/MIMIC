module fake_aes_8579_n_25 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_7;
BUFx10_ASAP7_75t_L g7 ( .A(n_2), .Y(n_7) );
INVx1_ASAP7_75t_SL g8 ( .A(n_3), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
AND2x2_ASAP7_75t_SL g10 ( .A(n_0), .B(n_5), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_1), .B(n_0), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_2), .B(n_3), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_1), .B(n_4), .Y(n_14) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_9), .A2(n_5), .B(n_6), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_9), .A2(n_6), .B(n_12), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_13), .B(n_7), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_16), .B(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_14), .B(n_15), .Y(n_21) );
AOI211xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_18), .B(n_8), .C(n_15), .Y(n_22) );
AOI211xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_18), .B(n_8), .C(n_12), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_7), .B1(n_10), .B2(n_22), .Y(n_24) );
OAI211xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_10), .B(n_23), .C(n_22), .Y(n_25) );
endmodule