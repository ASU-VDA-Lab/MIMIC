module fake_jpeg_22546_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_18),
.C(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_42),
.B1(n_33),
.B2(n_14),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_21),
.B1(n_24),
.B2(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_40),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_75),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_33),
.B1(n_42),
.B2(n_51),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_67),
.B1(n_50),
.B2(n_49),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_16),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_51),
.B1(n_69),
.B2(n_46),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_72),
.B1(n_68),
.B2(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_75),
.B1(n_59),
.B2(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_22),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.C(n_87),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_41),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_35),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_42),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_12),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_119),
.B1(n_93),
.B2(n_46),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_90),
.B(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_108),
.B1(n_114),
.B2(n_80),
.Y(n_129)
);

AO21x2_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_71),
.B(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_109),
.B1(n_93),
.B2(n_83),
.Y(n_131)
);

BUFx4f_ASAP7_75t_SL g107 ( 
.A(n_83),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_50),
.B1(n_49),
.B2(n_34),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_34),
.B1(n_29),
.B2(n_63),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_116),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_14),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_117),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_58),
.B1(n_38),
.B2(n_53),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_85),
.C(n_90),
.Y(n_126)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_91),
.C(n_87),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_128),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_130),
.C(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_96),
.C(n_80),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_140),
.Y(n_165)
);

OAI22x1_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_71),
.B1(n_43),
.B2(n_44),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_70),
.B(n_57),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_76),
.B(n_25),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_37),
.C(n_28),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_122),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_25),
.B(n_19),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_100),
.B(n_112),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_105),
.B(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_162),
.B1(n_168),
.B2(n_144),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_159),
.B1(n_163),
.B2(n_169),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_162)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_119),
.B1(n_45),
.B2(n_73),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_73),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_138),
.C(n_130),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_186),
.C(n_187),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_131),
.B(n_129),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_163),
.B(n_164),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_123),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_184),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_167),
.B1(n_163),
.B2(n_168),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_126),
.C(n_142),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_134),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_120),
.C(n_141),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_157),
.C(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_137),
.B(n_12),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_11),
.C(n_19),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_169),
.B1(n_145),
.B2(n_156),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_208),
.B1(n_184),
.B2(n_174),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_152),
.B1(n_162),
.B2(n_145),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_202),
.B1(n_207),
.B2(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_157),
.B1(n_167),
.B2(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_213),
.C(n_214),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_188),
.B1(n_181),
.B2(n_191),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_216),
.B(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_150),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_176),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_45),
.B1(n_70),
.B2(n_57),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_36),
.C(n_28),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_36),
.C(n_28),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_11),
.B(n_1),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_228),
.B1(n_214),
.B2(n_210),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_223),
.B(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_174),
.B1(n_195),
.B2(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_231),
.B1(n_220),
.B2(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_183),
.C(n_172),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_229),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_177),
.B1(n_45),
.B2(n_36),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_177),
.C(n_45),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_207),
.B1(n_203),
.B2(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_22),
.C(n_23),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_22),
.C(n_23),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_241),
.B1(n_221),
.B2(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_217),
.B1(n_11),
.B2(n_23),
.Y(n_241)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_218),
.B(n_0),
.C(n_2),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_22),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_235),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_0),
.Y(n_250)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_0),
.B(n_2),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_263),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_27),
.B1(n_15),
.B2(n_4),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_253),
.B1(n_249),
.B2(n_248),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_225),
.CI(n_27),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_22),
.C(n_23),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_268),
.C(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_27),
.B1(n_15),
.B2(n_4),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_246),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_27),
.C(n_15),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_256),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_269),
.A2(n_280),
.B1(n_261),
.B2(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_276),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_243),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_255),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_19),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_268),
.B(n_263),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_2),
.C(n_3),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_285),
.B1(n_280),
.B2(n_269),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_272),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_5),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_289),
.C(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_295),
.B(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_294),
.B(n_7),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_287),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_290),
.C(n_293),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_295),
.C(n_291),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_299),
.B(n_9),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_8),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_10),
.B(n_297),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_10),
.Y(n_305)
);


endmodule