module fake_jpeg_9358_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx5p33_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_16),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_11),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_6),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_20),
.B1(n_9),
.B2(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_15),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_10),
.B1(n_18),
.B2(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_25),
.C(n_14),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_23),
.C(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_28),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_37),
.C(n_33),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_30),
.C(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_17),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_26),
.C(n_8),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_8),
.B(n_41),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);


endmodule