module fake_ariane_1869_n_1685 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1685);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1685;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_25),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_10),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_65),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_8),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_35),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_44),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_97),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_23),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_7),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_40),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_64),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_32),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_140),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_136),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_53),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_17),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_54),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_3),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_21),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_92),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_17),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_34),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_33),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_19),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_113),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_68),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_19),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_80),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_69),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_125),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_122),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_123),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_145),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_142),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_101),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_50),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_46),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_28),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_50),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_43),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_139),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_16),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_148),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_147),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_32),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_99),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_112),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_55),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_86),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_9),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_31),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_37),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_45),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_151),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_126),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_124),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_59),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_138),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_115),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_22),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_78),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_23),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_40),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_116),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_67),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_60),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_41),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_95),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_9),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_146),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_105),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_178),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_152),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_194),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_170),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_180),
.B(n_1),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_180),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_246),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_211),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_199),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_247),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_184),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_187),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_271),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_187),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_184),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_201),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_157),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_201),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_189),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_199),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_212),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_212),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_228),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_204),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_234),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_234),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_164),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_243),
.B(n_4),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_217),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_287),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_204),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_204),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_260),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_182),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_227),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_161),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_183),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_288),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_291),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_5),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_204),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_296),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_198),
.B(n_205),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_204),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_161),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_169),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_190),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_154),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_154),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_169),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_163),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_210),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_169),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_R g377 ( 
.A(n_153),
.B(n_149),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_163),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_165),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_198),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_205),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_305),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_313),
.B(n_237),
.Y(n_394)
);

NAND2x1p5_ASAP7_75t_L g395 ( 
.A(n_314),
.B(n_185),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_197),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_308),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_337),
.B(n_237),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_369),
.B(n_209),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_215),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_299),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_330),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_335),
.A2(n_224),
.B(n_209),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_233),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_344),
.B(n_256),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_224),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_357),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_359),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_312),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_268),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_315),
.Y(n_443)
);

BUFx12f_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_365),
.B(n_277),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_320),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_302),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_394),
.A2(n_313),
.B1(n_350),
.B2(n_353),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_343),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_447),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_395),
.A2(n_350),
.B1(n_375),
.B2(n_356),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_395),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_426),
.B(n_368),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_415),
.B(n_320),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

INVx8_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_341),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_405),
.B(n_333),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_379),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_415),
.B(n_306),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_332),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_371),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_395),
.A2(n_316),
.B1(n_358),
.B2(n_216),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_425),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_388),
.B(n_226),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_396),
.B(n_322),
.Y(n_478)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_332),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_395),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_299),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_385),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_332),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_372),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_327),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_266),
.B1(n_219),
.B2(n_285),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_374),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_385),
.B(n_374),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_449),
.B(n_309),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_386),
.B(n_378),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_421),
.Y(n_497)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_386),
.B(n_378),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_449),
.B(n_380),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_446),
.Y(n_504)
);

BUFx4f_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_408),
.B(n_311),
.Y(n_506)
);

XOR2x2_ASAP7_75t_SL g507 ( 
.A(n_400),
.B(n_345),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_377),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_400),
.B(n_165),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_390),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_396),
.B(n_158),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_429),
.B(n_159),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_394),
.B(n_319),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_429),
.B(n_160),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_409),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_390),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_400),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_440),
.B(n_321),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_384),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_L g526 ( 
.A(n_409),
.B(n_156),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_391),
.B(n_226),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_402),
.B(n_318),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_400),
.B(n_406),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_444),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_406),
.B(n_410),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_402),
.B(n_373),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_427),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_406),
.B(n_155),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_384),
.B(n_376),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_387),
.B(n_323),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_427),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_387),
.B(n_325),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_434),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_406),
.A2(n_293),
.B1(n_297),
.B2(n_242),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_434),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_406),
.B(n_230),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_410),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

BUFx4f_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_391),
.B(n_155),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_416),
.A2(n_293),
.B1(n_297),
.B2(n_167),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_443),
.B(n_222),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_437),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_410),
.B(n_411),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_410),
.B(n_411),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_405),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_437),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_399),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

AND2x6_ASAP7_75t_L g573 ( 
.A(n_445),
.B(n_290),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_439),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_392),
.B(n_397),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_410),
.B(n_232),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_392),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_397),
.B(n_167),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_398),
.B(n_155),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_398),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_411),
.B(n_162),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_411),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_383),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_416),
.B(n_290),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_411),
.B(n_166),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_442),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_418),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_442),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_401),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_418),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_418),
.B(n_168),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_442),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_401),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_442),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_418),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_501),
.B(n_418),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_466),
.B(n_424),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_457),
.B(n_424),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_478),
.B(n_424),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_509),
.B(n_424),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_540),
.B(n_424),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_467),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_478),
.B(n_403),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_458),
.B(n_484),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_454),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_538),
.B(n_403),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_471),
.B(n_404),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_513),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_474),
.B(n_404),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_471),
.B(n_407),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_471),
.B(n_407),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_412),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_451),
.B(n_459),
.C(n_571),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_451),
.A2(n_432),
.B1(n_445),
.B2(n_438),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_412),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_460),
.A2(n_414),
.B(n_413),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_458),
.B(n_413),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_530),
.B(n_383),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_419),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_469),
.B(n_414),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_586),
.A2(n_416),
.B1(n_428),
.B2(n_423),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_580),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_546),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_473),
.A2(n_417),
.B1(n_438),
.B2(n_436),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_592),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_596),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_484),
.B(n_417),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_581),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_482),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_552),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_571),
.B(n_420),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_482),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_546),
.B(n_405),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_523),
.B(n_420),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_521),
.B(n_422),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_574),
.B(n_431),
.C(n_422),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_575),
.A2(n_593),
.B(n_589),
.C(n_579),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_497),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_530),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_515),
.B(n_516),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_574),
.B(n_431),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_569),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_492),
.B(n_435),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_581),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_488),
.A2(n_435),
.B1(n_436),
.B2(n_273),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_492),
.B(n_441),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_543),
.B(n_419),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_569),
.B(n_352),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_491),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_586),
.A2(n_416),
.B1(n_433),
.B2(n_430),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_450),
.B(n_441),
.C(n_433),
.Y(n_669)
);

BUFx5_ASAP7_75t_L g670 ( 
.A(n_475),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_557),
.B(n_419),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_579),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_488),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_495),
.B(n_423),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_488),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_518),
.B(n_529),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_483),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_493),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_560),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_529),
.B(n_489),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_496),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_494),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_492),
.B(n_537),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_499),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_534),
.B(n_423),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_494),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_578),
.B(n_428),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_563),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_564),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_428),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_578),
.B(n_430),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_578),
.B(n_430),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_537),
.B(n_433),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_531),
.B(n_441),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_475),
.A2(n_416),
.B1(n_382),
.B2(n_171),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_512),
.B(n_236),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_486),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_512),
.B(n_382),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_475),
.A2(n_269),
.B1(n_171),
.B2(n_172),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_560),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_472),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_512),
.B(n_249),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_485),
.Y(n_703)
);

BUFx6f_ASAP7_75t_SL g704 ( 
.A(n_485),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_585),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_464),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_463),
.B(n_251),
.Y(n_707)
);

INVx4_ASAP7_75t_SL g708 ( 
.A(n_475),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_481),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_487),
.Y(n_710)
);

BUFx6f_ASAP7_75t_SL g711 ( 
.A(n_485),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_549),
.B(n_470),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_485),
.B(n_355),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_528),
.B(n_517),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_576),
.B(n_172),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_453),
.B(n_254),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_559),
.B(n_173),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_476),
.Y(n_718)
);

AND2x4_ASAP7_75t_SL g719 ( 
.A(n_565),
.B(n_360),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_583),
.B(n_173),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_587),
.B(n_174),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_476),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_453),
.B(n_479),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_594),
.B(n_255),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_475),
.A2(n_265),
.B1(n_245),
.B2(n_244),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_472),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_472),
.B(n_174),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_477),
.B(n_175),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_506),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_514),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_507),
.A2(n_261),
.B1(n_177),
.B2(n_301),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_480),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_477),
.B(n_175),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_477),
.B(n_177),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_565),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_456),
.B(n_262),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_480),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_490),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_510),
.B(n_181),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_475),
.A2(n_527),
.B1(n_573),
.B2(n_462),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_464),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_507),
.B(n_363),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_527),
.B(n_181),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_524),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_524),
.B(n_156),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_519),
.B(n_272),
.C(n_274),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_510),
.B(n_206),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_527),
.A2(n_273),
.B1(n_301),
.B2(n_242),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_510),
.B(n_206),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_462),
.B(n_248),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_532),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_533),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_527),
.A2(n_186),
.B1(n_188),
.B2(n_295),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_453),
.B(n_156),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_479),
.B(n_156),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_479),
.B(n_156),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_527),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_532),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_533),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_522),
.B(n_544),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_535),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_522),
.B(n_248),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_535),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_608),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_662),
.B(n_456),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_672),
.A2(n_527),
.B1(n_573),
.B2(n_541),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_656),
.A2(n_597),
.B(n_536),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_606),
.A2(n_597),
.B(n_558),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_611),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_616),
.B(n_573),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_616),
.B(n_664),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_662),
.B(n_607),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_760),
.A2(n_548),
.B(n_536),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_605),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_664),
.B(n_573),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_602),
.A2(n_547),
.B(n_548),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_607),
.B(n_456),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_738),
.B(n_519),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_679),
.B(n_364),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_606),
.A2(n_547),
.B(n_554),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_685),
.B(n_573),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_601),
.A2(n_554),
.B(n_558),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_626),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_620),
.A2(n_562),
.B(n_591),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_598),
.A2(n_562),
.B(n_591),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_685),
.B(n_573),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_618),
.B(n_522),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_653),
.A2(n_252),
.B(n_282),
.C(n_275),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_544),
.Y(n_793)
);

BUFx4f_ASAP7_75t_SL g794 ( 
.A(n_655),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_598),
.A2(n_595),
.B(n_542),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_623),
.A2(n_595),
.B(n_542),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_676),
.A2(n_545),
.B(n_553),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_621),
.B(n_544),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_670),
.B(n_456),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_519),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_613),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_709),
.A2(n_550),
.B(n_553),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_672),
.A2(n_539),
.B1(n_541),
.B2(n_555),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_700),
.B(n_252),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_631),
.A2(n_668),
.B(n_636),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_680),
.A2(n_257),
.B(n_261),
.C(n_269),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_710),
.A2(n_550),
.B(n_545),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_604),
.A2(n_257),
.B(n_275),
.C(n_282),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_658),
.B(n_263),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_621),
.B(n_561),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_671),
.B(n_561),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_614),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_561),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_678),
.B(n_582),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_613),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_613),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_627),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_636),
.A2(n_567),
.B(n_566),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_699),
.B(n_500),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_697),
.A2(n_570),
.B(n_567),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_635),
.A2(n_572),
.B(n_570),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_617),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_703),
.B(n_462),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_660),
.A2(n_572),
.B(n_568),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_681),
.B(n_582),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_666),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_684),
.B(n_582),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_628),
.A2(n_651),
.B(n_663),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_693),
.A2(n_568),
.B(n_566),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_619),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_632),
.A2(n_539),
.B1(n_541),
.B2(n_555),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_652),
.A2(n_590),
.B(n_588),
.C(n_526),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_645),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_609),
.B(n_588),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_632),
.A2(n_539),
.B1(n_555),
.B2(n_588),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_642),
.A2(n_590),
.B(n_456),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_670),
.B(n_465),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_714),
.B(n_590),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_652),
.B(n_465),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_622),
.B(n_465),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_642),
.A2(n_465),
.B(n_500),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_634),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_R g844 ( 
.A(n_633),
.B(n_462),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_694),
.A2(n_556),
.B(n_505),
.C(n_502),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_648),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_650),
.B(n_465),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_667),
.A2(n_556),
.B(n_505),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_634),
.Y(n_849)
);

OAI321xp33_ASAP7_75t_L g850 ( 
.A1(n_699),
.A2(n_276),
.A3(n_284),
.B1(n_286),
.B2(n_294),
.C(n_298),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_716),
.A2(n_556),
.B(n_505),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_729),
.B(n_498),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_677),
.A2(n_502),
.B(n_500),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_650),
.B(n_498),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_624),
.A2(n_498),
.B1(n_502),
.B2(n_526),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_703),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_718),
.A2(n_292),
.B(n_283),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_722),
.A2(n_281),
.B(n_176),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_732),
.A2(n_225),
.B(n_279),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_674),
.B(n_280),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_615),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_629),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_694),
.A2(n_223),
.B(n_278),
.C(n_270),
.Y(n_863)
);

AO21x1_ASAP7_75t_L g864 ( 
.A1(n_754),
.A2(n_280),
.B(n_91),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_630),
.B(n_637),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_640),
.B(n_280),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_647),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_737),
.A2(n_267),
.B(n_253),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_751),
.A2(n_250),
.B(n_241),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_687),
.A2(n_692),
.B1(n_691),
.B2(n_641),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_657),
.A2(n_683),
.B(n_720),
.C(n_721),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_724),
.B(n_240),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_624),
.A2(n_239),
.B1(n_238),
.B2(n_235),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_615),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_724),
.A2(n_231),
.B1(n_229),
.B2(n_221),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_758),
.A2(n_220),
.B(n_214),
.Y(n_876)
);

AND2x2_ASAP7_75t_SL g877 ( 
.A(n_748),
.B(n_11),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_627),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_627),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_690),
.A2(n_213),
.B(n_208),
.C(n_203),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_639),
.B(n_202),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_690),
.A2(n_200),
.B(n_196),
.C(n_195),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_670),
.B(n_193),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_729),
.B(n_13),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_698),
.B(n_179),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_723),
.A2(n_52),
.B(n_131),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_682),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_719),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_686),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_688),
.B(n_14),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_627),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_689),
.B(n_14),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_705),
.B(n_20),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_703),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_670),
.B(n_20),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_649),
.B(n_21),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_707),
.B(n_26),
.C(n_27),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_750),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_727),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_643),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_670),
.B(n_654),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_701),
.A2(n_71),
.B(n_119),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_670),
.B(n_30),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_701),
.A2(n_70),
.B(n_118),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_728),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_654),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_673),
.B(n_36),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_696),
.B(n_36),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_750),
.B(n_38),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_754),
.A2(n_75),
.B(n_111),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_669),
.A2(n_39),
.B(n_41),
.C(n_44),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_654),
.B(n_47),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_675),
.B(n_48),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_644),
.B(n_49),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_733),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_734),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_739),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_668),
.A2(n_88),
.B(n_106),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_726),
.A2(n_85),
.B(n_104),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_746),
.A2(n_49),
.B1(n_51),
.B2(n_58),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_742),
.B(n_135),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_661),
.B(n_79),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_743),
.B(n_715),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_731),
.A2(n_93),
.B(n_712),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_603),
.A2(n_763),
.B(n_744),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_743),
.B(n_612),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_755),
.A2(n_756),
.B(n_761),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_702),
.A2(n_762),
.B(n_749),
.C(n_747),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_730),
.A2(n_752),
.B(n_759),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_646),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_659),
.Y(n_931)
);

NOR2x1p5_ASAP7_75t_L g932 ( 
.A(n_735),
.B(n_711),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_665),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_746),
.A2(n_625),
.B(n_748),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_731),
.B(n_741),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_713),
.B(n_610),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_740),
.B(n_610),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_612),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_731),
.B(n_717),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_750),
.B(n_695),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_755),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_757),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_736),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_695),
.B(n_725),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_846),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_774),
.B(n_706),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_775),
.A2(n_756),
.B(n_740),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_775),
.A2(n_753),
.B(n_708),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_786),
.B(n_704),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_767),
.B(n_704),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_861),
.B(n_711),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_794),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_846),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_861),
.B(n_708),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_884),
.B(n_708),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_934),
.A2(n_745),
.B(n_800),
.C(n_781),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_773),
.A2(n_745),
.B(n_780),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_764),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_781),
.A2(n_800),
.B(n_829),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_794),
.B(n_745),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_877),
.A2(n_745),
.B1(n_935),
.B2(n_782),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_877),
.A2(n_820),
.B1(n_896),
.B2(n_908),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_827),
.B(n_936),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_895),
.A2(n_903),
.B(n_918),
.C(n_780),
.Y(n_964)
);

INVx3_ASAP7_75t_SL g965 ( 
.A(n_888),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_936),
.B(n_865),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_765),
.B(n_772),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_768),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_932),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_856),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_872),
.A2(n_944),
.B1(n_820),
.B2(n_854),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_908),
.B(n_897),
.C(n_874),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_812),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_809),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_771),
.A2(n_778),
.B(n_811),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_844),
.B(n_852),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_911),
.A2(n_871),
.B(n_880),
.C(n_882),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_823),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_898),
.B(n_814),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_898),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_924),
.A2(n_921),
.B1(n_940),
.B2(n_939),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_813),
.A2(n_788),
.B(n_805),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_824),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_831),
.B(n_862),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_900),
.B(n_914),
.C(n_882),
.Y(n_985)
);

BUFx8_ASAP7_75t_L g986 ( 
.A(n_893),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_814),
.B(n_843),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_840),
.A2(n_769),
.B1(n_793),
.B2(n_810),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_839),
.A2(n_897),
.B(n_867),
.C(n_928),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_843),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_797),
.A2(n_798),
.B(n_790),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_844),
.B(n_852),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_849),
.B(n_856),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_894),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_850),
.B(n_942),
.Y(n_995)
);

O2A1O1Ixp5_ASAP7_75t_L g996 ( 
.A1(n_895),
.A2(n_903),
.B(n_912),
.C(n_883),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_784),
.A2(n_789),
.B1(n_885),
.B2(n_870),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_875),
.A2(n_873),
.B1(n_766),
.B2(n_926),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_923),
.B(n_804),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_777),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_849),
.B(n_894),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_909),
.B(n_866),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_911),
.A2(n_880),
.B(n_792),
.C(n_808),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_795),
.A2(n_770),
.B(n_842),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_821),
.A2(n_783),
.B(n_847),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_796),
.A2(n_837),
.B(n_779),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_860),
.B(n_931),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_785),
.A2(n_802),
.B(n_807),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_816),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_933),
.B(n_930),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_899),
.B(n_905),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_824),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_881),
.B(n_938),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_878),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_766),
.A2(n_839),
.B1(n_942),
.B2(n_937),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_SL g1017 ( 
.A1(n_920),
.A2(n_907),
.B1(n_913),
.B2(n_892),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_824),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_835),
.A2(n_815),
.B1(n_828),
.B2(n_826),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_878),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_890),
.B(n_915),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_834),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_916),
.B(n_917),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_879),
.B(n_906),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_806),
.B(n_841),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_879),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_791),
.B(n_801),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_791),
.B(n_801),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_SL g1029 ( 
.A1(n_943),
.A2(n_883),
.B(n_901),
.C(n_799),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_887),
.B(n_889),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_816),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_863),
.A2(n_803),
.B(n_833),
.C(n_845),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_816),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_830),
.A2(n_776),
.B(n_845),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_863),
.B(n_906),
.Y(n_1035)
);

XOR2xp5_ASAP7_75t_L g1036 ( 
.A(n_816),
.B(n_818),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_799),
.A2(n_838),
.B(n_925),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_818),
.B(n_891),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_818),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_848),
.A2(n_855),
.B(n_922),
.C(n_853),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_818),
.B(n_891),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_836),
.A2(n_832),
.B(n_822),
.C(n_876),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_891),
.B(n_910),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_787),
.A2(n_825),
.B(n_838),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_819),
.A2(n_851),
.B(n_927),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_901),
.A2(n_929),
.B(n_919),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_891),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_941),
.B(n_857),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_858),
.B(n_859),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_868),
.A2(n_869),
.B(n_886),
.C(n_902),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_904),
.A2(n_774),
.B(n_775),
.C(n_616),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_864),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_774),
.B(n_503),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_927),
.A2(n_925),
.B(n_821),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_764),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_774),
.B(n_616),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_846),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_774),
.B(n_616),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_774),
.B(n_616),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_774),
.A2(n_775),
.B(n_616),
.Y(n_1060)
);

BUFx8_ASAP7_75t_SL g1061 ( 
.A(n_786),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_774),
.B(n_616),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_774),
.A2(n_607),
.B(n_616),
.C(n_775),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_774),
.A2(n_775),
.B(n_773),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_774),
.B(n_616),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_764),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_774),
.A2(n_775),
.B(n_773),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_774),
.A2(n_775),
.B(n_616),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_846),
.Y(n_1069)
);

OAI22x1_ASAP7_75t_L g1070 ( 
.A1(n_908),
.A2(n_464),
.B1(n_405),
.B2(n_457),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_774),
.A2(n_775),
.B(n_773),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_774),
.B(n_309),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_767),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_861),
.B(n_679),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_774),
.B(n_503),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_774),
.B(n_616),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_794),
.B(n_530),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_774),
.B(n_616),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_856),
.B(n_894),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_774),
.B(n_616),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_954),
.Y(n_1081)
);

INVx5_ASAP7_75t_L g1082 ( 
.A(n_1024),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1056),
.B(n_1058),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1063),
.A2(n_959),
.B(n_1051),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1051),
.A2(n_1068),
.B(n_1060),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1079),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1059),
.A2(n_1065),
.B(n_1062),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1072),
.A2(n_1080),
.B(n_1078),
.C(n_1076),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_966),
.B(n_1064),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_956),
.A2(n_1067),
.B(n_1064),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_972),
.A2(n_989),
.B(n_1053),
.C(n_1075),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_1049),
.A2(n_955),
.B(n_1050),
.C(n_992),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_962),
.B(n_985),
.C(n_977),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1067),
.A2(n_1071),
.B(n_975),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_973),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1071),
.A2(n_975),
.B(n_997),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_946),
.B(n_963),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1021),
.B(n_1012),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_964),
.B(n_982),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1034),
.A2(n_1044),
.B(n_1046),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_1007),
.A2(n_1045),
.B(n_1004),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1023),
.B(n_1008),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_983),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1073),
.B(n_974),
.Y(n_1105)
);

NOR2xp67_ASAP7_75t_L g1106 ( 
.A(n_949),
.B(n_951),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1052),
.A2(n_982),
.A3(n_1007),
.B(n_1004),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_962),
.B(n_998),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_1036),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_964),
.A2(n_988),
.B(n_947),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_980),
.B(n_1011),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1019),
.A2(n_1040),
.B(n_991),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1061),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1005),
.A2(n_1009),
.B(n_1046),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_953),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1037),
.A2(n_1009),
.B(n_1005),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1016),
.B(n_999),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_957),
.A2(n_1029),
.B(n_1042),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_952),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1015),
.Y(n_1120)
);

AO22x2_ASAP7_75t_L g1121 ( 
.A1(n_1014),
.A2(n_1070),
.B1(n_947),
.B2(n_948),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1057),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_967),
.B(n_984),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_957),
.A2(n_948),
.A3(n_1048),
.B(n_1069),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1042),
.A2(n_1032),
.B(n_976),
.Y(n_1125)
);

INVx3_ASAP7_75t_SL g1126 ( 
.A(n_969),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_978),
.B(n_1066),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_950),
.B(n_1002),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_996),
.A2(n_1032),
.B(n_977),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1003),
.A2(n_1025),
.B(n_961),
.C(n_995),
.Y(n_1130)
);

AND2x6_ASAP7_75t_L g1131 ( 
.A(n_983),
.B(n_1018),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1041),
.A2(n_1038),
.B(n_1035),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1006),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_SL g1135 ( 
.A1(n_1027),
.A2(n_1028),
.B(n_1047),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_965),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1017),
.A2(n_979),
.B1(n_1055),
.B2(n_1013),
.C(n_1018),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_968),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_970),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1000),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_981),
.A2(n_1030),
.B(n_1022),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1041),
.A2(n_1024),
.B(n_1039),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1020),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1024),
.B(n_1026),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_970),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_990),
.Y(n_1146)
);

NOR2xp67_ASAP7_75t_L g1147 ( 
.A(n_993),
.B(n_1001),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_1043),
.A2(n_987),
.B(n_960),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1039),
.B(n_1010),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1010),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1031),
.A2(n_1033),
.B(n_1039),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_986),
.A2(n_994),
.B1(n_1031),
.B2(n_1033),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1033),
.A2(n_994),
.B(n_986),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_SL g1154 ( 
.A(n_1072),
.B(n_530),
.C(n_972),
.Y(n_1154)
);

INVx6_ASAP7_75t_L g1155 ( 
.A(n_986),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_1034),
.A2(n_1007),
.B(n_1045),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_958),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1052),
.A2(n_982),
.A3(n_1007),
.B(n_1034),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1063),
.A2(n_774),
.B(n_775),
.C(n_1056),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1061),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_952),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1072),
.B(n_946),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_L g1165 ( 
.A1(n_972),
.A2(n_924),
.B1(n_1060),
.B2(n_1068),
.C(n_1063),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1074),
.B(n_638),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1052),
.A2(n_982),
.A3(n_1007),
.B(n_1034),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_945),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1077),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1056),
.B(n_1058),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1060),
.A2(n_1068),
.B1(n_1063),
.B2(n_775),
.C(n_774),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_958),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1079),
.B(n_814),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1063),
.A2(n_775),
.B(n_1051),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_958),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_1063),
.A2(n_774),
.B(n_775),
.C(n_1056),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_774),
.B(n_1068),
.C(n_1058),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_958),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_1052),
.B(n_982),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1074),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1060),
.A2(n_1068),
.B1(n_1063),
.B2(n_775),
.C(n_774),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1072),
.A2(n_464),
.B1(n_457),
.B2(n_405),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1063),
.A2(n_775),
.B(n_1051),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_945),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1060),
.A2(n_774),
.B(n_1068),
.C(n_1058),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_952),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_958),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_952),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1063),
.A2(n_775),
.B(n_1051),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1051),
.A2(n_977),
.B(n_1064),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1061),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1074),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_972),
.B(n_1072),
.C(n_962),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1044),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1056),
.B(n_1058),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1061),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1056),
.B(n_1058),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1079),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_774),
.B(n_959),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1204),
.A2(n_1094),
.B(n_1154),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1161),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1121),
.A2(n_1195),
.B1(n_1188),
.B2(n_1176),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1087),
.Y(n_1215)
);

BUFx4f_ASAP7_75t_L g1216 ( 
.A(n_1155),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1127),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1179),
.A2(n_1190),
.B1(n_1195),
.B2(n_1188),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1108),
.A2(n_1187),
.B1(n_1163),
.B2(n_1103),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1121),
.A2(n_1098),
.B1(n_1103),
.B2(n_1099),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1099),
.A2(n_1117),
.B1(n_1105),
.B2(n_1138),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1096),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1176),
.A2(n_1202),
.B1(n_1197),
.B2(n_1191),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1166),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1170),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1090),
.B(n_1123),
.Y(n_1226)
);

BUFx10_ASAP7_75t_L g1227 ( 
.A(n_1155),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1117),
.A2(n_1110),
.B1(n_1196),
.B2(n_1123),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1140),
.A2(n_1183),
.B1(n_1203),
.B2(n_1141),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1192),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1162),
.A2(n_1201),
.B1(n_1211),
.B2(n_1210),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1136),
.Y(n_1232)
);

CKINVDCx6p67_ASAP7_75t_R g1233 ( 
.A(n_1126),
.Y(n_1233)
);

AOI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1172),
.A2(n_1185),
.B(n_1130),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1112),
.A2(n_1201),
.B(n_1162),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1157),
.Y(n_1236)
);

CKINVDCx11_ASAP7_75t_R g1237 ( 
.A(n_1192),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_1101),
.B(n_1199),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1120),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_1119),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1183),
.A2(n_1203),
.B1(n_1141),
.B2(n_1128),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1110),
.A2(n_1085),
.B1(n_1111),
.B2(n_1210),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1109),
.Y(n_1243)
);

BUFx8_ASAP7_75t_L g1244 ( 
.A(n_1113),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1084),
.A2(n_1171),
.B1(n_1208),
.B2(n_1206),
.Y(n_1245)
);

CKINVDCx11_ASAP7_75t_R g1246 ( 
.A(n_1160),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1211),
.A2(n_1091),
.B1(n_1086),
.B2(n_1129),
.Y(n_1247)
);

INVx5_ASAP7_75t_SL g1248 ( 
.A(n_1144),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1082),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1173),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1084),
.A2(n_1208),
.B1(n_1206),
.B2(n_1171),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1115),
.A2(n_1122),
.B1(n_1168),
.B2(n_1189),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_R g1253 ( 
.A1(n_1089),
.A2(n_1092),
.B1(n_1193),
.B2(n_1180),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1177),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1088),
.A2(n_1109),
.B1(n_1143),
.B2(n_1131),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1198),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1209),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1091),
.A2(n_1100),
.B1(n_1125),
.B2(n_1090),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1106),
.A2(n_1185),
.B1(n_1172),
.B2(n_1134),
.Y(n_1259)
);

CKINVDCx16_ASAP7_75t_R g1260 ( 
.A(n_1207),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1131),
.A2(n_1148),
.B1(n_1081),
.B2(n_1146),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1159),
.B(n_1178),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1165),
.A2(n_1137),
.B1(n_1134),
.B2(n_1209),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1081),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1131),
.A2(n_1148),
.B1(n_1082),
.B2(n_1144),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1174),
.A2(n_1147),
.B1(n_1152),
.B2(n_1131),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1100),
.A2(n_1082),
.B1(n_1153),
.B2(n_1133),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1082),
.A2(n_1144),
.B1(n_1153),
.B2(n_1135),
.Y(n_1268)
);

BUFx5_ASAP7_75t_L g1269 ( 
.A(n_1093),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1104),
.A2(n_1133),
.B1(n_1181),
.B2(n_1145),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1145),
.Y(n_1271)
);

CKINVDCx6p67_ASAP7_75t_R g1272 ( 
.A(n_1194),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1150),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1124),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1156),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1145),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1194),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1181),
.A2(n_1132),
.B1(n_1139),
.B2(n_1097),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1156),
.A2(n_1118),
.B1(n_1102),
.B2(n_1095),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1142),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1149),
.A2(n_1102),
.B1(n_1151),
.B2(n_1114),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1149),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1107),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1116),
.A2(n_1151),
.B1(n_1169),
.B2(n_1083),
.Y(n_1284)
);

BUFx4_ASAP7_75t_R g1285 ( 
.A(n_1158),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1164),
.A2(n_1182),
.B1(n_1200),
.B2(n_1186),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1158),
.Y(n_1287)
);

INVxp67_ASAP7_75t_SL g1288 ( 
.A(n_1175),
.Y(n_1288)
);

INVx8_ASAP7_75t_L g1289 ( 
.A(n_1158),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1184),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1205),
.A2(n_731),
.B1(n_1204),
.B2(n_877),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1167),
.A2(n_774),
.B1(n_1063),
.B2(n_962),
.Y(n_1292)
);

BUFx2_ASAP7_75t_R g1293 ( 
.A(n_1167),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1113),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1170),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1204),
.A2(n_962),
.B(n_1094),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_1155),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1124),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1161),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1187),
.A2(n_1070),
.B1(n_962),
.B2(n_1108),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1108),
.A2(n_962),
.B1(n_731),
.B2(n_1204),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1127),
.Y(n_1308)
);

BUFx8_ASAP7_75t_L g1309 ( 
.A(n_1113),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1204),
.A2(n_774),
.B1(n_1063),
.B2(n_962),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1204),
.A2(n_962),
.B(n_1094),
.Y(n_1311)
);

CKINVDCx8_ASAP7_75t_R g1312 ( 
.A(n_1113),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1082),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1166),
.Y(n_1314)
);

BUFx8_ASAP7_75t_L g1315 ( 
.A(n_1113),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1166),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1251),
.B(n_1245),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1273),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1275),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1287),
.B(n_1278),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1235),
.A2(n_1231),
.B(n_1223),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1307),
.A2(n_1291),
.B1(n_1306),
.B2(n_1304),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1251),
.B(n_1305),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1282),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1235),
.A2(n_1231),
.B(n_1223),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1289),
.B(n_1249),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1310),
.A2(n_1212),
.B(n_1218),
.Y(n_1327)
);

BUFx2_ASAP7_75t_SL g1328 ( 
.A(n_1269),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1214),
.B(n_1258),
.Y(n_1329)
);

BUFx2_ASAP7_75t_R g1330 ( 
.A(n_1312),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1280),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1269),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1275),
.Y(n_1333)
);

AOI221xp5_ASAP7_75t_L g1334 ( 
.A1(n_1298),
.A2(n_1311),
.B1(n_1310),
.B2(n_1292),
.C(n_1307),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1226),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1226),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1214),
.B(n_1258),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1225),
.B(n_1224),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1305),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1289),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1274),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1274),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1302),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1220),
.B(n_1217),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1302),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1281),
.A2(n_1238),
.B(n_1283),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1308),
.Y(n_1347)
);

INVx4_ASAP7_75t_SL g1348 ( 
.A(n_1249),
.Y(n_1348)
);

AO21x1_ASAP7_75t_L g1349 ( 
.A1(n_1218),
.A2(n_1234),
.B(n_1263),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_SL g1350 ( 
.A(n_1244),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1222),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1236),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1290),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1285),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1238),
.A2(n_1288),
.B(n_1262),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1269),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1242),
.B(n_1228),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1291),
.A2(n_1297),
.B1(n_1296),
.B2(n_1299),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1242),
.B(n_1228),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1250),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1234),
.A2(n_1262),
.B(n_1259),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1254),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1293),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1269),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1239),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1267),
.A2(n_1247),
.B(n_1288),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1269),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1247),
.B(n_1293),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1270),
.A2(n_1229),
.B(n_1241),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1268),
.A2(n_1265),
.B(n_1255),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1269),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1221),
.B(n_1219),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1279),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1261),
.B(n_1266),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1295),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1279),
.B(n_1264),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1267),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1276),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1271),
.A2(n_1257),
.B(n_1215),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1253),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1284),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1301),
.A2(n_1219),
.B1(n_1243),
.B2(n_1252),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1276),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1284),
.A2(n_1286),
.B(n_1313),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1347),
.B(n_1260),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1377),
.B(n_1318),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1377),
.B(n_1232),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1323),
.B(n_1339),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1339),
.B(n_1335),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1349),
.A2(n_1374),
.B(n_1327),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1357),
.B(n_1230),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1367),
.A2(n_1216),
.B(n_1303),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1369),
.B(n_1240),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1336),
.B(n_1272),
.Y(n_1397)
);

NAND4xp25_ASAP7_75t_SL g1398 ( 
.A(n_1334),
.B(n_1315),
.C(n_1294),
.D(n_1309),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1329),
.A2(n_1213),
.B(n_1277),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1360),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1340),
.B(n_1233),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1381),
.A2(n_1256),
.B1(n_1315),
.B2(n_1244),
.Y(n_1402)
);

NAND4xp25_ASAP7_75t_L g1403 ( 
.A(n_1381),
.B(n_1237),
.C(n_1294),
.D(n_1309),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1360),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1364),
.B(n_1246),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1336),
.B(n_1227),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1364),
.B(n_1227),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1357),
.A2(n_1300),
.B1(n_1359),
.B2(n_1337),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1355),
.A2(n_1382),
.B(n_1346),
.Y(n_1409)
);

AOI211xp5_ASAP7_75t_L g1410 ( 
.A1(n_1337),
.A2(n_1300),
.B(n_1359),
.C(n_1349),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1317),
.A2(n_1361),
.B(n_1373),
.C(n_1374),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1373),
.A2(n_1382),
.B(n_1386),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1321),
.A2(n_1325),
.B(n_1378),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1322),
.A2(n_1358),
.B1(n_1375),
.B2(n_1383),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1366),
.B(n_1324),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_L g1416 ( 
.A(n_1332),
.B(n_1341),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_R g1417 ( 
.A(n_1331),
.B(n_1350),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1386),
.A2(n_1380),
.B(n_1338),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1354),
.C(n_1320),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1375),
.A2(n_1344),
.B1(n_1331),
.B2(n_1352),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1380),
.A2(n_1341),
.B(n_1342),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1354),
.A2(n_1363),
.B1(n_1330),
.B2(n_1368),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1342),
.A2(n_1343),
.B(n_1345),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1376),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1362),
.Y(n_1425)
);

AO32x2_ASAP7_75t_L g1426 ( 
.A1(n_1332),
.A2(n_1379),
.A3(n_1384),
.B1(n_1344),
.B2(n_1362),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_L g1428 ( 
.A(n_1379),
.B(n_1384),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1326),
.B(n_1348),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1372),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1348),
.B(n_1387),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1343),
.B(n_1345),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1400),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1385),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1404),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1425),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1409),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1410),
.A2(n_1372),
.B1(n_1365),
.B2(n_1328),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1391),
.B(n_1333),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1426),
.B(n_1319),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1392),
.B(n_1333),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1432),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1426),
.B(n_1385),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1426),
.B(n_1385),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1427),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1389),
.B(n_1355),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1421),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1414),
.A2(n_1363),
.B1(n_1320),
.B2(n_1370),
.Y(n_1448)
);

NOR2x1_ASAP7_75t_L g1449 ( 
.A(n_1416),
.B(n_1332),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1423),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1393),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1393),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1430),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1429),
.B(n_1356),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1418),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1437),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1439),
.B(n_1388),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.B(n_1446),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1438),
.A2(n_1410),
.B1(n_1414),
.B2(n_1408),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1433),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1415),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1390),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1448),
.A2(n_1412),
.B1(n_1420),
.B2(n_1422),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1438),
.A2(n_1420),
.B1(n_1411),
.B2(n_1422),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1443),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1443),
.A2(n_1394),
.B(n_1419),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1406),
.Y(n_1467)
);

OAI211xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1453),
.A2(n_1397),
.B(n_1399),
.C(n_1405),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1446),
.B(n_1396),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1446),
.B(n_1353),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1433),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1431),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1433),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1435),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1435),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1441),
.B(n_1407),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1436),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1447),
.B(n_1412),
.Y(n_1478)
);

NAND2x1_ASAP7_75t_L g1479 ( 
.A(n_1449),
.B(n_1401),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1447),
.B(n_1395),
.C(n_1428),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1465),
.B(n_1454),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1460),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1469),
.B(n_1445),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1460),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1458),
.B(n_1444),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1471),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1458),
.B(n_1444),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1478),
.B(n_1447),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1469),
.B(n_1453),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1473),
.B(n_1450),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1472),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1473),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1474),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1474),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1475),
.B(n_1450),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1445),
.Y(n_1502)
);

INVx3_ASAP7_75t_SL g1503 ( 
.A(n_1472),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1465),
.B(n_1434),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1456),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1456),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1476),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_L g1509 ( 
.A(n_1479),
.B(n_1403),
.Y(n_1509)
);

OAI211xp5_ASAP7_75t_L g1510 ( 
.A1(n_1480),
.A2(n_1434),
.B(n_1403),
.C(n_1455),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1465),
.B(n_1434),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1465),
.B(n_1434),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1467),
.B(n_1442),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1482),
.Y(n_1514)
);

AOI21xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1510),
.A2(n_1503),
.B(n_1464),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1482),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1485),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1465),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1508),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1509),
.B(n_1417),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1485),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1488),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1499),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1488),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1484),
.B(n_1455),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1490),
.B(n_1455),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1510),
.A2(n_1465),
.B1(n_1464),
.B2(n_1459),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1499),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1499),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1424),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1513),
.B(n_1457),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1487),
.B(n_1465),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1503),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1496),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1487),
.B(n_1472),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1506),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1491),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1487),
.B(n_1461),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1505),
.B(n_1476),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_1467),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1503),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1491),
.B(n_1467),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1497),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1498),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1498),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1514),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1518),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1502),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1532),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1543),
.B(n_1494),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1481),
.Y(n_1561)
);

NAND2x1_ASAP7_75t_L g1562 ( 
.A(n_1547),
.B(n_1481),
.Y(n_1562)
);

NOR2xp67_ASAP7_75t_SL g1563 ( 
.A(n_1547),
.B(n_1480),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1538),
.B(n_1481),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1543),
.B(n_1495),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1528),
.B(n_1547),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1535),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1417),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1514),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1516),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1550),
.Y(n_1571)
);

INVx3_ASAP7_75t_SL g1572 ( 
.A(n_1535),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1516),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1550),
.B(n_1495),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1517),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1515),
.B(n_1459),
.C(n_1463),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1526),
.A2(n_1463),
.B1(n_1466),
.B2(n_1448),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1521),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1523),
.B(n_1519),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1521),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1524),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.B(n_1495),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1524),
.B(n_1402),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1502),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1548),
.B(n_1505),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1527),
.A2(n_1466),
.B1(n_1452),
.B2(n_1451),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1533),
.B(n_1493),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1563),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1577),
.B(n_1559),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1552),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1578),
.A2(n_1504),
.B(n_1512),
.C(n_1511),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1566),
.A2(n_1540),
.B(n_1533),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1568),
.B(n_1398),
.Y(n_1595)
);

NOR4xp75_ASAP7_75t_L g1596 ( 
.A(n_1566),
.B(n_1479),
.C(n_1504),
.D(n_1511),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1544),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1572),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1544),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_SL g1603 ( 
.A(n_1580),
.B(n_1402),
.C(n_1468),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1534),
.Y(n_1604)
);

CKINVDCx16_ASAP7_75t_R g1605 ( 
.A(n_1584),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1556),
.B(n_1553),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1587),
.A2(n_1534),
.B1(n_1504),
.B2(n_1511),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1555),
.B(n_1534),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1584),
.A2(n_1512),
.B1(n_1489),
.B2(n_1486),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1584),
.A2(n_1500),
.B(n_1493),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1584),
.A2(n_1501),
.B(n_1500),
.Y(n_1611)
);

O2A1O1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1572),
.A2(n_1512),
.B(n_1468),
.C(n_1525),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1569),
.Y(n_1613)
);

OAI321xp33_ASAP7_75t_L g1614 ( 
.A1(n_1590),
.A2(n_1555),
.A3(n_1557),
.B1(n_1567),
.B2(n_1588),
.C(n_1582),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1591),
.B(n_1572),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1591),
.B(n_1604),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1590),
.B(n_1558),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1597),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1598),
.B(n_1586),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1599),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1605),
.A2(n_1609),
.B1(n_1611),
.B2(n_1610),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1612),
.A2(n_1594),
.B(n_1600),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1613),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1593),
.B(n_1585),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1606),
.B(n_1573),
.Y(n_1627)
);

OAI211xp5_ASAP7_75t_L g1628 ( 
.A1(n_1603),
.A2(n_1562),
.B(n_1574),
.C(n_1581),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1558),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1607),
.A2(n_1558),
.B1(n_1486),
.B2(n_1489),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1593),
.B(n_1601),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1615),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1621),
.B(n_1616),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1616),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1632),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1627),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1622),
.A2(n_1582),
.B1(n_1451),
.B2(n_1452),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1621),
.B(n_1602),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1592),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1628),
.B(n_1596),
.C(n_1595),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1486),
.C(n_1489),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1615),
.B(n_1561),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1635),
.B(n_1629),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1634),
.B(n_1623),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1636),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_SL g1647 ( 
.A1(n_1641),
.A2(n_1617),
.B(n_1619),
.C(n_1624),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1633),
.B(n_1617),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1643),
.B(n_1626),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1637),
.B(n_1631),
.C(n_1620),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1639),
.B(n_1627),
.Y(n_1651)
);

NAND5xp2_ASAP7_75t_L g1652 ( 
.A(n_1640),
.B(n_1630),
.C(n_1625),
.D(n_1618),
.E(n_1565),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1642),
.B(n_1561),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1647),
.A2(n_1641),
.B(n_1574),
.C(n_1570),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1645),
.A2(n_1581),
.B(n_1579),
.C(n_1569),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1651),
.A2(n_1564),
.B1(n_1561),
.B2(n_1562),
.Y(n_1657)
);

AOI31xp33_ASAP7_75t_L g1658 ( 
.A1(n_1648),
.A2(n_1564),
.A3(n_1579),
.B(n_1570),
.Y(n_1658)
);

O2A1O1Ixp5_ASAP7_75t_L g1659 ( 
.A1(n_1654),
.A2(n_1649),
.B(n_1650),
.C(n_1653),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1657),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1646),
.B1(n_1576),
.B2(n_1564),
.Y(n_1661)
);

OAI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1655),
.A2(n_1646),
.B(n_1652),
.C(n_1638),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_L g1663 ( 
.A(n_1656),
.B(n_1539),
.C(n_1529),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1654),
.A2(n_1530),
.B1(n_1522),
.B2(n_1536),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1661),
.B(n_1565),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1659),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1660),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1662),
.B(n_1522),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1664),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1666),
.A2(n_1663),
.B1(n_1541),
.B2(n_1531),
.Y(n_1670)
);

AND3x1_ASAP7_75t_L g1671 ( 
.A(n_1668),
.B(n_1583),
.C(n_1575),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1667),
.A2(n_1542),
.B1(n_1530),
.B2(n_1551),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1671),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1673),
.Y(n_1674)
);

XNOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1674),
.B(n_1669),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1674),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1676),
.B(n_1670),
.C(n_1672),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1675),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1677),
.A2(n_1665),
.B1(n_1525),
.B2(n_1551),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1541),
.B(n_1537),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1545),
.B1(n_1537),
.B2(n_1539),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1681),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1679),
.B1(n_1529),
.B2(n_1531),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1542),
.B1(n_1536),
.B2(n_1549),
.C(n_1545),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1583),
.B(n_1575),
.C(n_1401),
.Y(n_1685)
);


endmodule