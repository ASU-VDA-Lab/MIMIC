module fake_jpeg_30155_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_14),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_35),
.B(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_51),
.Y(n_79)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_8),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_77),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_22),
.B1(n_28),
.B2(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_36),
.A2(n_29),
.B1(n_33),
.B2(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_28),
.B1(n_32),
.B2(n_29),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_48),
.B1(n_28),
.B2(n_47),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_21),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_55),
.Y(n_103)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_19),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_24),
.B(n_30),
.C(n_21),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_49),
.B1(n_37),
.B2(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_109),
.B1(n_86),
.B2(n_81),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_102),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_27),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_110),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_83),
.C(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_116),
.C(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_2),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_61),
.B(n_58),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_74),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_130),
.C(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_99),
.B1(n_113),
.B2(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_114),
.B(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_68),
.B1(n_86),
.B2(n_87),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_125),
.B1(n_93),
.B2(n_62),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_98),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_58),
.C(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_105),
.B1(n_95),
.B2(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_152),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_100),
.B(n_97),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_26),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_69),
.B1(n_26),
.B2(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_59),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_122),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_2),
.B(n_3),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_4),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_118),
.A3(n_125),
.B1(n_134),
.B2(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_136),
.Y(n_164)
);

NAND2xp67_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_137),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_169),
.C(n_132),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_151),
.C(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_177),
.C(n_5),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_143),
.B(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_151),
.C(n_141),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_160),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_178),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_147),
.C(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_149),
.B1(n_139),
.B2(n_140),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_168),
.B1(n_165),
.B2(n_159),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_155),
.C(n_148),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_158),
.A3(n_132),
.B1(n_153),
.B2(n_122),
.C1(n_119),
.C2(n_8),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_186),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_185),
.B1(n_170),
.B2(n_180),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_163),
.B1(n_158),
.B2(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_181),
.C(n_186),
.Y(n_196)
);

OAI221xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_187),
.B1(n_173),
.B2(n_193),
.C(n_182),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_190),
.B(n_171),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_193),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_174),
.B(n_196),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_195),
.B(n_5),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_6),
.B(n_202),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_6),
.Y(n_205)
);


endmodule