module real_aes_16839_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g462 ( .A(n_0), .Y(n_462) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1), .Y(n_1088) );
AOI221x1_ASAP7_75t_SL g1104 ( .A1(n_1), .A2(n_2), .B1(n_547), .B2(n_716), .C(n_1105), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_2), .A2(n_23), .B1(n_323), .B2(n_1092), .Y(n_1096) );
AOI221x1_ASAP7_75t_SL g477 ( .A1(n_3), .A2(n_240), .B1(n_478), .B2(n_482), .C(n_483), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_3), .A2(n_568), .B(n_569), .Y(n_567) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_4), .B(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_5), .Y(n_734) );
INVx1_ASAP7_75t_L g914 ( .A(n_6), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_7), .A2(n_96), .B1(n_307), .B2(n_310), .C(n_315), .Y(n_306) );
INVx1_ASAP7_75t_L g388 ( .A(n_7), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g1019 ( .A1(n_8), .A2(n_205), .B1(n_1020), .B2(n_1023), .C(n_1024), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_8), .A2(n_205), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_9), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_9), .A2(n_28), .B1(n_318), .B2(n_355), .Y(n_992) );
INVx1_ASAP7_75t_L g1018 ( .A(n_10), .Y(n_1018) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_10), .A2(n_241), .B1(n_1037), .B2(n_1039), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_11), .A2(n_235), .B1(n_315), .B2(n_956), .C(n_1013), .Y(n_1012) );
AOI222xp33_ASAP7_75t_L g1049 ( .A1(n_11), .A2(n_62), .B1(n_135), .B2(n_373), .C1(n_731), .C2(n_929), .Y(n_1049) );
AOI21xp33_ASAP7_75t_L g1095 ( .A1(n_12), .A2(n_657), .B(n_658), .Y(n_1095) );
INVx1_ASAP7_75t_L g1114 ( .A(n_12), .Y(n_1114) );
INVx1_ASAP7_75t_L g263 ( .A(n_13), .Y(n_263) );
AND2x2_ASAP7_75t_L g288 ( .A(n_13), .B(n_215), .Y(n_288) );
AND2x2_ASAP7_75t_L g328 ( .A(n_13), .B(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_13), .B(n_273), .Y(n_497) );
INVx1_ASAP7_75t_L g1125 ( .A(n_14), .Y(n_1125) );
OAI211xp5_ASAP7_75t_L g1162 ( .A1(n_14), .A2(n_782), .B(n_821), .C(n_1163), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_15), .A2(n_170), .B1(n_592), .B2(n_728), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_15), .A2(n_81), .B1(n_340), .B2(n_341), .C(n_756), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g875 ( .A1(n_16), .A2(n_876), .B(n_877), .C(n_883), .Y(n_875) );
INVx1_ASAP7_75t_L g893 ( .A(n_16), .Y(n_893) );
INVx1_ASAP7_75t_L g1455 ( .A(n_17), .Y(n_1455) );
INVx1_ASAP7_75t_L g825 ( .A(n_18), .Y(n_825) );
INVx1_ASAP7_75t_L g778 ( .A(n_19), .Y(n_778) );
INVx1_ASAP7_75t_L g721 ( .A(n_20), .Y(n_721) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_21), .B(n_1182), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_21), .B(n_92), .Y(n_1184) );
INVx2_ASAP7_75t_L g1188 ( .A(n_21), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_22), .A2(n_151), .B1(n_867), .B2(n_869), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_22), .A2(n_151), .B1(n_702), .B2(n_895), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_23), .A2(n_174), .B1(n_547), .B2(n_1110), .C(n_1112), .Y(n_1109) );
INVx1_ASAP7_75t_L g1428 ( .A(n_24), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_25), .A2(n_129), .B1(n_284), .B2(n_518), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_25), .A2(n_219), .B1(n_530), .B2(n_532), .C(n_534), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_26), .A2(n_165), .B1(n_1183), .B2(n_1189), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_27), .A2(n_41), .B1(n_265), .B2(n_874), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_27), .A2(n_41), .B1(n_886), .B2(n_888), .Y(n_885) );
INVxp67_ASAP7_75t_SL g973 ( .A(n_28), .Y(n_973) );
OAI211xp5_ASAP7_75t_L g817 ( .A1(n_29), .A2(n_818), .B(n_821), .C(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g852 ( .A(n_29), .Y(n_852) );
INVx1_ASAP7_75t_L g1432 ( .A(n_30), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_31), .A2(n_200), .B1(n_718), .B2(n_719), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_31), .A2(n_57), .B1(n_667), .B2(n_740), .C(n_742), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_32), .A2(n_69), .B1(n_318), .B2(n_323), .Y(n_317) );
INVx1_ASAP7_75t_L g397 ( .A(n_32), .Y(n_397) );
INVx1_ASAP7_75t_L g957 ( .A(n_33), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_34), .A2(n_199), .B1(n_1179), .B2(n_1186), .Y(n_1236) );
INVx1_ASAP7_75t_L g1145 ( .A(n_35), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_36), .A2(n_243), .B1(n_867), .B2(n_869), .Y(n_1403) );
OAI22xp33_ASAP7_75t_L g1411 ( .A1(n_36), .A2(n_243), .B1(n_895), .B2(n_1166), .Y(n_1411) );
INVx1_ASAP7_75t_L g643 ( .A(n_37), .Y(n_643) );
INVx1_ASAP7_75t_L g913 ( .A(n_38), .Y(n_913) );
INVx1_ASAP7_75t_L g1124 ( .A(n_39), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_40), .A2(n_214), .B1(n_338), .B2(n_341), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_40), .A2(n_96), .B1(n_399), .B2(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g1427 ( .A(n_42), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_43), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_44), .A2(n_72), .B1(n_550), .B2(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g633 ( .A(n_44), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_45), .A2(n_154), .B1(n_874), .B2(n_962), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_45), .A2(n_154), .B1(n_1159), .B2(n_1161), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g1208 ( .A1(n_46), .A2(n_208), .B1(n_1179), .B2(n_1189), .Y(n_1208) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_47), .A2(n_101), .B1(n_1179), .B2(n_1186), .Y(n_1218) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_48), .A2(n_89), .B1(n_1179), .B2(n_1186), .Y(n_1220) );
INVx1_ASAP7_75t_L g975 ( .A(n_49), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_49), .A2(n_121), .B1(n_338), .B2(n_988), .Y(n_987) );
OAI22xp5_ASAP7_75t_SL g1078 ( .A1(n_50), .A2(n_172), .B1(n_292), .B2(n_424), .Y(n_1078) );
INVx1_ASAP7_75t_L g1082 ( .A(n_50), .Y(n_1082) );
INVx1_ASAP7_75t_L g909 ( .A(n_51), .Y(n_909) );
INVx1_ASAP7_75t_L g296 ( .A(n_52), .Y(n_296) );
INVx1_ASAP7_75t_L g369 ( .A(n_52), .Y(n_369) );
INVxp67_ASAP7_75t_SL g1028 ( .A(n_53), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_53), .A2(n_235), .B1(n_537), .B2(n_588), .Y(n_1057) );
INVx1_ASAP7_75t_L g827 ( .A(n_54), .Y(n_827) );
OAI211xp5_ASAP7_75t_L g839 ( .A1(n_54), .A2(n_840), .B(n_843), .C(n_846), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_55), .Y(n_492) );
INVx1_ASAP7_75t_L g356 ( .A(n_56), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_57), .A2(n_177), .B1(n_588), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g256 ( .A(n_58), .Y(n_256) );
INVx2_ASAP7_75t_L g302 ( .A(n_59), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_60), .A2(n_76), .B1(n_1186), .B2(n_1193), .Y(n_1209) );
OAI22xp33_ASAP7_75t_L g1457 ( .A1(n_61), .A2(n_138), .B1(n_895), .B2(n_1458), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_61), .A2(n_138), .B1(n_1128), .B2(n_1466), .Y(n_1465) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_62), .A2(n_146), .B1(n_338), .B2(n_1015), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_63), .A2(n_145), .B1(n_874), .B2(n_962), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_63), .A2(n_145), .B1(n_815), .B2(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g955 ( .A(n_64), .Y(n_955) );
INVx1_ASAP7_75t_L g920 ( .A(n_65), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_66), .A2(n_93), .B1(n_307), .B2(n_334), .C(n_335), .Y(n_333) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_66), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g1451 ( .A1(n_67), .A2(n_117), .B1(n_1003), .B2(n_1407), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_67), .A2(n_117), .B1(n_874), .B2(n_1461), .Y(n_1460) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_68), .A2(n_115), .B1(n_1179), .B2(n_1186), .Y(n_1202) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_69), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g1121 ( .A1(n_70), .A2(n_986), .B(n_1122), .C(n_1123), .Y(n_1121) );
INVx1_ASAP7_75t_L g1164 ( .A(n_70), .Y(n_1164) );
XOR2xp5_ASAP7_75t_L g1421 ( .A(n_71), .B(n_1422), .Y(n_1421) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_72), .A2(n_110), .B1(n_341), .B2(n_609), .C(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g882 ( .A(n_73), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g889 ( .A1(n_73), .A2(n_821), .B(n_890), .C(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g725 ( .A(n_74), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_75), .A2(n_163), .B1(n_485), .B2(n_487), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_75), .B(n_702), .Y(n_701) );
XOR2x2_ASAP7_75t_L g862 ( .A(n_76), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g1059 ( .A(n_77), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_78), .Y(n_1383) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_79), .Y(n_604) );
INVx1_ASAP7_75t_L g1094 ( .A(n_80), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_81), .A2(n_111), .B1(n_594), .B2(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_82), .A2(n_116), .B1(n_1179), .B2(n_1186), .Y(n_1206) );
OA222x2_ASAP7_75t_L g464 ( .A1(n_83), .A2(n_201), .B1(n_219), .B2(n_465), .C1(n_467), .C2(n_473), .Y(n_464) );
INVx1_ASAP7_75t_L g546 ( .A(n_83), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_84), .A2(n_1118), .B1(n_1119), .B2(n_1167), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_84), .Y(n_1167) );
AOI22xp5_ASAP7_75t_SL g1205 ( .A1(n_84), .A2(n_242), .B1(n_1189), .B2(n_1193), .Y(n_1205) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_85), .Y(n_258) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_85), .B(n_256), .Y(n_1180) );
OAI211xp5_ASAP7_75t_SL g1009 ( .A1(n_86), .A2(n_1010), .B(n_1011), .C(n_1016), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_86), .A2(n_206), .B1(n_447), .B2(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g1007 ( .A(n_88), .B(n_1008), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_90), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g1217 ( .A1(n_91), .A2(n_102), .B1(n_1183), .B2(n_1189), .Y(n_1217) );
INVx1_ASAP7_75t_L g1182 ( .A(n_92), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_92), .B(n_1188), .Y(n_1190) );
INVx1_ASAP7_75t_L g395 ( .A(n_93), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_94), .A2(n_184), .B1(n_340), .B2(n_355), .Y(n_659) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_94), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_95), .A2(n_100), .B1(n_547), .B2(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g636 ( .A(n_95), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_97), .Y(n_1027) );
INVx1_ASAP7_75t_L g581 ( .A(n_98), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_98), .A2(n_223), .B1(n_486), .B2(n_490), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_99), .A2(n_245), .B1(n_1179), .B2(n_1183), .Y(n_1178) );
INVx1_ASAP7_75t_L g614 ( .A(n_100), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g1390 ( .A(n_103), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_104), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g380 ( .A(n_104), .Y(n_380) );
INVx1_ASAP7_75t_L g414 ( .A(n_104), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_105), .A2(n_226), .B1(n_1179), .B2(n_1186), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1404 ( .A1(n_106), .A2(n_168), .B1(n_874), .B2(n_962), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g1406 ( .A1(n_106), .A2(n_168), .B1(n_1003), .B2(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1133 ( .A(n_107), .Y(n_1133) );
INVx1_ASAP7_75t_L g781 ( .A(n_108), .Y(n_781) );
INVx1_ASAP7_75t_L g1434 ( .A(n_109), .Y(n_1434) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_110), .A2(n_148), .B1(n_588), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g744 ( .A(n_111), .Y(n_744) );
INVx1_ASAP7_75t_L g958 ( .A(n_112), .Y(n_958) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_113), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_113), .A2(n_220), .B1(n_486), .B2(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_114), .A2(n_239), .B1(n_471), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_114), .A2(n_222), .B1(n_548), .B2(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_118), .B(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_118), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_119), .Y(n_1384) );
OAI211xp5_ASAP7_75t_SL g1399 ( .A1(n_120), .A2(n_804), .B(n_1122), .C(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1410 ( .A(n_120), .Y(n_1410) );
INVxp67_ASAP7_75t_SL g967 ( .A(n_121), .Y(n_967) );
INVx1_ASAP7_75t_L g1456 ( .A(n_122), .Y(n_1456) );
OAI211xp5_ASAP7_75t_L g1462 ( .A1(n_122), .A2(n_883), .B(n_986), .C(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g770 ( .A(n_123), .Y(n_770) );
INVx1_ASAP7_75t_L g1141 ( .A(n_124), .Y(n_1141) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_125), .Y(n_1387) );
INVx1_ASAP7_75t_L g666 ( .A(n_126), .Y(n_666) );
INVx1_ASAP7_75t_L g1064 ( .A(n_127), .Y(n_1064) );
INVx1_ASAP7_75t_L g789 ( .A(n_128), .Y(n_789) );
INVx1_ASAP7_75t_L g549 ( .A(n_129), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g828 ( .A1(n_130), .A2(n_147), .B1(n_829), .B2(n_830), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_130), .A2(n_147), .B1(n_854), .B2(n_856), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_131), .Y(n_506) );
INVx1_ASAP7_75t_L g344 ( .A(n_132), .Y(n_344) );
INVx1_ASAP7_75t_L g735 ( .A(n_133), .Y(n_735) );
INVx1_ASAP7_75t_L g919 ( .A(n_134), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_135), .A2(n_211), .B1(n_334), .B2(n_335), .C(n_1030), .Y(n_1029) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_136), .A2(n_232), .B1(n_1189), .B2(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1437 ( .A(n_137), .Y(n_1437) );
INVx1_ASAP7_75t_L g353 ( .A(n_139), .Y(n_353) );
OAI322xp33_ASAP7_75t_L g361 ( .A1(n_139), .A2(n_362), .A3(n_376), .B1(n_381), .B2(n_391), .C1(n_408), .C2(n_415), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_140), .Y(n_1389) );
BUFx3_ASAP7_75t_L g298 ( .A(n_141), .Y(n_298) );
INVx1_ASAP7_75t_L g1144 ( .A(n_142), .Y(n_1144) );
INVx1_ASAP7_75t_L g303 ( .A(n_143), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_144), .A2(n_247), .B1(n_340), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_144), .A2(n_186), .B1(n_404), .B2(n_536), .Y(n_678) );
INVx1_ASAP7_75t_L g1056 ( .A(n_146), .Y(n_1056) );
AOI211xp5_ASAP7_75t_SL g630 ( .A1(n_148), .A2(n_631), .B(n_632), .C(n_635), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_149), .Y(n_723) );
INVx1_ASAP7_75t_L g759 ( .A(n_150), .Y(n_759) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_152), .Y(n_270) );
INVx1_ASAP7_75t_L g968 ( .A(n_153), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_155), .A2(n_188), .B1(n_592), .B2(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g613 ( .A(n_155), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_156), .A2(n_190), .B1(n_669), .B2(n_671), .C(n_672), .Y(n_668) );
INVx1_ASAP7_75t_L g689 ( .A(n_156), .Y(n_689) );
OAI22xp33_ASAP7_75t_SL g653 ( .A1(n_157), .A2(n_204), .B1(n_504), .B2(n_634), .Y(n_653) );
INVx1_ASAP7_75t_L g692 ( .A(n_157), .Y(n_692) );
AOI21xp5_ASAP7_75t_SL g662 ( .A1(n_158), .A2(n_335), .B(n_657), .Y(n_662) );
INVx1_ASAP7_75t_L g676 ( .A(n_158), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g1401 ( .A(n_159), .Y(n_1401) );
INVx1_ASAP7_75t_L g655 ( .A(n_160), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_160), .A2(n_247), .B1(n_536), .B2(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g791 ( .A(n_161), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_162), .Y(n_661) );
INVx1_ASAP7_75t_L g691 ( .A(n_163), .Y(n_691) );
INVx1_ASAP7_75t_L g785 ( .A(n_164), .Y(n_785) );
INVx1_ASAP7_75t_L g980 ( .A(n_166), .Y(n_980) );
INVx1_ASAP7_75t_L g902 ( .A(n_167), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_169), .Y(n_421) );
INVx1_ASAP7_75t_L g743 ( .A(n_170), .Y(n_743) );
INVx1_ASAP7_75t_L g949 ( .A(n_171), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g1086 ( .A(n_172), .Y(n_1086) );
INVx1_ASAP7_75t_L g951 ( .A(n_173), .Y(n_951) );
AOI21xp33_ASAP7_75t_L g1089 ( .A1(n_174), .A2(n_334), .B(n_1090), .Y(n_1089) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_175), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_176), .Y(n_579) );
INVx1_ASAP7_75t_L g757 ( .A(n_177), .Y(n_757) );
INVx1_ASAP7_75t_L g880 ( .A(n_178), .Y(n_880) );
INVx1_ASAP7_75t_L g330 ( .A(n_179), .Y(n_330) );
OAI222xp33_ASAP7_75t_L g1066 ( .A1(n_180), .A2(n_217), .B1(n_229), .B2(n_447), .C1(n_1067), .C2(n_1070), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_181), .A2(n_248), .B1(n_1189), .B2(n_1193), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_182), .A2(n_189), .B1(n_1183), .B2(n_1189), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_183), .A2(n_246), .B1(n_323), .B2(n_1092), .Y(n_1091) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_183), .Y(n_1113) );
INVxp67_ASAP7_75t_L g681 ( .A(n_184), .Y(n_681) );
INVx1_ASAP7_75t_L g1430 ( .A(n_185), .Y(n_1430) );
AOI21xp33_ASAP7_75t_L g656 ( .A1(n_186), .A2(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g1402 ( .A(n_187), .Y(n_1402) );
OAI211xp5_ASAP7_75t_L g1408 ( .A1(n_187), .A2(n_782), .B(n_821), .C(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g639 ( .A(n_188), .Y(n_639) );
XOR2x2_ASAP7_75t_L g1374 ( .A(n_189), .B(n_1375), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_189), .A2(n_1418), .B1(n_1420), .B2(n_1467), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_190), .Y(n_695) );
INVx1_ASAP7_75t_L g976 ( .A(n_191), .Y(n_976) );
INVx1_ASAP7_75t_L g905 ( .A(n_192), .Y(n_905) );
INVx1_ASAP7_75t_L g1139 ( .A(n_193), .Y(n_1139) );
INVx1_ASAP7_75t_L g786 ( .A(n_194), .Y(n_786) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_195), .Y(n_269) );
OAI22xp33_ASAP7_75t_L g811 ( .A1(n_196), .A2(n_213), .B1(n_812), .B2(n_815), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_196), .A2(n_213), .B1(n_265), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1135 ( .A(n_197), .Y(n_1135) );
INVx1_ASAP7_75t_L g1148 ( .A(n_198), .Y(n_1148) );
INVx1_ASAP7_75t_L g758 ( .A(n_200), .Y(n_758) );
INVx1_ASAP7_75t_L g535 ( .A(n_201), .Y(n_535) );
INVx1_ASAP7_75t_L g971 ( .A(n_202), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_203), .Y(n_522) );
INVx1_ASAP7_75t_L g698 ( .A(n_204), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g1127 ( .A1(n_207), .A2(n_218), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_207), .A2(n_218), .B1(n_895), .B2(n_1166), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_209), .Y(n_1076) );
INVx1_ASAP7_75t_L g772 ( .A(n_210), .Y(n_772) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_211), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1379 ( .A(n_212), .Y(n_1379) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_214), .Y(n_382) );
BUFx3_ASAP7_75t_L g273 ( .A(n_215), .Y(n_273) );
INVx1_ASAP7_75t_L g329 ( .A(n_215), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_216), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_220), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_221), .Y(n_500) );
INVx1_ASAP7_75t_L g484 ( .A(n_222), .Y(n_484) );
INVx1_ASAP7_75t_L g642 ( .A(n_223), .Y(n_642) );
INVx1_ASAP7_75t_L g911 ( .A(n_224), .Y(n_911) );
INVx1_ASAP7_75t_L g1147 ( .A(n_225), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_227), .Y(n_1386) );
INVx1_ASAP7_75t_L g291 ( .A(n_228), .Y(n_291) );
INVx2_ASAP7_75t_L g360 ( .A(n_228), .Y(n_360) );
INVx1_ASAP7_75t_L g413 ( .A(n_228), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_229), .A2(n_233), .B1(n_1098), .B2(n_1100), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_230), .Y(n_525) );
INVx1_ASAP7_75t_L g1438 ( .A(n_231), .Y(n_1438) );
INVx1_ASAP7_75t_L g646 ( .A(n_232), .Y(n_646) );
INVx1_ASAP7_75t_L g1077 ( .A(n_233), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_234), .A2(n_236), .B1(n_1186), .B2(n_1189), .Y(n_1185) );
INVx1_ASAP7_75t_L g1435 ( .A(n_237), .Y(n_1435) );
OAI211xp5_ASAP7_75t_L g1452 ( .A1(n_238), .A2(n_890), .B(n_1453), .C(n_1454), .Y(n_1452) );
INVx1_ASAP7_75t_L g1464 ( .A(n_238), .Y(n_1464) );
INVx1_ASAP7_75t_L g563 ( .A(n_239), .Y(n_563) );
INVx1_ASAP7_75t_L g562 ( .A(n_240), .Y(n_562) );
INVx1_ASAP7_75t_L g1017 ( .A(n_241), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_244), .Y(n_583) );
INVx1_ASAP7_75t_L g1106 ( .A(n_246), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_274), .B(n_1171), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_259), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_253), .B(n_262), .Y(n_1416) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_255), .B(n_258), .Y(n_1419) );
INVx1_ASAP7_75t_L g1468 ( .A(n_255), .Y(n_1468) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g1470 ( .A(n_258), .B(n_1468), .Y(n_1470) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g860 ( .A(n_262), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g316 ( .A(n_263), .B(n_273), .Y(n_316) );
AND2x4_ASAP7_75t_L g336 ( .A(n_263), .B(n_272), .Y(n_336) );
INVx1_ASAP7_75t_L g962 ( .A(n_264), .Y(n_962) );
AND2x4_ASAP7_75t_SL g1415 ( .A(n_264), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1461 ( .A(n_264), .Y(n_1461) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
BUFx4f_ASAP7_75t_L g794 ( .A(n_266), .Y(n_794) );
OR2x6_ASAP7_75t_L g855 ( .A(n_266), .B(n_838), .Y(n_855) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g486 ( .A(n_267), .Y(n_486) );
BUFx4f_ASAP7_75t_L g638 ( .A(n_267), .Y(n_638) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
AND2x2_ASAP7_75t_L g309 ( .A(n_269), .B(n_270), .Y(n_309) );
AND2x2_ASAP7_75t_L g313 ( .A(n_269), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g321 ( .A(n_269), .Y(n_321) );
INVx2_ASAP7_75t_L g325 ( .A(n_269), .Y(n_325) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_269), .B(n_270), .Y(n_475) );
INVx2_ASAP7_75t_L g314 ( .A(n_270), .Y(n_314) );
INVx1_ASAP7_75t_L g322 ( .A(n_270), .Y(n_322) );
AND2x2_ASAP7_75t_L g324 ( .A(n_270), .B(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_270), .B(n_325), .Y(n_491) );
OR2x2_ASAP7_75t_L g503 ( .A(n_270), .B(n_321), .Y(n_503) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g845 ( .A(n_272), .Y(n_845) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g848 ( .A(n_273), .Y(n_848) );
AND2x4_ASAP7_75t_L g851 ( .A(n_273), .B(n_286), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_762), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_456), .B1(n_457), .B2(n_761), .Y(n_275) );
INVx1_ASAP7_75t_L g761 ( .A(n_276), .Y(n_761) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
XNOR2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_455), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_281), .B(n_420), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_303), .B1(n_304), .B2(n_357), .C(n_361), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_292), .Y(n_283) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_284), .B(n_292), .Y(n_1035) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x6_ASAP7_75t_L g331 ( .A(n_288), .B(n_308), .Y(n_331) );
INVx1_ASAP7_75t_L g350 ( .A(n_288), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_288), .B(n_320), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_288), .B(n_360), .Y(n_516) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_288), .Y(n_629) );
INVxp67_ASAP7_75t_L g449 ( .A(n_289), .Y(n_449) );
INVx1_ASAP7_75t_L g524 ( .A(n_289), .Y(n_524) );
INVx1_ASAP7_75t_L g861 ( .A(n_289), .Y(n_861) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g300 ( .A(n_290), .Y(n_300) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g578 ( .A(n_292), .Y(n_578) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_299), .Y(n_292) );
INVx4_ASAP7_75t_L g557 ( .A(n_293), .Y(n_557) );
INVx3_ASAP7_75t_L g566 ( .A(n_293), .Y(n_566) );
BUFx6f_ASAP7_75t_L g978 ( .A(n_293), .Y(n_978) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g390 ( .A(n_294), .Y(n_390) );
BUFx2_ASAP7_75t_L g820 ( .A(n_294), .Y(n_820) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
BUFx2_ASAP7_75t_L g700 ( .A(n_295), .Y(n_700) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_296), .B(n_298), .Y(n_375) );
INVx2_ASAP7_75t_L g407 ( .A(n_296), .Y(n_407) );
INVx2_ASAP7_75t_L g436 ( .A(n_297), .Y(n_436) );
AND2x4_ASAP7_75t_L g548 ( .A(n_297), .B(n_442), .Y(n_548) );
BUFx2_ASAP7_75t_L g697 ( .A(n_297), .Y(n_697) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g370 ( .A(n_298), .Y(n_370) );
OR2x2_ASAP7_75t_L g386 ( .A(n_298), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g406 ( .A(n_298), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
OR2x2_ASAP7_75t_L g424 ( .A(n_299), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g454 ( .A(n_299), .Y(n_454) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
OR2x2_ASAP7_75t_L g378 ( .A(n_300), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g512 ( .A(n_300), .Y(n_512) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_300), .Y(n_710) );
INVx1_ASAP7_75t_L g553 ( .A(n_301), .Y(n_553) );
NAND2xp33_ASAP7_75t_SL g379 ( .A(n_302), .B(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g411 ( .A(n_302), .Y(n_411) );
BUFx3_ASAP7_75t_L g586 ( .A(n_302), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_332), .C(n_351), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_317), .B1(n_326), .B2(n_330), .C(n_331), .Y(n_305) );
BUFx2_ASAP7_75t_L g482 ( .A(n_307), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_307), .A2(n_600), .B1(n_606), .B2(n_621), .C(n_623), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_307), .A2(n_621), .B1(n_721), .B2(n_735), .C(n_748), .Y(n_747) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_SL g327 ( .A(n_308), .B(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g631 ( .A(n_308), .Y(n_631) );
AND2x2_ASAP7_75t_L g844 ( .A(n_308), .B(n_845), .Y(n_844) );
BUFx3_ASAP7_75t_L g956 ( .A(n_308), .Y(n_956) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_308), .Y(n_1030) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g352 ( .A(n_312), .B(n_328), .Y(n_352) );
AND2x2_ASAP7_75t_L g527 ( .A(n_312), .B(n_328), .Y(n_527) );
INVx2_ASAP7_75t_L g622 ( .A(n_312), .Y(n_622) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_312), .Y(n_657) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g334 ( .A(n_313), .Y(n_334) );
INVx2_ASAP7_75t_L g481 ( .A(n_313), .Y(n_481) );
AND2x4_ASAP7_75t_L g837 ( .A(n_313), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g510 ( .A(n_316), .B(n_511), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_316), .A2(n_633), .B(n_634), .Y(n_632) );
INVx4_ASAP7_75t_L g658 ( .A(n_316), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_316), .A2(n_505), .B1(n_634), .B2(n_757), .C(n_758), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_316), .B(n_511), .Y(n_917) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g508 ( .A(n_319), .Y(n_508) );
INVx1_ASAP7_75t_L g1092 ( .A(n_319), .Y(n_1092) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_320), .Y(n_340) );
AND2x2_ASAP7_75t_L g343 ( .A(n_320), .B(n_328), .Y(n_343) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_321), .Y(n_628) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g341 ( .A(n_324), .Y(n_341) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
INVx2_ASAP7_75t_L g472 ( .A(n_324), .Y(n_472) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g1022 ( .A(n_327), .Y(n_1022) );
AND2x4_ASAP7_75t_L g354 ( .A(n_328), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_328), .B(n_413), .Y(n_470) );
BUFx2_ASAP7_75t_L g619 ( .A(n_328), .Y(n_619) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_328), .B(n_471), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_329), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_330), .A2(n_431), .B1(n_437), .B2(n_438), .C(n_443), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_331), .A2(n_1012), .B(n_1014), .Y(n_1011) );
AOI221xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_337), .B1(n_342), .B2(n_344), .C(n_345), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_336), .A2(n_611), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_336), .A2(n_611), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_742) );
INVx2_ASAP7_75t_L g1090 ( .A(n_336), .Y(n_1090) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g609 ( .A(n_339), .Y(n_609) );
INVx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_340), .A2(n_583), .B(n_625), .C(n_629), .Y(n_624) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_340), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g750 ( .A1(n_340), .A2(n_725), .B(n_751), .C(n_754), .Y(n_750) );
AND2x2_ASAP7_75t_L g950 ( .A(n_340), .B(n_848), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_342), .A2(n_352), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g523 ( .A(n_343), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_344), .B(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_346), .Y(n_1023) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g670 ( .A(n_348), .Y(n_670) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g520 ( .A(n_349), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_349), .A2(n_579), .B1(n_604), .B2(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g753 ( .A(n_349), .Y(n_753) );
AND2x2_ASAP7_75t_L g847 ( .A(n_349), .B(n_848), .Y(n_847) );
AND2x4_ASAP7_75t_L g879 ( .A(n_349), .B(n_848), .Y(n_879) );
INVx1_ASAP7_75t_L g754 ( .A(n_350), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_354), .B2(n_356), .Y(n_351) );
INVx3_ASAP7_75t_L g1010 ( .A(n_354), .Y(n_1010) );
INVx1_ASAP7_75t_L g741 ( .A(n_355), .Y(n_741) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_355), .Y(n_988) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_355), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_356), .B(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI31xp33_ASAP7_75t_L g607 ( .A1(n_358), .A2(n_608), .A3(n_617), .B(n_630), .Y(n_607) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_358), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g738 ( .A1(n_358), .A2(n_739), .A3(n_746), .B(n_755), .Y(n_738) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_358), .Y(n_1102) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND3x4_ASAP7_75t_L g585 ( .A(n_359), .B(n_380), .C(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g496 ( .A(n_360), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_371), .B2(n_372), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_364), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx8_ASAP7_75t_L g716 ( .A(n_365), .Y(n_716) );
INVx5_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g544 ( .A(n_366), .Y(n_544) );
INVx2_ASAP7_75t_SL g593 ( .A(n_366), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_366), .A2(n_588), .B1(n_691), .B2(n_692), .Y(n_690) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_366), .Y(n_933) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
INVx2_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
BUFx8_ASAP7_75t_L g568 ( .A(n_367), .Y(n_568) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
AND2x4_ASAP7_75t_L g402 ( .A(n_370), .B(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_372), .A2(n_392), .B1(n_562), .B2(n_563), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_372), .A2(n_675), .B1(n_676), .B2(n_677), .C(n_678), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_372), .A2(n_661), .B1(n_680), .B2(n_681), .C(n_682), .Y(n_679) );
CKINVDCx8_ASAP7_75t_R g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g396 ( .A(n_373), .Y(n_396) );
INVx3_ASAP7_75t_L g930 ( .A(n_373), .Y(n_930) );
INVx3_ASAP7_75t_L g934 ( .A(n_373), .Y(n_934) );
INVx3_ASAP7_75t_L g983 ( .A(n_373), .Y(n_983) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g776 ( .A(n_375), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_376), .A2(n_674), .B1(n_679), .B2(n_684), .Y(n_673) );
OAI33xp33_ASAP7_75t_L g768 ( .A1(n_376), .A2(n_769), .A3(n_777), .B1(n_784), .B2(n_787), .B3(n_788), .Y(n_768) );
OAI33xp33_ASAP7_75t_L g965 ( .A1(n_376), .A2(n_787), .A3(n_966), .B1(n_970), .B2(n_974), .B3(n_979), .Y(n_965) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_376), .A2(n_1050), .A3(n_1132), .B1(n_1138), .B2(n_1142), .B3(n_1146), .Y(n_1131) );
OAI33xp33_ASAP7_75t_L g1377 ( .A1(n_376), .A2(n_1050), .A3(n_1378), .B1(n_1382), .B2(n_1385), .B3(n_1388), .Y(n_1377) );
OAI33xp33_ASAP7_75t_L g1425 ( .A1(n_376), .A2(n_1050), .A3(n_1426), .B1(n_1429), .B2(n_1433), .B3(n_1436), .Y(n_1425) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx4f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_L g922 ( .A(n_378), .Y(n_922) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_378), .Y(n_1045) );
BUFx2_ASAP7_75t_L g569 ( .A(n_379), .Y(n_569) );
INVx1_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_380), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B1(n_388), .B2(n_389), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g558 ( .A(n_386), .Y(n_558) );
OR2x4_ASAP7_75t_L g703 ( .A(n_386), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g780 ( .A(n_386), .Y(n_780) );
OR2x4_ASAP7_75t_L g814 ( .A(n_386), .B(n_411), .Y(n_814) );
BUFx4f_ASAP7_75t_L g926 ( .A(n_386), .Y(n_926) );
INVx1_ASAP7_75t_L g403 ( .A(n_387), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_389), .A2(n_905), .B1(n_914), .B2(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_389), .A2(n_1140), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g783 ( .A(n_390), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B1(n_396), .B2(n_397), .C(n_398), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g675 ( .A(n_393), .Y(n_675) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_394), .Y(n_590) );
AND2x4_ASAP7_75t_L g816 ( .A(n_394), .B(n_704), .Y(n_816) );
INVx2_ASAP7_75t_L g972 ( .A(n_394), .Y(n_972) );
INVx1_ASAP7_75t_L g981 ( .A(n_394), .Y(n_981) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_401), .Y(n_1048) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_402), .B(n_433), .Y(n_448) );
INVx8_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_402), .Y(n_542) );
BUFx3_ASAP7_75t_L g718 ( .A(n_402), .Y(n_718) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g596 ( .A(n_405), .Y(n_596) );
INVx1_ASAP7_75t_L g719 ( .A(n_405), .Y(n_719) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
BUFx3_ASAP7_75t_L g537 ( .A(n_406), .Y(n_537) );
BUFx2_ASAP7_75t_L g550 ( .A(n_406), .Y(n_550) );
BUFx2_ASAP7_75t_L g683 ( .A(n_406), .Y(n_683) );
AND2x4_ASAP7_75t_L g705 ( .A(n_406), .B(n_411), .Y(n_705) );
BUFx2_ASAP7_75t_L g731 ( .A(n_406), .Y(n_731) );
BUFx2_ASAP7_75t_L g998 ( .A(n_406), .Y(n_998) );
INVx1_ASAP7_75t_L g442 ( .A(n_407), .Y(n_442) );
OAI33xp33_ASAP7_75t_L g921 ( .A1(n_408), .A2(n_922), .A3(n_923), .B1(n_927), .B2(n_931), .B3(n_935), .Y(n_921) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g684 ( .A(n_409), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_409), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_409), .A2(n_443), .B1(n_1104), .B2(n_1109), .C(n_1115), .Y(n_1103) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g1052 ( .A(n_410), .Y(n_1052) );
NAND3x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_414), .Y(n_410) );
AND2x4_ASAP7_75t_L g433 ( .A(n_411), .B(n_434), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_411), .B(n_414), .Y(n_560) );
INVx1_ASAP7_75t_L g704 ( .A(n_411), .Y(n_704) );
OR2x6_ASAP7_75t_L g832 ( .A(n_411), .B(n_776), .Y(n_832) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g427 ( .A(n_413), .Y(n_427) );
NAND2x1_ASAP7_75t_L g1071 ( .A(n_415), .B(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g680 ( .A(n_417), .Y(n_680) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g929 ( .A(n_418), .Y(n_929) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_418), .Y(n_1431) );
INVxp67_ASAP7_75t_L g1038 ( .A(n_419), .Y(n_1038) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_429), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g1058 ( .A1(n_422), .A2(n_1059), .B(n_1060), .Y(n_1058) );
INVx8_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g582 ( .A(n_424), .Y(n_582) );
INVx1_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
AND2x4_ASAP7_75t_L g432 ( .A(n_427), .B(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_445), .C(n_450), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_431), .A2(n_443), .B1(n_604), .B2(n_605), .C(n_606), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_431), .A2(n_443), .B1(n_605), .B2(n_734), .C(n_735), .Y(n_733) );
AND2x4_ASAP7_75t_SL g431 ( .A(n_432), .B(n_435), .Y(n_431) );
AND2x4_ASAP7_75t_L g438 ( .A(n_432), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g443 ( .A(n_432), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_432), .B(n_439), .Y(n_605) );
NAND2x1_ASAP7_75t_L g1042 ( .A(n_432), .B(n_435), .Y(n_1042) );
AND2x6_ASAP7_75t_L g531 ( .A(n_433), .B(n_435), .Y(n_531) );
AND2x2_ASAP7_75t_L g533 ( .A(n_433), .B(n_441), .Y(n_533) );
INVx1_ASAP7_75t_L g539 ( .A(n_433), .Y(n_539) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g1043 ( .A(n_438), .Y(n_1043) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_438), .A2(n_1075), .B1(n_1076), .B2(n_1077), .C(n_1078), .Y(n_1074) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_443), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_446), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_446), .B(n_737), .Y(n_736) );
INVx5_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
AND2x4_ASAP7_75t_L g580 ( .A(n_452), .B(n_454), .Y(n_580) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_453), .Y(n_536) );
INVx3_ASAP7_75t_L g571 ( .A(n_453), .Y(n_571) );
INVx8_ASAP7_75t_L g588 ( .A(n_453), .Y(n_588) );
AND2x4_ASAP7_75t_L g601 ( .A(n_454), .B(n_568), .Y(n_601) );
INVx3_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_644), .B2(n_760), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XOR2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_574), .Y(n_460) );
XNOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
NAND4xp75_ASAP7_75t_L g463 ( .A(n_464), .B(n_476), .C(n_521), .D(n_528), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g473 ( .A(n_470), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g664 ( .A(n_472), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_474), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_474), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g801 ( .A(n_474), .Y(n_801) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_474), .Y(n_804) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_475), .Y(n_505) );
AOI211x1_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_493), .B(n_498), .C(n_517), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g1013 ( .A(n_481), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_487), .B2(n_492), .Y(n_483) );
INVx1_ASAP7_75t_L g904 ( .A(n_485), .Y(n_904) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx3_ASAP7_75t_L g806 ( .A(n_486), .Y(n_806) );
INVx2_ASAP7_75t_SL g1026 ( .A(n_486), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g640 ( .A(n_489), .Y(n_640) );
INVx2_ASAP7_75t_L g749 ( .A(n_489), .Y(n_749) );
INVx1_ASAP7_75t_L g795 ( .A(n_489), .Y(n_795) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_489), .Y(n_808) );
INVx1_ASAP7_75t_L g1444 ( .A(n_489), .Y(n_1444) );
INVx8_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g858 ( .A(n_490), .B(n_848), .Y(n_858) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_492), .A2(n_506), .B1(n_556), .B2(n_558), .C(n_559), .Y(n_555) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_494), .A2(n_793), .A3(n_796), .B1(n_802), .B2(n_805), .B3(n_809), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g1149 ( .A1(n_494), .A2(n_915), .A3(n_1150), .B1(n_1154), .B2(n_1155), .B3(n_1156), .Y(n_1149) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g900 ( .A(n_495), .Y(n_900) );
INVx2_ASAP7_75t_L g990 ( .A(n_495), .Y(n_990) );
INVx4_ASAP7_75t_L g1392 ( .A(n_495), .Y(n_1392) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
OR2x6_ASAP7_75t_L g598 ( .A(n_496), .B(n_560), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_509), .B(n_513), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_504), .B2(n_506), .C(n_507), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g564 ( .A1(n_500), .A2(n_565), .B(n_567), .C(n_570), .Y(n_564) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g616 ( .A(n_503), .Y(n_616) );
BUFx3_ASAP7_75t_L g634 ( .A(n_503), .Y(n_634) );
BUFx2_ASAP7_75t_L g799 ( .A(n_503), .Y(n_799) );
BUFx2_ASAP7_75t_L g1395 ( .A(n_503), .Y(n_1395) );
OAI211xp5_ASAP7_75t_SL g654 ( .A1(n_504), .A2(n_655), .B(n_656), .C(n_659), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_504), .A2(n_661), .B(n_662), .C(n_663), .Y(n_660) );
BUFx4f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x6_ASAP7_75t_L g513 ( .A(n_505), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g612 ( .A(n_505), .Y(n_612) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_505), .Y(n_672) );
BUFx4f_ASAP7_75t_L g842 ( .A(n_505), .Y(n_842) );
BUFx4f_ASAP7_75t_L g910 ( .A(n_505), .Y(n_910) );
BUFx4f_ASAP7_75t_L g986 ( .A(n_505), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_509), .A2(n_985), .B1(n_989), .B2(n_991), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g809 ( .A(n_510), .Y(n_809) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2x2_ASAP7_75t_L g518 ( .A(n_515), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_525), .B2(n_526), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_522), .A2(n_525), .B1(n_542), .B2(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g1069 ( .A(n_523), .Y(n_1069) );
AND2x4_ASAP7_75t_L g526 ( .A(n_524), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g1072 ( .A(n_526), .Y(n_1072) );
OAI31xp67_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_540), .A3(n_554), .B(n_572), .Y(n_528) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_537), .C(n_538), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_537), .A2(n_666), .B1(n_688), .B2(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI21xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_545), .B(n_551), .Y(n_540) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_549), .B2(n_550), .Y(n_545) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
BUFx12f_ASAP7_75t_L g688 ( .A(n_548), .Y(n_688) );
INVx5_ASAP7_75t_L g729 ( .A(n_548), .Y(n_729) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI21xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_561), .B(n_564), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g890 ( .A(n_557), .Y(n_890) );
INVx2_ASAP7_75t_L g1108 ( .A(n_557), .Y(n_1108) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_558), .A2(n_782), .B1(n_785), .B2(n_786), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_558), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_558), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_565), .A2(n_926), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
OAI22xp33_ASAP7_75t_L g1378 ( .A1(n_565), .A2(n_1379), .B1(n_1380), .B2(n_1381), .Y(n_1378) );
OAI22xp33_ASAP7_75t_L g1426 ( .A1(n_565), .A2(n_938), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_568), .Y(n_1111) );
INVx3_ASAP7_75t_L g1143 ( .A(n_568), .Y(n_1143) );
INVx1_ASAP7_75t_L g1031 ( .A(n_572), .Y(n_1031) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_643), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_602), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_584), .C(n_599), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_580), .B2(n_581), .C1(n_582), .C2(n_583), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_578), .A2(n_580), .B1(n_582), .B2(n_723), .C1(n_724), .C2(n_725), .Y(n_722) );
AOI33xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .A3(n_589), .B1(n_591), .B2(n_595), .B3(n_597), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_585), .B(n_715), .C(n_717), .Y(n_714) );
BUFx3_ASAP7_75t_L g1115 ( .A(n_585), .Y(n_1115) );
INVx3_ASAP7_75t_L g693 ( .A(n_586), .Y(n_693) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_597), .B(n_727), .C(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_601), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g1039 ( .A(n_601), .Y(n_1039) );
NAND3xp33_ASAP7_75t_SL g602 ( .A(n_603), .B(n_607), .C(n_641), .Y(n_602) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_611), .A2(n_1094), .B(n_1095), .C(n_1096), .Y(n_1093) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g876 ( .A(n_612), .Y(n_876) );
INVx1_ASAP7_75t_L g1084 ( .A(n_612), .Y(n_1084) );
INVx2_ASAP7_75t_L g1446 ( .A(n_612), .Y(n_1446) );
OAI221xp5_ASAP7_75t_SL g985 ( .A1(n_615), .A2(n_971), .B1(n_980), .B2(n_986), .C(n_987), .Y(n_985) );
OAI221xp5_ASAP7_75t_SL g991 ( .A1(n_615), .A2(n_968), .B1(n_976), .B2(n_986), .C(n_992), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_615), .A2(n_1430), .B1(n_1434), .B2(n_1446), .Y(n_1445) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g745 ( .A(n_616), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B(n_624), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g746 ( .A1(n_618), .A2(n_747), .B(n_750), .Y(n_746) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_619), .A2(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_627), .A2(n_723), .B1(n_734), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_627), .A2(n_753), .B1(n_1076), .B2(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_SL g665 ( .A1(n_629), .A2(n_666), .B(n_667), .C(n_668), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g1081 ( .A1(n_629), .A2(n_667), .B(n_1082), .C(n_1083), .Y(n_1081) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_639), .B2(n_640), .Y(n_635) );
INVx4_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g1153 ( .A(n_638), .Y(n_1153) );
BUFx6f_ASAP7_75t_L g1442 ( .A(n_638), .Y(n_1442) );
INVx2_ASAP7_75t_L g907 ( .A(n_640), .Y(n_907) );
XNOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_711), .Y(n_644) );
XOR2xp5_ASAP7_75t_L g760 ( .A(n_645), .B(n_711), .Y(n_760) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_685), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B(n_673), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .C(n_660), .D(n_665), .Y(n_650) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g1448 ( .A(n_672), .Y(n_1448) );
OAI31xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_701), .A3(n_705), .B(n_706), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B(n_693), .C(n_694), .Y(n_686) );
AND2x4_ASAP7_75t_L g696 ( .A(n_693), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g699 ( .A(n_693), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g824 ( .A(n_693), .B(n_697), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_699), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_696), .A2(n_699), .B1(n_1455), .B2(n_1456), .Y(n_1454) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_699), .Y(n_826) );
BUFx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g829 ( .A(n_703), .Y(n_829) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_703), .Y(n_1000) );
CKINVDCx8_ASAP7_75t_R g821 ( .A(n_705), .Y(n_821) );
CKINVDCx8_ASAP7_75t_R g1453 ( .A(n_705), .Y(n_1453) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
AND2x2_ASAP7_75t_L g833 ( .A(n_707), .B(n_709), .Y(n_833) );
AND2x4_ASAP7_75t_L g897 ( .A(n_707), .B(n_709), .Y(n_897) );
AND2x2_ASAP7_75t_SL g1005 ( .A(n_707), .B(n_709), .Y(n_1005) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
XNOR2x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_759), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_732), .Y(n_712) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_714), .B(n_720), .C(n_722), .D(n_726), .Y(n_713) );
INVx1_ASAP7_75t_L g771 ( .A(n_716), .Y(n_771) );
INVx2_ASAP7_75t_L g1140 ( .A(n_716), .Y(n_1140) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND3xp33_ASAP7_75t_SL g732 ( .A(n_733), .B(n_736), .C(n_738), .Y(n_732) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_745), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_745), .A2(n_800), .B1(n_913), .B2(n_914), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_745), .A2(n_910), .B1(n_1139), .B2(n_1144), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_745), .A2(n_910), .B1(n_1135), .B2(n_1148), .Y(n_1155) );
OAI22xp33_ASAP7_75t_SL g1447 ( .A1(n_745), .A2(n_1428), .B1(n_1438), .B2(n_1448), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_941), .B1(n_1169), .B2(n_1170), .Y(n_762) );
INVxp67_ASAP7_75t_SL g1169 ( .A(n_763), .Y(n_1169) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_862), .B1(n_939), .B2(n_940), .Y(n_763) );
INVx1_ASAP7_75t_L g939 ( .A(n_764), .Y(n_939) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_810), .C(n_834), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_792), .Y(n_767) );
OAI22xp33_ASAP7_75t_SL g769 ( .A1(n_770), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_770), .A2(n_789), .B1(n_797), .B2(n_800), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_772), .A2(n_791), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx3_ASAP7_75t_L g790 ( .A(n_776), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_781), .B2(n_782), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_778), .A2(n_785), .B1(n_794), .B2(n_795), .Y(n_793) );
BUFx4f_ASAP7_75t_SL g1107 ( .A(n_779), .Y(n_1107) );
INVx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_SL g938 ( .A(n_780), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_781), .A2(n_786), .B1(n_803), .B2(n_804), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_782), .A2(n_902), .B1(n_913), .B2(n_924), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_782), .A2(n_1134), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g969 ( .A(n_783), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_790), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
INVx4_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g803 ( .A(n_798), .Y(n_803) );
INVx4_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_800), .A2(n_1383), .B1(n_1386), .B2(n_1395), .Y(n_1394) );
INVx5_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g1397 ( .A1(n_804), .A2(n_1025), .B1(n_1384), .B2(n_1387), .Y(n_1397) );
INVx6_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI31xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_817), .A3(n_828), .B(n_833), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_SL g887 ( .A(n_814), .Y(n_887) );
INVx1_ASAP7_75t_L g1004 ( .A(n_814), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_814), .Y(n_1160) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g888 ( .A(n_816), .Y(n_888) );
INVx2_ASAP7_75t_L g1161 ( .A(n_816), .Y(n_1161) );
INVx1_ASAP7_75t_L g1407 ( .A(n_816), .Y(n_1407) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g994 ( .A(n_821), .B(n_995), .C(n_999), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_822) );
AOI222xp33_ASAP7_75t_L g995 ( .A1(n_823), .A2(n_826), .B1(n_955), .B2(n_957), .C1(n_958), .C2(n_996), .Y(n_995) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx3_ASAP7_75t_L g892 ( .A(n_824), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_825), .A2(n_847), .B1(n_849), .B2(n_852), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_826), .A2(n_880), .B1(n_892), .B2(n_893), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_826), .A2(n_892), .B1(n_1124), .B2(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_826), .A2(n_892), .B1(n_1401), .B2(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx3_ASAP7_75t_L g895 ( .A(n_832), .Y(n_895) );
INVx2_ASAP7_75t_L g1001 ( .A(n_832), .Y(n_1001) );
OAI31xp33_ASAP7_75t_SL g1405 ( .A1(n_833), .A2(n_1406), .A3(n_1408), .B(n_1411), .Y(n_1405) );
OAI31xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_839), .A3(n_853), .B(n_859), .Y(n_834) );
CKINVDCx16_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
INVx3_ASAP7_75t_SL g874 ( .A(n_837), .Y(n_874) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx3_ASAP7_75t_L g883 ( .A(n_844), .Y(n_883) );
INVx1_ASAP7_75t_L g1122 ( .A(n_844), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_849), .A2(n_878), .B1(n_1455), .B2(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx3_ASAP7_75t_L g881 ( .A(n_851), .Y(n_881) );
INVx2_ASAP7_75t_L g960 ( .A(n_851), .Y(n_960) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g868 ( .A(n_855), .Y(n_868) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_855), .Y(n_1128) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g1129 ( .A(n_857), .Y(n_1129) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g872 ( .A(n_858), .Y(n_872) );
BUFx2_ASAP7_75t_L g953 ( .A(n_858), .Y(n_953) );
OAI31xp33_ASAP7_75t_SL g1398 ( .A1(n_859), .A2(n_1399), .A3(n_1403), .B(n_1404), .Y(n_1398) );
OAI31xp33_ASAP7_75t_SL g1459 ( .A1(n_859), .A2(n_1460), .A3(n_1462), .B(n_1465), .Y(n_1459) );
BUFx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g864 ( .A(n_860), .Y(n_864) );
BUFx2_ASAP7_75t_L g963 ( .A(n_860), .Y(n_963) );
OAI31xp33_ASAP7_75t_L g1120 ( .A1(n_860), .A2(n_1121), .A3(n_1126), .B(n_1127), .Y(n_1120) );
INVx1_ASAP7_75t_L g940 ( .A(n_862), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_884), .B2(n_896), .C(n_898), .Y(n_863) );
NOR3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_873), .C(n_875), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g1087 ( .A1(n_876), .A2(n_1088), .B(n_1089), .C(n_1091), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_880), .B1(n_881), .B2(n_882), .Y(n_877) );
AOI222xp33_ASAP7_75t_L g954 ( .A1(n_878), .A2(n_955), .B1(n_956), .B2(n_957), .C1(n_958), .C2(n_959), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_878), .A2(n_881), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_878), .A2(n_881), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
BUFx3_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_883), .B(n_948), .C(n_954), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_889), .C(n_894), .Y(n_884) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
CKINVDCx14_ASAP7_75t_R g896 ( .A(n_897), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_921), .Y(n_898) );
OAI33xp33_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .A3(n_908), .B1(n_912), .B2(n_915), .B3(n_918), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B1(n_905), .B2(n_906), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_903), .A2(n_906), .B1(n_919), .B2(n_920), .Y(n_918) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_906), .A2(n_1025), .B1(n_1027), .B2(n_1028), .C(n_1029), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_906), .A2(n_1133), .B1(n_1147), .B2(n_1151), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_906), .A2(n_1141), .B1(n_1145), .B2(n_1151), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_906), .A2(n_1151), .B1(n_1379), .B2(n_1389), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_906), .A2(n_1381), .B1(n_1390), .B2(n_1395), .Y(n_1396) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_909), .A2(n_919), .B1(n_928), .B2(n_930), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_911), .A2(n_920), .B1(n_932), .B2(n_934), .Y(n_931) );
OAI33xp33_ASAP7_75t_L g1391 ( .A1(n_915), .A2(n_1392), .A3(n_1393), .B1(n_1394), .B2(n_1396), .B3(n_1397), .Y(n_1391) );
OAI33xp33_ASAP7_75t_L g1439 ( .A1(n_915), .A2(n_989), .A3(n_1440), .B1(n_1445), .B2(n_1447), .B3(n_1449), .Y(n_1439) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
HB1xp67_ASAP7_75t_L g1380 ( .A(n_926), .Y(n_1380) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g1054 ( .A(n_929), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g1053 ( .A1(n_930), .A2(n_1054), .B1(n_1055), .B2(n_1056), .C(n_1057), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_930), .A2(n_1139), .B1(n_1140), .B2(n_1141), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_930), .A2(n_1143), .B1(n_1144), .B2(n_1145), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_930), .A2(n_972), .B1(n_1383), .B2(n_1384), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_930), .A2(n_1111), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1134 ( .A(n_937), .Y(n_1134) );
INVx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
OR2x6_ASAP7_75t_L g1037 ( .A(n_938), .B(n_1038), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1436 ( .A1(n_938), .A2(n_977), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
INVx1_ASAP7_75t_L g1170 ( .A(n_941), .Y(n_1170) );
OA22x2_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_943), .B1(n_1061), .B2(n_1062), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
XNOR2x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_1007), .Y(n_943) );
XOR2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_1006), .Y(n_944) );
NAND3x1_ASAP7_75t_L g945 ( .A(n_946), .B(n_964), .C(n_993), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_961), .B(n_963), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_950), .B1(n_951), .B2(n_952), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_949), .A2(n_951), .B1(n_1000), .B2(n_1001), .Y(n_999) );
INVx1_ASAP7_75t_L g1466 ( .A(n_952), .Y(n_1466) );
INVx2_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NOR2x1_ASAP7_75t_L g964 ( .A(n_965), .B(n_984), .Y(n_964) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1137 ( .A(n_978), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_983), .A2(n_1380), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
OAI22xp5_ASAP7_75t_L g1429 ( .A1(n_983), .A2(n_1430), .B1(n_1431), .B2(n_1432), .Y(n_1429) );
BUFx6f_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
OAI21xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_1002), .B(n_1005), .Y(n_993) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1000), .Y(n_1166) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1000), .Y(n_1458) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_1005), .A2(n_1158), .A3(n_1162), .B(n_1165), .Y(n_1157) );
OAI31xp33_ASAP7_75t_L g1450 ( .A1(n_1005), .A2(n_1451), .A3(n_1452), .B(n_1457), .Y(n_1450) );
O2A1O1Ixp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1019), .B(n_1031), .C(n_1032), .Y(n_1008) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1021), .Y(n_1100) );
INVx4_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
OAI21xp5_ASAP7_75t_L g1046 ( .A1(n_1027), .A2(n_1047), .B(n_1049), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1040), .C(n_1058), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1036), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1037), .B(n_1069), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1044), .Y(n_1040) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1042), .Y(n_1075) );
OAI22xp5_ASAP7_75t_SL g1044 ( .A1(n_1045), .A2(n_1046), .B1(n_1050), .B2(n_1053), .Y(n_1044) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
AO22x2_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1116), .B1(n_1117), .B2(n_1168), .Y(n_1062) );
INVx1_ASAP7_75t_SL g1168 ( .A(n_1063), .Y(n_1168) );
XNOR2x1_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NOR2x1_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1073), .Y(n_1065) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NAND3xp33_ASAP7_75t_SL g1073 ( .A(n_1074), .B(n_1079), .C(n_1103), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1097), .B(n_1101), .Y(n_1079) );
NAND3xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1087), .C(n_1093), .Y(n_1080) );
NAND2xp5_ASAP7_75t_SL g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_1094), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1105) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1130), .C(n_1157), .Y(n_1119) );
NOR2xp33_ASAP7_75t_SL g1130 ( .A(n_1131), .B(n_1149), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1134), .B1(n_1135), .B2(n_1136), .Y(n_1132) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx2_ASAP7_75t_SL g1152 ( .A(n_1153), .Y(n_1152) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_1160), .Y(n_1159) );
OAI221xp5_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1371), .B1(n_1374), .B2(n_1412), .C(n_1417), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1326), .Y(n_1172) );
NAND3xp33_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1265), .C(n_1295), .Y(n_1173) );
AOI211xp5_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1195), .B(n_1228), .C(n_1245), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1175), .B(n_1269), .Y(n_1268) );
AOI322xp5_ASAP7_75t_L g1277 ( .A1(n_1175), .A2(n_1203), .A3(n_1226), .B1(n_1230), .B2(n_1273), .C1(n_1278), .C2(n_1281), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1191), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1176), .B(n_1307), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1176), .B(n_1308), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1176), .B(n_1219), .Y(n_1363) );
INVx3_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1177), .B(n_1233), .Y(n_1232) );
INVx3_ASAP7_75t_L g1244 ( .A(n_1177), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1177), .B(n_1191), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1177), .B(n_1294), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1177), .B(n_1269), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1177), .B(n_1274), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1177), .B(n_1253), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1177), .B(n_1191), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1177), .B(n_1367), .Y(n_1366) );
AND2x4_ASAP7_75t_SL g1177 ( .A(n_1178), .B(n_1185), .Y(n_1177) );
AND2x6_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1181), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1180), .B(n_1184), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_1180), .B(n_1187), .Y(n_1186) );
AND2x6_ASAP7_75t_L g1189 ( .A(n_1180), .B(n_1190), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1180), .B(n_1184), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1180), .B(n_1184), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1182), .B(n_1188), .Y(n_1187) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1189), .Y(n_1373) );
OAI21xp5_ASAP7_75t_L g1467 ( .A1(n_1190), .A2(n_1468), .B(n_1469), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1191), .B(n_1225), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1191), .B(n_1216), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1191), .B(n_1216), .Y(n_1308) );
OAI221xp5_ASAP7_75t_SL g1332 ( .A1(n_1191), .A2(n_1196), .B1(n_1333), .B2(n_1334), .C(n_1335), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1194), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1231 ( .A(n_1192), .B(n_1194), .Y(n_1231) );
A2O1A1Ixp33_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1210), .B(n_1214), .C(n_1222), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1196), .B(n_1238), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1196), .B(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1197), .B(n_1226), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1203), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1198), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1198), .B(n_1248), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1198), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1198), .B(n_1303), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1198), .B(n_1319), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1198), .B(n_1240), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1199), .B(n_1203), .Y(n_1227) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_1199), .B(n_1219), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1199), .B(n_1207), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1199), .B(n_1240), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1199), .B(n_1219), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1199), .B(n_1303), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1202), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1200), .B(n_1202), .Y(n_1285) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1203), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1203), .B(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1207), .Y(n_1203) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1204), .Y(n_1213) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1204), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1206), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1207), .B(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1207), .Y(n_1249) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1207), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1207), .B(n_1213), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
NOR2xp33_ASAP7_75t_L g1351 ( .A(n_1210), .B(n_1352), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1211), .B(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1212), .B(n_1259), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1213), .B(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1213), .Y(n_1303) );
INVxp33_ASAP7_75t_SL g1301 ( .A(n_1214), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1219), .Y(n_1214) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1215), .Y(n_1260) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1215), .Y(n_1329) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1216), .Y(n_1225) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1216), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
INVx3_ASAP7_75t_L g1226 ( .A(n_1219), .Y(n_1226) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1219), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1219), .B(n_1225), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1219), .B(n_1310), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1227), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1224), .B(n_1300), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1226), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1225), .B(n_1231), .Y(n_1230) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1226), .B(n_1233), .C(n_1239), .Y(n_1254) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1226), .Y(n_1259) );
NOR2xp33_ASAP7_75t_L g1281 ( .A(n_1226), .B(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1226), .B(n_1316), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1226), .B(n_1302), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1227), .B(n_1242), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1227), .B(n_1270), .Y(n_1276) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1227), .Y(n_1313) );
OAI21xp5_ASAP7_75t_L g1359 ( .A1(n_1227), .A2(n_1360), .B(n_1361), .Y(n_1359) );
OAI21xp33_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1239), .B(n_1241), .Y(n_1228) );
NAND3xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1232), .C(n_1237), .Y(n_1229) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1230), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_1231), .A2(n_1299), .B1(n_1301), .B2(n_1302), .Y(n_1298) );
OAI211xp5_ASAP7_75t_L g1317 ( .A1(n_1231), .A2(n_1318), .B(n_1320), .C(n_1324), .Y(n_1317) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1231), .Y(n_1367) );
OAI21xp33_ASAP7_75t_L g1327 ( .A1(n_1232), .A2(n_1328), .B(n_1332), .Y(n_1327) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1234), .Y(n_1243) );
OAI31xp33_ASAP7_75t_SL g1295 ( .A1(n_1234), .A2(n_1296), .A3(n_1305), .B(n_1317), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1237), .B(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
NAND2xp5_ASAP7_75t_SL g1319 ( .A(n_1238), .B(n_1279), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1238), .B(n_1307), .Y(n_1358) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1242), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1243), .Y(n_1262) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1244), .Y(n_1304) );
OAI221xp5_ASAP7_75t_L g1245 ( .A1(n_1246), .A2(n_1251), .B1(n_1252), .B2(n_1254), .C(n_1255), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1250), .Y(n_1247) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1248), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1248), .B(n_1285), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1250), .B(n_1279), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1250), .B(n_1264), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_1251), .Y(n_1294) );
OAI322xp33_ASAP7_75t_L g1283 ( .A1(n_1252), .A2(n_1284), .A3(n_1286), .B1(n_1287), .B2(n_1288), .C1(n_1290), .C2(n_1292), .Y(n_1283) );
CKINVDCx14_ASAP7_75t_R g1252 ( .A(n_1253), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1253), .B(n_1259), .Y(n_1322) );
NAND4xp25_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1258), .C(n_1261), .D(n_1263), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1314 ( .A1(n_1256), .A2(n_1315), .B(n_1316), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1256), .B(n_1331), .Y(n_1353) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1259), .B(n_1275), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1259), .B(n_1294), .Y(n_1340) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1259), .B(n_1369), .Y(n_1368) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_1261), .A2(n_1266), .B1(n_1268), .B2(n_1271), .C(n_1283), .Y(n_1265) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_1263), .A2(n_1273), .B1(n_1279), .B2(n_1294), .C(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI21xp33_ASAP7_75t_L g1272 ( .A1(n_1268), .A2(n_1273), .B(n_1275), .Y(n_1272) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1269), .Y(n_1334) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NAND3xp33_ASAP7_75t_SL g1271 ( .A(n_1272), .B(n_1276), .C(n_1277), .Y(n_1271) );
CKINVDCx14_ASAP7_75t_R g1273 ( .A(n_1274), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1278), .B(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1279), .B(n_1285), .Y(n_1291) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1282), .Y(n_1323) );
OAI21xp33_ASAP7_75t_L g1356 ( .A1(n_1282), .A2(n_1357), .B(n_1359), .Y(n_1356) );
OAI321xp33_ASAP7_75t_L g1305 ( .A1(n_1285), .A2(n_1306), .A3(n_1309), .B1(n_1311), .B2(n_1313), .C(n_1314), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1285), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
AOI21xp33_ASAP7_75t_L g1296 ( .A1(n_1297), .A2(n_1298), .B(n_1304), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1300), .B(n_1310), .Y(n_1309) );
AOI211xp5_ASAP7_75t_L g1354 ( .A1(n_1307), .A2(n_1355), .B(n_1356), .C(n_1364), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1307), .B(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_1311), .A2(n_1365), .B1(n_1368), .B2(n_1370), .Y(n_1364) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1316), .Y(n_1339) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1322), .B(n_1323), .Y(n_1320) );
NAND4xp25_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1337), .C(n_1350), .D(n_1354), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1334), .B(n_1348), .Y(n_1347) );
AOI211xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1340), .B(n_1341), .C(n_1346), .Y(n_1337) );
AOI21xp33_ASAP7_75t_SL g1341 ( .A1(n_1342), .A2(n_1344), .B(n_1345), .Y(n_1341) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1342), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1345), .B(n_1347), .Y(n_1346) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1353), .Y(n_1350) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
CKINVDCx20_ASAP7_75t_R g1371 ( .A(n_1372), .Y(n_1371) );
CKINVDCx20_ASAP7_75t_R g1372 ( .A(n_1373), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1398), .C(n_1405), .Y(n_1375) );
NOR2xp33_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1391), .Y(n_1376) );
CKINVDCx20_ASAP7_75t_R g1412 ( .A(n_1413), .Y(n_1412) );
CKINVDCx20_ASAP7_75t_R g1413 ( .A(n_1414), .Y(n_1413) );
INVx3_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
HB1xp67_ASAP7_75t_SL g1418 ( .A(n_1419), .Y(n_1418) );
INVxp33_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
NAND3xp33_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1450), .C(n_1459), .Y(n_1423) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1439), .Y(n_1424) );
OAI22xp33_ASAP7_75t_L g1440 ( .A1(n_1427), .A2(n_1437), .B1(n_1441), .B2(n_1443), .Y(n_1440) );
OAI22xp33_ASAP7_75t_L g1449 ( .A1(n_1432), .A2(n_1435), .B1(n_1441), .B2(n_1443), .Y(n_1449) );
INVx2_ASAP7_75t_SL g1441 ( .A(n_1442), .Y(n_1441) );
BUFx3_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
endmodule