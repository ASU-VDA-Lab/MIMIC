module fake_ariane_1873_n_89 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_89);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_89;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_47;
wire n_86;
wire n_75;
wire n_67;
wire n_69;
wire n_74;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_46;
wire n_84;
wire n_72;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_55;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_63;
wire n_59;
wire n_54;

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_7),
.Y(n_46)
);

OAI21x1_ASAP7_75t_L g47 ( 
.A1(n_18),
.A2(n_38),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_6),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_31),
.B1(n_21),
.B2(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_35),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_1),
.B(n_11),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_15),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_22),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_55),
.B1(n_43),
.B2(n_52),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_47),
.B(n_50),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_56),
.C(n_51),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_48),
.B(n_46),
.C(n_51),
.Y(n_69)
);

AO31x2_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_41),
.A3(n_56),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_23),
.B(n_26),
.Y(n_72)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_76),
.Y(n_80)
);

NAND2x1p5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_74),
.Y(n_82)
);

OAI222xp33_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_78),
.B1(n_79),
.B2(n_74),
.C1(n_72),
.C2(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_86),
.Y(n_88)
);

OR2x6_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_32),
.Y(n_89)
);


endmodule