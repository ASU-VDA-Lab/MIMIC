module real_aes_6493_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g481 ( .A1(n_0), .A2(n_164), .B(n_482), .C(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_1), .B(n_476), .Y(n_487) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_91), .C(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g202 ( .A(n_3), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_4), .B(n_165), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g142 ( .A1(n_5), .A2(n_143), .B1(n_144), .B2(n_450), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_5), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_5), .A2(n_98), .B1(n_450), .B2(n_750), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_6), .A2(n_461), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_7), .A2(n_171), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_8), .A2(n_38), .B1(n_168), .B2(n_220), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_9), .B(n_171), .Y(n_188) );
AND2x6_ASAP7_75t_L g173 ( .A(n_10), .B(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_11), .A2(n_173), .B(n_464), .C(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_12), .B(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
INVx1_ASAP7_75t_L g194 ( .A(n_14), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_15), .B(n_161), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_16), .A2(n_41), .B1(n_536), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_16), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_17), .B(n_165), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_18), .B(n_151), .Y(n_150) );
AO32x2_ASAP7_75t_L g231 ( .A1(n_19), .A2(n_171), .A3(n_172), .B1(n_191), .B2(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_20), .B(n_168), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_21), .B(n_151), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_22), .A2(n_54), .B1(n_168), .B2(n_220), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g228 ( .A1(n_23), .A2(n_83), .B1(n_161), .B2(n_168), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_24), .B(n_168), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_25), .A2(n_172), .B(n_464), .C(n_466), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_26), .A2(n_172), .B(n_464), .C(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_27), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_28), .A2(n_99), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_28), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_29), .B(n_210), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_30), .A2(n_461), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_31), .B(n_210), .Y(n_247) );
INVx2_ASAP7_75t_L g163 ( .A(n_32), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_33), .A2(n_496), .B(n_497), .C(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_34), .B(n_168), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_35), .B(n_210), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_36), .A2(n_135), .B1(n_138), .B2(n_139), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_36), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_37), .B(n_216), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_40), .B(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_41), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_42), .B(n_165), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_43), .B(n_461), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_44), .A2(n_496), .B(n_501), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_45), .B(n_168), .Y(n_181) );
INVx1_ASAP7_75t_L g483 ( .A(n_46), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_47), .A2(n_752), .B1(n_753), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g755 ( .A(n_47), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_48), .A2(n_92), .B1(n_220), .B2(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g522 ( .A(n_49), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_50), .B(n_168), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_51), .B(n_168), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_52), .B(n_461), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_53), .B(n_186), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g167 ( .A1(n_55), .A2(n_60), .B1(n_161), .B2(n_168), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_56), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_56), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_57), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_58), .B(n_168), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_59), .B(n_168), .Y(n_267) );
INVx1_ASAP7_75t_L g174 ( .A(n_61), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_62), .B(n_461), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_63), .B(n_476), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_64), .A2(n_186), .B(n_197), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_65), .B(n_168), .Y(n_203) );
INVx1_ASAP7_75t_L g154 ( .A(n_66), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_68), .B(n_165), .Y(n_499) );
AO32x2_ASAP7_75t_L g224 ( .A1(n_69), .A2(n_171), .A3(n_172), .B1(n_225), .B2(n_229), .Y(n_224) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_70), .A2(n_130), .B1(n_131), .B2(n_140), .C1(n_735), .C2(n_741), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_71), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_72), .B(n_166), .Y(n_533) );
INVx1_ASAP7_75t_L g266 ( .A(n_73), .Y(n_266) );
INVx1_ASAP7_75t_L g242 ( .A(n_74), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_75), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_76), .B(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_77), .A2(n_464), .B(n_501), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_78), .B(n_161), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_79), .Y(n_509) );
INVx1_ASAP7_75t_L g114 ( .A(n_80), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_81), .A2(n_106), .B1(n_115), .B2(n_757), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_82), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_84), .B(n_220), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_85), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_86), .B(n_161), .Y(n_246) );
INVx2_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_88), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_89), .B(n_158), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_90), .B(n_161), .Y(n_182) );
OR2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g451 ( .A(n_91), .B(n_125), .Y(n_451) );
INVx2_ASAP7_75t_L g734 ( .A(n_91), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_93), .A2(n_104), .B1(n_161), .B2(n_162), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_94), .B(n_461), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_95), .Y(n_498) );
INVxp67_ASAP7_75t_L g512 ( .A(n_96), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_97), .B(n_161), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_98), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_99), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g529 ( .A(n_101), .Y(n_529) );
INVx1_ASAP7_75t_L g558 ( .A(n_102), .Y(n_558) );
AND2x2_ASAP7_75t_L g524 ( .A(n_103), .B(n_210), .Y(n_524) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_107), .Y(n_758) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_129), .B1(n_744), .B2(n_745), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g744 ( .A(n_118), .Y(n_744) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_120), .A2(n_746), .B(n_756), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_128), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_123), .Y(n_756) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_124), .B(n_734), .Y(n_743) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g733 ( .A(n_125), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_135), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_451), .B1(n_452), .B2(n_733), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_142), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_144), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_384), .Y(n_144) );
NOR5xp2_ASAP7_75t_L g145 ( .A(n_146), .B(n_297), .C(n_343), .D(n_356), .E(n_368), .Y(n_145) );
OAI211xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_205), .B(n_251), .C(n_278), .Y(n_146) );
INVx1_ASAP7_75t_SL g379 ( .A(n_147), .Y(n_379) );
OR2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_175), .Y(n_147) );
AND2x2_ASAP7_75t_L g303 ( .A(n_148), .B(n_176), .Y(n_303) );
AND2x2_ASAP7_75t_L g331 ( .A(n_148), .B(n_277), .Y(n_331) );
AND2x2_ASAP7_75t_L g339 ( .A(n_148), .B(n_282), .Y(n_339) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g269 ( .A(n_149), .B(n_177), .Y(n_269) );
INVx2_ASAP7_75t_L g281 ( .A(n_149), .Y(n_281) );
AND2x2_ASAP7_75t_L g406 ( .A(n_149), .B(n_348), .Y(n_406) );
OR2x2_ASAP7_75t_L g408 ( .A(n_149), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_156), .Y(n_149) );
INVx1_ASAP7_75t_L g275 ( .A(n_150), .Y(n_275) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx1_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_152), .B(n_153), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NAND3xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_170), .C(n_172), .Y(n_156) );
AO21x1_ASAP7_75t_L g274 ( .A1(n_157), .A2(n_170), .B(n_275), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B1(n_164), .B2(n_167), .Y(n_157) );
INVx2_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g225 ( .A1(n_158), .A2(n_166), .B1(n_226), .B2(n_228), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_158), .A2(n_164), .B1(n_233), .B2(n_234), .Y(n_232) );
INVx4_ASAP7_75t_L g484 ( .A(n_158), .Y(n_484) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
INVx1_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
AND2x2_ASAP7_75t_L g462 ( .A(n_159), .B(n_187), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_159), .Y(n_465) );
INVx2_ASAP7_75t_L g195 ( .A(n_161), .Y(n_195) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
INVx1_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_184), .B(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_202), .C(n_203), .Y(n_200) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_181), .B(n_182), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_SL g240 ( .A1(n_165), .A2(n_241), .B(n_242), .C(n_243), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_165), .A2(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_165), .B(n_512), .Y(n_511) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_168), .Y(n_560) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
BUFx3_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
AND2x6_ASAP7_75t_L g464 ( .A(n_169), .B(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g476 ( .A(n_170), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_170), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_170), .A2(n_528), .B(n_535), .Y(n_527) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_170), .A2(n_555), .B(n_562), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_170), .B(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_171), .A2(n_179), .B(n_188), .Y(n_178) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_171), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_171), .A2(n_540), .B(n_541), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_172), .A2(n_262), .B(n_265), .Y(n_261) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_173), .A2(n_180), .B(n_183), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_173), .A2(n_193), .B(n_200), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_173), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_173), .A2(n_240), .B(n_244), .Y(n_239) );
AND2x4_ASAP7_75t_L g461 ( .A(n_173), .B(n_462), .Y(n_461) );
INVx4_ASAP7_75t_SL g486 ( .A(n_173), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_173), .B(n_462), .Y(n_530) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g319 ( .A(n_176), .B(n_291), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_176), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g433 ( .A(n_176), .B(n_273), .Y(n_433) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_189), .Y(n_176) );
AND2x2_ASAP7_75t_L g276 ( .A(n_177), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g323 ( .A(n_177), .Y(n_323) );
AND2x2_ASAP7_75t_L g348 ( .A(n_177), .B(n_260), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_177), .B(n_381), .Y(n_418) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g282 ( .A(n_178), .B(n_260), .Y(n_282) );
AND2x2_ASAP7_75t_L g296 ( .A(n_178), .B(n_259), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_178), .B(n_189), .Y(n_313) );
AND2x2_ASAP7_75t_L g370 ( .A(n_178), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_178), .B(n_277), .Y(n_383) );
AND2x2_ASAP7_75t_L g435 ( .A(n_178), .B(n_360), .Y(n_435) );
INVx2_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g258 ( .A(n_189), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_189), .B(n_260), .Y(n_354) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_204), .Y(n_189) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_190), .A2(n_261), .B(n_268), .Y(n_260) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_191), .B(n_536), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .C(n_197), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_195), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_195), .A2(n_543), .B(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_197), .A2(n_558), .B(n_559), .C(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_245), .B(n_246), .Y(n_244) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g468 ( .A(n_199), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g265 ( .A1(n_201), .A2(n_221), .B(n_266), .C(n_267), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_201), .A2(n_467), .B(n_469), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_235), .B(n_248), .Y(n_205) );
INVx1_ASAP7_75t_SL g367 ( .A(n_206), .Y(n_367) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_223), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_208), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g250 ( .A(n_209), .Y(n_250) );
INVx1_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
AND2x2_ASAP7_75t_L g308 ( .A(n_209), .B(n_230), .Y(n_308) );
AND2x2_ASAP7_75t_L g342 ( .A(n_209), .B(n_231), .Y(n_342) );
OR2x2_ASAP7_75t_L g361 ( .A(n_209), .B(n_237), .Y(n_361) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_209), .Y(n_375) );
AND2x2_ASAP7_75t_L g388 ( .A(n_209), .B(n_389), .Y(n_388) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_222), .Y(n_209) );
INVx2_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_210), .A2(n_239), .B(n_247), .Y(n_238) );
INVx1_ASAP7_75t_L g474 ( .A(n_210), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_210), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_210), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_221), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_223), .A2(n_310), .B1(n_311), .B2(n_320), .Y(n_309) );
AND2x2_ASAP7_75t_L g393 ( .A(n_223), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
INVx1_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
INVx1_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
AND2x2_ASAP7_75t_L g317 ( .A(n_224), .B(n_231), .Y(n_317) );
INVx2_ASAP7_75t_L g485 ( .A(n_227), .Y(n_485) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_227), .Y(n_500) );
INVx1_ASAP7_75t_L g471 ( .A(n_229), .Y(n_471) );
OR2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_256), .Y(n_271) );
AND2x2_ASAP7_75t_L g301 ( .A(n_230), .B(n_302), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_230), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g249 ( .A(n_231), .B(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g358 ( .A(n_231), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_235), .B(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g336 ( .A(n_236), .B(n_302), .Y(n_336) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g248 ( .A(n_237), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g307 ( .A(n_237), .Y(n_307) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g256 ( .A(n_238), .Y(n_256) );
OR2x2_ASAP7_75t_L g286 ( .A(n_238), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_238), .Y(n_341) );
AOI32xp33_ASAP7_75t_L g378 ( .A1(n_248), .A2(n_308), .A3(n_379), .B1(n_380), .B2(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g304 ( .A(n_249), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_249), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_249), .B(n_336), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_249), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_257), .B1(n_270), .B2(n_272), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_254), .B(n_256), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_255), .A2(n_279), .B1(n_283), .B2(n_293), .Y(n_278) );
AND2x2_ASAP7_75t_L g300 ( .A(n_255), .B(n_301), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_255), .A2(n_269), .B(n_317), .C(n_352), .Y(n_351) );
OAI332xp33_ASAP7_75t_L g356 ( .A1(n_255), .A2(n_357), .A3(n_359), .B1(n_361), .B2(n_362), .B3(n_364), .C1(n_365), .C2(n_367), .Y(n_356) );
INVx2_ASAP7_75t_L g397 ( .A(n_255), .Y(n_397) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
INVx1_ASAP7_75t_L g390 ( .A(n_256), .Y(n_390) );
AND2x2_ASAP7_75t_L g444 ( .A(n_256), .B(n_308), .Y(n_444) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_269), .Y(n_257) );
AND2x2_ASAP7_75t_L g324 ( .A(n_259), .B(n_274), .Y(n_324) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_260), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g372 ( .A(n_260), .B(n_274), .Y(n_372) );
INVx1_ASAP7_75t_L g381 ( .A(n_260), .Y(n_381) );
INVx1_ASAP7_75t_L g355 ( .A(n_269), .Y(n_355) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g439 ( .A(n_271), .B(n_291), .Y(n_439) );
INVx1_ASAP7_75t_SL g350 ( .A(n_272), .Y(n_350) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
AND2x2_ASAP7_75t_L g377 ( .A(n_273), .B(n_335), .Y(n_377) );
INVx1_ASAP7_75t_L g396 ( .A(n_273), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_273), .B(n_363), .Y(n_398) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
AND2x2_ASAP7_75t_L g299 ( .A(n_276), .B(n_280), .Y(n_299) );
AND2x2_ASAP7_75t_L g366 ( .A(n_276), .B(n_324), .Y(n_366) );
INVx2_ASAP7_75t_L g409 ( .A(n_276), .Y(n_409) );
INVx2_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
AND2x2_ASAP7_75t_L g294 ( .A(n_277), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_281), .B(n_354), .Y(n_360) );
OR2x2_ASAP7_75t_L g424 ( .A(n_281), .B(n_383), .Y(n_424) );
INVx1_ASAP7_75t_L g448 ( .A(n_281), .Y(n_448) );
INVx1_ASAP7_75t_L g404 ( .A(n_282), .Y(n_404) );
AND2x2_ASAP7_75t_L g449 ( .A(n_282), .B(n_292), .Y(n_449) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_286), .A2(n_312), .B1(n_314), .B2(n_318), .Y(n_311) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI322xp33_ASAP7_75t_SL g395 ( .A1(n_289), .A2(n_396), .A3(n_397), .B1(n_398), .B2(n_399), .C1(n_402), .C2(n_404), .Y(n_395) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x2_ASAP7_75t_L g392 ( .A(n_290), .B(n_308), .Y(n_392) );
OR2x2_ASAP7_75t_L g426 ( .A(n_290), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g429 ( .A(n_290), .B(n_361), .Y(n_429) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g374 ( .A(n_291), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g430 ( .A(n_291), .B(n_361), .Y(n_430) );
INVx3_ASAP7_75t_L g363 ( .A(n_292), .Y(n_363) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g419 ( .A(n_294), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g298 ( .A1(n_296), .A2(n_299), .B1(n_300), .B2(n_303), .C1(n_304), .C2(n_306), .Y(n_298) );
INVx1_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
NAND3xp33_ASAP7_75t_SL g297 ( .A(n_298), .B(n_309), .C(n_326), .Y(n_297) );
AND2x2_ASAP7_75t_L g414 ( .A(n_301), .B(n_315), .Y(n_414) );
BUFx2_ASAP7_75t_L g305 ( .A(n_302), .Y(n_305) );
INVx1_ASAP7_75t_L g346 ( .A(n_302), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_303), .A2(n_339), .B1(n_392), .B2(n_393), .C(n_395), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_305), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_313), .B(n_324), .Y(n_325) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
OAI21xp33_ASAP7_75t_L g320 ( .A1(n_315), .A2(n_321), .B(n_325), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_315), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g412 ( .A(n_317), .B(n_394), .Y(n_412) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g335 ( .A(n_323), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_324), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g441 ( .A(n_324), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_332), .B1(n_333), .B2(n_336), .C(n_337), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_328), .B(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g437 ( .A(n_336), .B(n_342), .Y(n_437) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OAI31xp33_ASAP7_75t_SL g405 ( .A1(n_340), .A2(n_379), .A3(n_406), .B(n_407), .Y(n_405) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g394 ( .A(n_341), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_342), .B(n_346), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_351), .Y(n_343) );
INVx1_ASAP7_75t_L g349 ( .A(n_345), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_348), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g364 ( .A(n_357), .Y(n_364) );
INVx2_ASAP7_75t_L g400 ( .A(n_358), .Y(n_400) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g386 ( .A(n_363), .B(n_372), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_363), .A2(n_380), .B(n_437), .C(n_438), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g368 ( .A1(n_364), .A2(n_369), .B1(n_373), .B2(n_376), .C(n_378), .Y(n_368) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_367), .A2(n_432), .B(n_434), .C(n_436), .Y(n_431) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_428), .Y(n_420) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NOR4xp25_ASAP7_75t_L g384 ( .A(n_385), .B(n_410), .C(n_431), .D(n_442), .Y(n_384) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .B(n_391), .C(n_405), .Y(n_385) );
INVx1_ASAP7_75t_SL g440 ( .A(n_392), .Y(n_440) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_SL g403 ( .A(n_401), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_408), .A2(n_417), .B1(n_429), .B2(n_430), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_415), .C(n_420), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI31xp33_ASAP7_75t_L g442 ( .A1(n_413), .A2(n_443), .A3(n_445), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g737 ( .A(n_451), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_452), .Y(n_738) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_453), .B(n_669), .Y(n_452) );
NOR5xp2_ASAP7_75t_L g453 ( .A(n_454), .B(n_600), .C(n_629), .D(n_649), .E(n_656), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_488), .B(n_545), .C(n_587), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_456), .A2(n_672), .B1(n_674), .B2(n_675), .Y(n_671) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_475), .Y(n_456) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_457), .Y(n_548) );
AND2x4_ASAP7_75t_L g580 ( .A(n_457), .B(n_581), .Y(n_580) );
INVx5_ASAP7_75t_L g598 ( .A(n_457), .Y(n_598) );
AND2x2_ASAP7_75t_L g607 ( .A(n_457), .B(n_599), .Y(n_607) );
AND2x2_ASAP7_75t_L g619 ( .A(n_457), .B(n_492), .Y(n_619) );
AND2x2_ASAP7_75t_L g715 ( .A(n_457), .B(n_583), .Y(n_715) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_472), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_463), .B(n_471), .Y(n_458) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx5_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
INVx2_ASAP7_75t_L g470 ( .A(n_468), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_470), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_470), .A2(n_500), .B(n_522), .C(n_523), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g581 ( .A(n_475), .Y(n_581) );
AND2x2_ASAP7_75t_L g599 ( .A(n_475), .B(n_554), .Y(n_599) );
AND2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_553), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_475), .B(n_598), .Y(n_658) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_487), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B(n_481), .C(n_486), .Y(n_478) );
INVx2_ASAP7_75t_L g496 ( .A(n_480), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_480), .A2(n_486), .B(n_509), .C(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g501 ( .A(n_486), .Y(n_501) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_514), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI322xp5_ASAP7_75t_L g717 ( .A1(n_491), .A2(n_525), .A3(n_572), .B1(n_580), .B2(n_634), .C1(n_718), .C2(n_721), .Y(n_717) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_504), .Y(n_491) );
INVx5_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
AND2x2_ASAP7_75t_L g566 ( .A(n_492), .B(n_552), .Y(n_566) );
BUFx2_ASAP7_75t_L g644 ( .A(n_492), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_492), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g721 ( .A(n_492), .B(n_628), .Y(n_721) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_504), .B(n_516), .Y(n_575) );
INVx1_ASAP7_75t_L g602 ( .A(n_504), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_504), .B(n_537), .Y(n_615) );
AND2x2_ASAP7_75t_L g716 ( .A(n_504), .B(n_634), .Y(n_716) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_516), .Y(n_570) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_505), .Y(n_578) );
OR2x2_ASAP7_75t_L g585 ( .A(n_505), .B(n_537), .Y(n_585) );
AND2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_505), .B(n_527), .Y(n_624) );
INVxp67_ASAP7_75t_L g648 ( .A(n_505), .Y(n_648) );
AND2x2_ASAP7_75t_L g655 ( .A(n_505), .B(n_525), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_505), .B(n_537), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_505), .B(n_526), .Y(n_681) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_516), .B(n_538), .Y(n_625) );
OR2x2_ASAP7_75t_L g647 ( .A(n_516), .B(n_526), .Y(n_647) );
AND2x2_ASAP7_75t_L g660 ( .A(n_516), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_516), .B(n_615), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_516), .A2(n_671), .B(n_676), .C(n_685), .Y(n_670) );
AND2x2_ASAP7_75t_L g731 ( .A(n_516), .B(n_537), .Y(n_731) );
INVx5_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g584 ( .A(n_517), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_517), .B(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_517), .B(n_579), .Y(n_591) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_517), .Y(n_593) );
OR2x2_ASAP7_75t_L g604 ( .A(n_517), .B(n_526), .Y(n_604) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_517), .B(n_595), .Y(n_609) );
AND2x2_ASAP7_75t_L g634 ( .A(n_517), .B(n_526), .Y(n_634) );
AND2x2_ASAP7_75t_L g654 ( .A(n_517), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g692 ( .A(n_517), .B(n_525), .Y(n_692) );
OR2x2_ASAP7_75t_L g695 ( .A(n_517), .B(n_681), .Y(n_695) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_526), .A2(n_639), .B(n_642), .C(n_648), .Y(n_638) );
INVx5_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_527), .B(n_537), .Y(n_569) );
AND2x2_ASAP7_75t_L g573 ( .A(n_527), .B(n_538), .Y(n_573) );
OR2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_537), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_SL g596 ( .A(n_537), .Y(n_596) );
OR2x2_ASAP7_75t_L g724 ( .A(n_537), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_564), .B(n_567), .C(n_576), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI31xp33_ASAP7_75t_L g649 ( .A1(n_547), .A2(n_650), .A3(n_652), .B(n_653), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_548), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_549), .B(n_580), .Y(n_586) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_550), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g606 ( .A(n_550), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_550), .B(n_581), .Y(n_611) );
AND2x2_ASAP7_75t_L g621 ( .A(n_550), .B(n_580), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_550), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_550), .B(n_598), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_550), .B(n_618), .Y(n_646) );
OR2x2_ASAP7_75t_L g665 ( .A(n_550), .B(n_552), .Y(n_665) );
OR2x2_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_550), .Y(n_714) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g614 ( .A(n_552), .B(n_581), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_552), .B(n_598), .Y(n_637) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g583 ( .A(n_554), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g674 ( .A(n_566), .B(n_598), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_566), .A2(n_580), .A3(n_618), .B1(n_677), .B2(n_678), .C1(n_679), .C2(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_SL g678 ( .A(n_568), .Y(n_678) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
OR2x2_ASAP7_75t_L g630 ( .A(n_569), .B(n_575), .Y(n_630) );
INVx1_ASAP7_75t_L g661 ( .A(n_569), .Y(n_661) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI32xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .A3(n_582), .B1(n_584), .B2(n_586), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI21xp33_ASAP7_75t_SL g616 ( .A1(n_579), .A2(n_594), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g631 ( .A(n_580), .Y(n_631) );
AND2x4_ASAP7_75t_L g628 ( .A(n_581), .B(n_598), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_581), .B(n_664), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_582), .A2(n_609), .A3(n_628), .B1(n_661), .B2(n_694), .C1(n_696), .C2(n_697), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_582), .A2(n_659), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_722) );
AND2x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g590 ( .A(n_585), .Y(n_590) );
OR2x2_ASAP7_75t_L g662 ( .A(n_585), .B(n_647), .Y(n_662) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .A3(n_592), .B(n_597), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_621), .B1(n_622), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g633 ( .A(n_590), .B(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_592), .A2(n_633), .B1(n_686), .B2(n_689), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g675 ( .A(n_595), .B(n_644), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_595), .B(n_634), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_596), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g709 ( .A(n_596), .B(n_647), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_597), .A2(n_692), .B1(n_705), .B2(n_708), .Y(n_704) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g613 ( .A(n_598), .Y(n_613) );
AND2x2_ASAP7_75t_L g696 ( .A(n_598), .B(n_618), .Y(n_696) );
OR2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_665), .Y(n_698) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_598), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_599), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_599), .B(n_644), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B(n_608), .C(n_620), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_612), .B2(n_615), .C(n_616), .Y(n_608) );
INVxp67_ASAP7_75t_L g720 ( .A(n_611), .Y(n_720) );
INVx1_ASAP7_75t_L g687 ( .A(n_612), .Y(n_687) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g651 ( .A(n_613), .B(n_618), .Y(n_651) );
INVx1_ASAP7_75t_L g668 ( .A(n_614), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_614), .B(n_641), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g683 ( .A(n_618), .Y(n_683) );
AND2x2_ASAP7_75t_L g689 ( .A(n_618), .B(n_644), .Y(n_689) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_SL g677 ( .A(n_625), .Y(n_677) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_628), .B(n_664), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_635), .C(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g725 ( .A(n_634), .Y(n_725) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g643 ( .A(n_637), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_641), .B(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_647), .Y(n_642) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_645), .A2(n_691), .B(n_693), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g702 ( .A(n_647), .Y(n_702) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B1(n_662), .B2(n_663), .C1(n_666), .C2(n_667), .Y(n_656) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g732 ( .A(n_663), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_664), .B(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_664), .A2(n_711), .B1(n_713), .B2(n_716), .Y(n_710) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_690), .C(n_703), .D(n_722), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_672), .B(n_702), .Y(n_712) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g679 ( .A(n_677), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_680), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .C(n_717), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_L g719 ( .A(n_715), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_729), .B(n_732), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g740 ( .A(n_733), .Y(n_740) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
XOR2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
endmodule