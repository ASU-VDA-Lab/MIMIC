module real_jpeg_24935_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_0),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_87),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

INVx8_ASAP7_75t_SL g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_28),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_8),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_12),
.A2(n_58),
.B1(n_75),
.B2(n_78),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_27),
.B1(n_63),
.B2(n_78),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_15),
.B(n_69),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_15),
.B(n_36),
.C(n_38),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_15),
.A2(n_28),
.B1(n_31),
.B2(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_15),
.B(n_41),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_15),
.B(n_49),
.C(n_53),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_15),
.A2(n_83),
.B(n_172),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_95),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_21),
.A2(n_22),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_25),
.B(n_44),
.C(n_59),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_31),
.B1(n_65),
.B2(n_66),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_28),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_28),
.B(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_31),
.A2(n_63),
.A3(n_66),
.B1(n_73),
.B2(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_33),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_33),
.A2(n_111),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_34),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_36),
.B(n_179),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_41),
.B(n_99),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_42),
.Y(n_110)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_46),
.A2(n_48),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_48),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_48),
.A2(n_54),
.B(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_48),
.B(n_71),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_50),
.B(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_55),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_57),
.B(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_70),
.B(n_76),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_113),
.B(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_71),
.B(n_199),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_80),
.B(n_95),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_93),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_93),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_82),
.A2(n_183),
.B1(n_185),
.B2(n_187),
.Y(n_182)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_86),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_89),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_117),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_126),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_124),
.A2(n_160),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_211),
.B(n_216),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_161),
.B(n_210),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_150),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_150),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_142),
.C(n_147),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_133),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_136),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_157),
.C(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_204),
.B(n_209),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_180),
.B(n_203),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_174),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_174),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_178),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B(n_202),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_188),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_196),
.B(n_201),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_193),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_208),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);


endmodule