module fake_aes_10120_n_31 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx3_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
NAND2xp33_ASAP7_75t_SL g12 ( .A(n_8), .B(n_4), .Y(n_12) );
CKINVDCx8_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_7), .B(n_5), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_1), .B(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_11), .B(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_19), .B(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AOI21xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_12), .B(n_17), .Y(n_26) );
OAI31xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_21), .A3(n_15), .B(n_14), .Y(n_27) );
NAND3x1_ASAP7_75t_L g28 ( .A(n_26), .B(n_27), .C(n_14), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_29), .B(n_10), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
endmodule