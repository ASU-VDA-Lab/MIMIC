module fake_netlist_6_2996_n_1747 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1747);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1747;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_57),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_79),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_40),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_48),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_78),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_37),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_45),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_107),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_35),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_58),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_112),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_116),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_98),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_96),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_91),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_71),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_7),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_67),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_64),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_28),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_141),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_36),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_63),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_92),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_26),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_29),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_19),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_99),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_90),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_146),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_47),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_42),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_147),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_52),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_5),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_75),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_125),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_41),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_148),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_113),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_95),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_87),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_30),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_83),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_123),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_21),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_32),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_55),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_81),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_106),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_6),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_11),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_138),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_68),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_118),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_46),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_121),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_41),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_47),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_82),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_132),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_126),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_10),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_4),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_101),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_37),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_28),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_89),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_129),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_127),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_94),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_32),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_111),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_163),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_168),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_225),
.Y(n_303)
);

BUFx6f_ASAP7_75t_SL g304 ( 
.A(n_241),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_171),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_171),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_153),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_171),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_171),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_169),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_160),
.B(n_0),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_171),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_154),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_171),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_220),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_171),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_223),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_155),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_165),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_157),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_157),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_170),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_172),
.B(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_159),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_156),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_165),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_206),
.B(n_159),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_233),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_173),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_161),
.B(n_1),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_183),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_254),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_156),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_161),
.B(n_1),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_191),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_184),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_177),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_177),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_186),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_191),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_189),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_190),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_193),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_257),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_224),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_224),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_239),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_201),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_205),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_239),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_207),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_208),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_273),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_178),
.B(n_4),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_214),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_228),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_229),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_152),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_152),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_258),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_178),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_307),
.B(n_200),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_336),
.B(n_185),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_309),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_200),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_236),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_180),
.Y(n_391)
);

NOR2x1_ASAP7_75t_L g392 ( 
.A(n_310),
.B(n_236),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_308),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_252),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_326),
.B(n_327),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_313),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_339),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_185),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_301),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_312),
.B(n_241),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_187),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_187),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_329),
.B(n_241),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_252),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_358),
.B(n_188),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_355),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_364),
.B(n_188),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_250),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_366),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_264),
.B1(n_298),
.B2(n_265),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_199),
.B1(n_263),
.B2(n_279),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_314),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_384),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_384),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_431),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_386),
.B(n_324),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_393),
.B(n_303),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_328),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_342),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_202),
.C(n_197),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_391),
.B(n_350),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_386),
.B(n_352),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_202),
.C(n_197),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_378),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_421),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_410),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_383),
.B(n_354),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_360),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_372),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_386),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_436),
.A2(n_264),
.B1(n_242),
.B2(n_213),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_366),
.Y(n_479)
);

AND3x2_ASAP7_75t_L g480 ( 
.A(n_394),
.B(n_300),
.C(n_250),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_431),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_391),
.B(n_365),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_391),
.A2(n_371),
.B1(n_340),
.B2(n_347),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_391),
.B(n_369),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_372),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_409),
.B(n_370),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_409),
.B(n_192),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_368),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_277),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_394),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_391),
.B(n_167),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_372),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_424),
.B(n_343),
.C(n_221),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_393),
.B(n_353),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_368),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_411),
.B(n_231),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_424),
.B(n_361),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_372),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_396),
.B(n_363),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_372),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_396),
.B(n_321),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_372),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_411),
.B(n_232),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_408),
.B(n_166),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_372),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_396),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_203),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_378),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_372),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_398),
.B(n_302),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_395),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_406),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_378),
.B(n_243),
.Y(n_528)
);

INVx6_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_408),
.B(n_419),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_408),
.B(n_203),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_378),
.Y(n_532)
);

AND2x2_ASAP7_75t_SL g533 ( 
.A(n_377),
.B(n_300),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_419),
.B(n_304),
.Y(n_534)
);

AND2x2_ASAP7_75t_SL g535 ( 
.A(n_377),
.B(n_167),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_419),
.B(n_304),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_406),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_378),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_395),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_419),
.A2(n_204),
.B1(n_198),
.B2(n_299),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_416),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_395),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_378),
.B(n_304),
.Y(n_543)
);

AO21x2_ASAP7_75t_L g544 ( 
.A1(n_377),
.A2(n_267),
.B(n_256),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_422),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_397),
.B(n_245),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_397),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_397),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_406),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_397),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_397),
.B(n_246),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_428),
.B(n_210),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_407),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

OAI21xp33_ASAP7_75t_L g559 ( 
.A1(n_428),
.A2(n_255),
.B(n_297),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_395),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_407),
.B(n_249),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_407),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_410),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_388),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_428),
.B(n_158),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_373),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g570 ( 
.A(n_379),
.B(n_167),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_398),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_373),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_427),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_388),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_373),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_428),
.B(n_259),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_413),
.B(n_417),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_435),
.B(n_266),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_374),
.B(n_269),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_427),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_374),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_435),
.B(n_210),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_374),
.B(n_271),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_471),
.B(n_311),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_520),
.B(n_435),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_517),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_530),
.B(n_392),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_530),
.B(n_392),
.Y(n_591)
);

NOR2xp67_ASAP7_75t_L g592 ( 
.A(n_455),
.B(n_413),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_457),
.Y(n_593)
);

NOR2x1p5_ASAP7_75t_L g594 ( 
.A(n_451),
.B(n_162),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_547),
.B(n_379),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_533),
.A2(n_392),
.B1(n_388),
.B2(n_390),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_449),
.B(n_450),
.Y(n_597)
);

NAND2x1_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_388),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_533),
.A2(n_388),
.B1(n_390),
.B2(n_385),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_569),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_530),
.B(n_379),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_547),
.B(n_385),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_569),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_437),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_530),
.B(n_385),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_437),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_440),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_528),
.A2(n_390),
.B(n_388),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_440),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_449),
.B(n_388),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_450),
.B(n_390),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_475),
.B(n_167),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_492),
.B(n_315),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_456),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_475),
.B(n_390),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_448),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_535),
.B(n_570),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_535),
.B(n_390),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_494),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_535),
.B(n_390),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_570),
.B(n_429),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_481),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_448),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_441),
.B(n_435),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_441),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_446),
.A2(n_320),
.B1(n_317),
.B2(n_287),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_453),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_453),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_451),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_494),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_452),
.A2(n_235),
.B(n_194),
.C(n_209),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_570),
.B(n_429),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_429),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_459),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_574),
.B(n_167),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_462),
.A2(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_459),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_461),
.A2(n_296),
.B1(n_219),
.B2(n_274),
.Y(n_642)
);

NOR3xp33_ASAP7_75t_L g643 ( 
.A(n_483),
.B(n_416),
.C(n_260),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_465),
.B(n_429),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_482),
.B(n_164),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_464),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_481),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_464),
.B(n_429),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_429),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_474),
.Y(n_652)
);

NAND2x1p5_ASAP7_75t_L g653 ( 
.A(n_574),
.B(n_215),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_488),
.B(n_489),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_567),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_485),
.B(n_174),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_518),
.B(n_176),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_511),
.B(n_175),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_556),
.A2(n_518),
.B1(n_460),
.B2(n_463),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_500),
.A2(n_215),
.B1(n_280),
.B2(n_267),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_430),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_496),
.B(n_430),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_496),
.B(n_430),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_507),
.B(n_430),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_574),
.B(n_427),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_430),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_582),
.B(n_521),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_572),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_582),
.B(n_430),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_521),
.B(n_531),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_575),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_575),
.Y(n_675)
);

O2A1O1Ixp5_ASAP7_75t_L g676 ( 
.A1(n_582),
.A2(n_400),
.B(n_375),
.C(n_376),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_550),
.B(n_427),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_582),
.B(n_375),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_521),
.A2(n_280),
.B1(n_217),
.B2(n_219),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_514),
.B(n_226),
.C(n_238),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_499),
.B(n_182),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_521),
.B(n_375),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_581),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_499),
.B(n_211),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_550),
.B(n_427),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_581),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

BUFx12f_ASAP7_75t_L g688 ( 
.A(n_571),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_522),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_376),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_495),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_531),
.B(n_376),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_532),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_532),
.B(n_217),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_499),
.B(n_212),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_467),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_538),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_495),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_538),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_444),
.B(n_176),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_546),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_550),
.B(n_427),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_497),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_568),
.A2(n_240),
.B1(n_283),
.B2(n_274),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_540),
.A2(n_240),
.B1(n_247),
.B2(n_256),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_380),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_SL g707 ( 
.A(n_504),
.B(n_254),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_497),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_501),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_571),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_460),
.B(n_413),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_556),
.A2(n_284),
.B1(n_247),
.B2(n_283),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_417),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_556),
.A2(n_284),
.B1(n_427),
.B2(n_434),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_501),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_509),
.B(n_216),
.Y(n_716)
);

BUFx6f_ASAP7_75t_SL g717 ( 
.A(n_556),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_467),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_529),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_545),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_508),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_546),
.B(n_380),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_529),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_463),
.B(n_417),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_549),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_454),
.B(n_222),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_503),
.B(n_276),
.C(n_227),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_508),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_553),
.B(n_380),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_534),
.A2(n_423),
.B1(n_420),
.B2(n_432),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_553),
.B(n_382),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_493),
.B(n_382),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_467),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_486),
.B(n_427),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_498),
.B(n_382),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_577),
.B(n_400),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_540),
.B(n_234),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_486),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_445),
.B(n_237),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_512),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_562),
.B(n_400),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_579),
.B(n_401),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_486),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_556),
.A2(n_434),
.B1(n_427),
.B2(n_195),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_420),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_583),
.B(n_401),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_487),
.B(n_401),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_512),
.Y(n_749)
);

BUFx5_ASAP7_75t_L g750 ( 
.A(n_563),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_487),
.B(n_434),
.Y(n_751)
);

AND2x4_ASAP7_75t_SL g752 ( 
.A(n_444),
.B(n_536),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_487),
.B(n_412),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_606),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_609),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_593),
.B(n_490),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_738),
.A2(n_559),
.B(n_443),
.C(n_476),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_601),
.A2(n_555),
.B(n_548),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_587),
.B(n_490),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_601),
.A2(n_506),
.B(n_490),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_597),
.B(n_506),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_607),
.A2(n_506),
.B(n_502),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_597),
.B(n_576),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_587),
.B(n_543),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_636),
.A2(n_564),
.B(n_563),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_595),
.B(n_578),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_659),
.A2(n_559),
.B(n_544),
.C(n_564),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_710),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_707),
.A2(n_525),
.B(n_541),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_696),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_615),
.B(n_545),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_602),
.B(n_438),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_592),
.B(n_438),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_705),
.A2(n_537),
.B(n_527),
.C(n_552),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_619),
.A2(n_527),
.B(n_537),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_627),
.B(n_438),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_628),
.A2(n_275),
.B(n_255),
.C(n_261),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_275),
.B1(n_265),
.B2(n_261),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_720),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_607),
.A2(n_561),
.B(n_502),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_669),
.B(n_445),
.Y(n_783)
);

BUFx8_ASAP7_75t_L g784 ( 
.A(n_720),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_627),
.B(n_491),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_587),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_552),
.B(n_557),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_609),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_616),
.Y(n_789)
);

OAI21xp33_ASAP7_75t_L g790 ( 
.A1(n_658),
.A2(n_278),
.B(n_290),
.Y(n_790)
);

AOI21x1_ASAP7_75t_L g791 ( 
.A1(n_666),
.A2(n_557),
.B(n_439),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_590),
.A2(n_561),
.B(n_502),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_618),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_590),
.A2(n_561),
.B(n_502),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_591),
.A2(n_561),
.B(n_526),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_621),
.A2(n_529),
.B1(n_491),
.B2(n_510),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_591),
.A2(n_598),
.B(n_665),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_628),
.A2(n_439),
.B(n_442),
.C(n_447),
.Y(n_798)
);

INVx6_ASAP7_75t_L g799 ( 
.A(n_688),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_635),
.A2(n_478),
.B(n_442),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_584),
.B(n_491),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_598),
.A2(n_526),
.B(n_510),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_586),
.B(n_510),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_668),
.A2(n_523),
.B(n_526),
.Y(n_804)
);

OAI21xp33_ASAP7_75t_L g805 ( 
.A1(n_716),
.A2(n_253),
.B(n_248),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_623),
.A2(n_529),
.B1(n_523),
.B2(n_539),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_523),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_672),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_672),
.A2(n_539),
.B1(n_468),
.B2(n_566),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_718),
.A2(n_539),
.B(n_445),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_632),
.B(n_480),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_672),
.B(n_445),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_625),
.B(n_254),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_608),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_736),
.B(n_447),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_608),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_676),
.A2(n_469),
.B(n_458),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_589),
.B(n_458),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_603),
.B(n_466),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_604),
.B(n_466),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_647),
.B(n_469),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

AOI21x1_ASAP7_75t_L g823 ( 
.A1(n_666),
.A2(n_478),
.B(n_484),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_585),
.B(n_470),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_588),
.B(n_470),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_657),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_620),
.B(n_477),
.Y(n_827)
);

OAI321xp33_ASAP7_75t_L g828 ( 
.A1(n_642),
.A2(n_213),
.A3(n_194),
.B1(n_209),
.B2(n_218),
.C(n_230),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_622),
.B(n_420),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_718),
.A2(n_551),
.B(n_445),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_633),
.B(n_477),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_718),
.A2(n_513),
.B(n_473),
.Y(n_832)
);

INVx11_ASAP7_75t_L g833 ( 
.A(n_688),
.Y(n_833)
);

BUFx4f_ASAP7_75t_L g834 ( 
.A(n_657),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_671),
.A2(n_513),
.B(n_473),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_618),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_637),
.A2(n_179),
.B(n_230),
.C(n_235),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_SL g838 ( 
.A1(n_710),
.A2(n_285),
.B1(n_262),
.B2(n_289),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_681),
.B(n_423),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_651),
.B(n_484),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_650),
.B(n_473),
.Y(n_841)
);

INVx11_ASAP7_75t_L g842 ( 
.A(n_594),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_742),
.A2(n_747),
.B(n_743),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_612),
.A2(n_515),
.B(n_473),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_752),
.B(n_179),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_650),
.B(n_473),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_613),
.A2(n_542),
.B(n_513),
.Y(n_847)
);

AO21x1_ASAP7_75t_L g848 ( 
.A1(n_653),
.A2(n_218),
.B(n_242),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_614),
.A2(n_244),
.B(n_268),
.C(n_291),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_670),
.B(n_513),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_674),
.B(n_513),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_686),
.B(n_515),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_713),
.A2(n_580),
.B(n_573),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_617),
.A2(n_551),
.B(n_515),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_684),
.B(n_515),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_626),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_626),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_753),
.A2(n_678),
.B(n_682),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_752),
.B(n_244),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_690),
.A2(n_551),
.B(n_515),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_611),
.B(n_542),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_630),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_735),
.A2(n_412),
.B(n_415),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_560),
.B(n_542),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_744),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_630),
.B(n_542),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_631),
.B(n_542),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_631),
.B(n_551),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_629),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_638),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_638),
.B(n_641),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_744),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_746),
.A2(n_580),
.B(n_573),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_641),
.B(n_551),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_735),
.A2(n_412),
.B(n_415),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_727),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_746),
.A2(n_580),
.B(n_573),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_650),
.B(n_560),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_646),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_646),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_652),
.B(n_560),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_706),
.A2(n_560),
.B(n_558),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_652),
.B(n_560),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_653),
.A2(n_268),
.B(n_291),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_614),
.A2(n_294),
.B(n_297),
.C(n_432),
.Y(n_885)
);

CKINVDCx10_ASAP7_75t_R g886 ( 
.A(n_717),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_695),
.B(n_270),
.C(n_281),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_748),
.A2(n_558),
.B(n_554),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_644),
.A2(n_558),
.B(n_554),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_645),
.A2(n_286),
.B(n_288),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_662),
.B(n_565),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_700),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_700),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_SL g894 ( 
.A(n_717),
.B(n_294),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_704),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_654),
.A2(n_558),
.B(n_554),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_610),
.A2(n_558),
.B(n_554),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_662),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_673),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_599),
.A2(n_565),
.B1(n_423),
.B2(n_432),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_673),
.B(n_565),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_648),
.A2(n_558),
.B(n_554),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_655),
.B(n_414),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_675),
.B(n_433),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_675),
.B(n_433),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_656),
.A2(n_415),
.B(n_426),
.C(n_414),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_683),
.B(n_433),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_683),
.B(n_433),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_751),
.A2(n_554),
.B(n_524),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_719),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_751),
.A2(n_737),
.B(n_639),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_639),
.A2(n_524),
.B(n_519),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_677),
.A2(n_524),
.B(n_519),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_667),
.A2(n_426),
.B1(n_415),
.B2(n_414),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_750),
.B(n_524),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_677),
.A2(n_702),
.B(n_685),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_687),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_712),
.A2(n_414),
.B1(n_426),
.B2(n_415),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_685),
.A2(n_702),
.B(n_653),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_649),
.A2(n_524),
.B(n_519),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_689),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_734),
.A2(n_524),
.B(n_519),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_600),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_711),
.B(n_426),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_426),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_739),
.A2(n_519),
.B(n_399),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_634),
.A2(n_434),
.B(n_519),
.C(n_12),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_693),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_600),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_605),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_697),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_680),
.B(n_104),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_SL g933 ( 
.A1(n_661),
.A2(n_8),
.B(n_9),
.C(n_12),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_719),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_699),
.B(n_434),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_701),
.Y(n_936)
);

CKINVDCx6p67_ASAP7_75t_R g937 ( 
.A(n_717),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_750),
.B(n_434),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_596),
.A2(n_663),
.B(n_664),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_719),
.A2(n_399),
.B(n_434),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_728),
.B(n_105),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_770),
.B(n_643),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_824),
.B(n_839),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_773),
.B(n_640),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_799),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_754),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_756),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_781),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_833),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_834),
.B(n_731),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_834),
.B(n_750),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_789),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_764),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_791),
.A2(n_605),
.B(n_722),
.Y(n_954)
);

AO22x1_ASAP7_75t_L g955 ( 
.A1(n_773),
.A2(n_726),
.B1(n_724),
.B2(n_723),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_788),
.Y(n_956)
);

OR2x6_ASAP7_75t_SL g957 ( 
.A(n_887),
.B(n_732),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_893),
.Y(n_958)
);

CKINVDCx8_ASAP7_75t_R g959 ( 
.A(n_886),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_758),
.A2(n_660),
.B(n_679),
.C(n_730),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_784),
.Y(n_961)
);

OA22x2_ASAP7_75t_L g962 ( 
.A1(n_826),
.A2(n_691),
.B1(n_698),
.B2(n_703),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_824),
.B(n_750),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_814),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_797),
.A2(n_723),
.B(n_714),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_843),
.A2(n_723),
.B(n_749),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_793),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_855),
.A2(n_694),
.B(n_740),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_786),
.A2(n_740),
.B1(n_694),
.B2(n_750),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_772),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_842),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_783),
.A2(n_709),
.B(n_749),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_876),
.B(n_715),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_892),
.B(n_750),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_757),
.A2(n_745),
.B1(n_709),
.B2(n_741),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_869),
.A2(n_691),
.B1(n_698),
.B2(n_703),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_816),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_845),
.A2(n_750),
.B1(n_741),
.B2(n_729),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_768),
.B(n_729),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_784),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_765),
.A2(n_721),
.B(n_715),
.C(n_708),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_779),
.A2(n_721),
.B(n_708),
.C(n_20),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_865),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_434),
.B1(n_399),
.B2(n_149),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_813),
.B(n_434),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_858),
.A2(n_399),
.B(n_434),
.Y(n_987)
);

INVx6_ASAP7_75t_L g988 ( 
.A(n_799),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_939),
.A2(n_399),
.B(n_145),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_845),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_990)
);

BUFx8_ASAP7_75t_SL g991 ( 
.A(n_941),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_895),
.B(n_18),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_837),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_837),
.A2(n_790),
.B(n_890),
.C(n_805),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_872),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_821),
.B(n_23),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_921),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_836),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_822),
.A2(n_399),
.B1(n_143),
.B2(n_128),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_828),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_859),
.B(n_25),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_872),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_859),
.B(n_31),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_771),
.B(n_31),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_927),
.A2(n_33),
.B(n_38),
.C(n_39),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_766),
.A2(n_399),
.B(n_56),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_921),
.B(n_399),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_911),
.A2(n_399),
.B(n_59),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_755),
.Y(n_1010)
);

OA21x2_ASAP7_75t_L g1011 ( 
.A1(n_853),
.A2(n_399),
.B(n_124),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_821),
.B(n_33),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_825),
.B(n_38),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_825),
.B(n_39),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_811),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_766),
.A2(n_40),
.B(n_43),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_759),
.A2(n_794),
.B(n_792),
.Y(n_1017)
);

OA21x2_ASAP7_75t_L g1018 ( 
.A1(n_873),
.A2(n_399),
.B(n_69),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_829),
.B(n_44),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_829),
.B(n_44),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_856),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_917),
.B(n_49),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_755),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_870),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_808),
.B(n_70),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_762),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_755),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_838),
.B(n_50),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_880),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_774),
.A2(n_84),
.B(n_108),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_928),
.B(n_52),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_871),
.A2(n_62),
.B(n_86),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_906),
.A2(n_97),
.B(n_119),
.C(n_53),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_919),
.A2(n_53),
.B(n_54),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_799),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_830),
.A2(n_54),
.B(n_832),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_811),
.B(n_941),
.C(n_932),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_755),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_763),
.A2(n_782),
.B(n_761),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_809),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_857),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_769),
.A2(n_877),
.B(n_916),
.C(n_780),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_772),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_910),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_937),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_SL g1046 ( 
.A(n_927),
.B(n_760),
.C(n_936),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_931),
.B(n_780),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_760),
.A2(n_899),
.B1(n_815),
.B2(n_812),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_808),
.B(n_894),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_932),
.B(n_862),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_933),
.A2(n_849),
.B(n_885),
.C(n_827),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_879),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_778),
.B(n_785),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_775),
.A2(n_810),
.B(n_767),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_SL g1055 ( 
.A1(n_841),
.A2(n_878),
.B(n_846),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_807),
.A2(n_878),
.B(n_846),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_902),
.A2(n_920),
.B(n_777),
.C(n_817),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_903),
.B(n_898),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_848),
.B(n_884),
.C(n_906),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_923),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_820),
.B(n_831),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_795),
.A2(n_776),
.B(n_798),
.C(n_903),
.Y(n_1062)
);

AND2x2_ASAP7_75t_SL g1063 ( 
.A(n_861),
.B(n_840),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_910),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_812),
.B(n_910),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_850),
.A2(n_852),
.B1(n_851),
.B2(n_841),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_910),
.B(n_934),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_929),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_930),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_818),
.B(n_819),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_934),
.B(n_925),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_801),
.B(n_803),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_891),
.B(n_901),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_900),
.B(n_868),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_904),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_934),
.Y(n_1076)
);

AND2x6_ASAP7_75t_L g1077 ( 
.A(n_934),
.B(n_883),
.Y(n_1077)
);

AO32x1_ASAP7_75t_L g1078 ( 
.A1(n_914),
.A2(n_796),
.A3(n_806),
.B1(n_933),
.B2(n_875),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_924),
.B(n_874),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_866),
.B(n_867),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_881),
.B(n_907),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_860),
.B(n_864),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_787),
.B(n_800),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_SL g1084 ( 
.A1(n_935),
.A2(n_918),
.B1(n_908),
.B2(n_905),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_844),
.B(n_854),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_863),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_918),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_847),
.A2(n_835),
.B(n_804),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_944),
.A2(n_938),
.B1(n_915),
.B2(n_802),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_948),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_968),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_952),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_943),
.A2(n_882),
.B(n_938),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_954),
.A2(n_966),
.B(n_1088),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1085),
.A2(n_823),
.B(n_897),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_998),
.B(n_1037),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1015),
.B(n_915),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_945),
.B(n_913),
.Y(n_1099)
);

BUFx10_ASAP7_75t_L g1100 ( 
.A(n_988),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_SL g1101 ( 
.A(n_1035),
.B(n_909),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_946),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1054),
.A2(n_889),
.B(n_896),
.Y(n_1103)
);

CKINVDCx11_ASAP7_75t_R g1104 ( 
.A(n_959),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_988),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_965),
.A2(n_888),
.B(n_922),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_972),
.B(n_926),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_1062),
.A2(n_912),
.A3(n_940),
.B(n_1016),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_953),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_962),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_944),
.B(n_1015),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1026),
.B(n_968),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1056),
.A2(n_973),
.B(n_1082),
.Y(n_1113)
);

AO21x1_ASAP7_75t_L g1114 ( 
.A1(n_995),
.A2(n_1034),
.B(n_1009),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1074),
.A2(n_1053),
.B(n_960),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_963),
.A2(n_1057),
.B(n_1061),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_1066),
.A2(n_985),
.A3(n_989),
.B(n_1036),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_SL g1118 ( 
.A1(n_1050),
.A2(n_1025),
.B(n_950),
.C(n_951),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_975),
.B(n_958),
.Y(n_1119)
);

BUFx2_ASAP7_75t_R g1120 ( 
.A(n_949),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1002),
.A2(n_1004),
.B1(n_1005),
.B2(n_1040),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1026),
.B(n_1053),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_974),
.B(n_980),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_962),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_SL g1125 ( 
.A(n_1002),
.B(n_1004),
.C(n_992),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_987),
.A2(n_1086),
.B(n_1071),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1048),
.A2(n_1007),
.B(n_1073),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1083),
.A2(n_1070),
.B(n_1080),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_976),
.A2(n_1081),
.A3(n_982),
.B(n_980),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_964),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1081),
.A2(n_1072),
.B(n_1079),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1084),
.A2(n_970),
.B(n_1063),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_978),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1005),
.A2(n_1014),
.B(n_1001),
.C(n_997),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_984),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1063),
.A2(n_1055),
.B(n_971),
.Y(n_1136)
);

AO32x2_ASAP7_75t_L g1137 ( 
.A1(n_977),
.A2(n_990),
.A3(n_1078),
.B1(n_1046),
.B2(n_1000),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1028),
.B(n_974),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_955),
.A2(n_1018),
.B(n_1011),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1012),
.A2(n_1078),
.A3(n_1047),
.B(n_1075),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_971),
.A2(n_1078),
.B(n_1018),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1022),
.A2(n_1031),
.A3(n_1030),
.B(n_1029),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_993),
.B(n_996),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1033),
.A2(n_1046),
.B(n_979),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1049),
.A2(n_1059),
.B(n_1008),
.C(n_1019),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1024),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1051),
.A2(n_986),
.B(n_1059),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1020),
.A2(n_1060),
.A3(n_1021),
.B(n_947),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_956),
.A2(n_1052),
.A3(n_967),
.B(n_999),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_993),
.B(n_1003),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1011),
.A2(n_1032),
.B(n_1043),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1065),
.A2(n_983),
.B(n_1033),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1087),
.B(n_1058),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_1069),
.B(n_1065),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1044),
.A2(n_1064),
.B(n_1006),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_994),
.A2(n_958),
.B(n_1068),
.C(n_996),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1043),
.A2(n_1027),
.B(n_1068),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1027),
.A2(n_1064),
.B(n_1044),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1003),
.B(n_957),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_981),
.A2(n_1045),
.B1(n_1023),
.B2(n_991),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1010),
.A2(n_1038),
.B(n_1023),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1076),
.A2(n_1077),
.A3(n_1067),
.B(n_1010),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1077),
.A2(n_1010),
.A3(n_1038),
.B(n_942),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1038),
.A2(n_945),
.B(n_1077),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1038),
.A2(n_1077),
.B(n_988),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_961),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_962),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1042),
.A2(n_1009),
.B(n_1088),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1035),
.Y(n_1169)
);

O2A1O1Ixp5_ASAP7_75t_L g1170 ( 
.A1(n_969),
.A2(n_593),
.B(n_944),
.C(n_1013),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_954),
.A2(n_1017),
.B(n_1039),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1015),
.B(n_834),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_943),
.A2(n_593),
.B1(n_944),
.B2(n_1087),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_944),
.A2(n_593),
.B1(n_425),
.B2(n_394),
.C(n_738),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_L g1177 ( 
.A(n_944),
.B(n_593),
.C(n_707),
.Y(n_1177)
);

INVxp67_ASAP7_75t_SL g1178 ( 
.A(n_968),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_948),
.B(n_468),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_948),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_954),
.A2(n_1017),
.B(n_1039),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_962),
.Y(n_1182)
);

AO32x2_ASAP7_75t_L g1183 ( 
.A1(n_977),
.A2(n_990),
.A3(n_659),
.B1(n_1048),
.B2(n_1066),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_943),
.B(n_593),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_948),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_945),
.B(n_1023),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_948),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_943),
.B(n_593),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1010),
.Y(n_1189)
);

AO32x2_ASAP7_75t_L g1190 ( 
.A1(n_977),
.A2(n_990),
.A3(n_659),
.B1(n_1048),
.B2(n_1066),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_834),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_954),
.A2(n_1017),
.B(n_1039),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_943),
.A2(n_593),
.B1(n_944),
.B2(n_1087),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_946),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_946),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1198)
);

CKINVDCx11_ASAP7_75t_R g1199 ( 
.A(n_959),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_955),
.A2(n_1082),
.B(n_1054),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_943),
.A2(n_593),
.B(n_944),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_1023),
.B(n_770),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_948),
.B(n_468),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1015),
.B(n_834),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1010),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_998),
.B(n_1037),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_944),
.A2(n_593),
.B1(n_585),
.B2(n_1037),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_944),
.A2(n_593),
.B1(n_1037),
.B2(n_738),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_948),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_943),
.B(n_593),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_SL g1214 ( 
.A(n_1050),
.B(n_951),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1042),
.A2(n_758),
.B(n_593),
.C(n_1050),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_943),
.B(n_593),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_998),
.B(n_1037),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_944),
.B(n_593),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_944),
.A2(n_593),
.B(n_585),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_969),
.A2(n_1042),
.A3(n_1017),
.B(n_1039),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_998),
.B(n_1037),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_962),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_954),
.A2(n_1017),
.B(n_1039),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_943),
.B(n_593),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1035),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1035),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_SL g1228 ( 
.A(n_952),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1054),
.A2(n_593),
.B(n_843),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1076),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_943),
.A2(n_593),
.B(n_944),
.Y(n_1231)
);

INVx6_ASAP7_75t_L g1232 ( 
.A(n_1100),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1110),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1130),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1090),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1104),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1184),
.B(n_1188),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_SL g1238 ( 
.A(n_1100),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1125),
.A2(n_1219),
.B1(n_1231),
.B2(n_1204),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1133),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1180),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1199),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1121),
.A2(n_1193),
.B1(n_1174),
.B2(n_1111),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1115),
.A2(n_1216),
.B1(n_1213),
.B2(n_1225),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1114),
.A2(n_1138),
.B1(n_1168),
.B2(n_1218),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1168),
.A2(n_1209),
.B1(n_1218),
.B2(n_1222),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1187),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1097),
.A2(n_1222),
.B1(n_1209),
.B2(n_1132),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1133),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_1228),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1220),
.A2(n_1173),
.B1(n_1207),
.B2(n_1191),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1097),
.A2(n_1122),
.B1(n_1147),
.B2(n_1123),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1194),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1144),
.A2(n_1128),
.B1(n_1159),
.B2(n_1153),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1105),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1162),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1169),
.A2(n_1227),
.B1(n_1179),
.B2(n_1206),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1134),
.A2(n_1205),
.B(n_1229),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1228),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1162),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1144),
.A2(n_1197),
.B1(n_1131),
.B2(n_1146),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1169),
.A2(n_1227),
.B1(n_1185),
.B2(n_1212),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1214),
.A2(n_1227),
.B1(n_1169),
.B2(n_1135),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1102),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1119),
.A2(n_1156),
.B1(n_1098),
.B2(n_1092),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1226),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1093),
.A2(n_1112),
.B1(n_1160),
.B2(n_1166),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1143),
.B(n_1150),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1163),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1109),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1186),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1178),
.B(n_1146),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1149),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1167),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1162),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1120),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1170),
.B(n_1148),
.Y(n_1278)
);

BUFx2_ASAP7_75t_R g1279 ( 
.A(n_1230),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1182),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1182),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1089),
.A2(n_1107),
.B1(n_1164),
.B2(n_1157),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1223),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1189),
.Y(n_1284)
);

BUFx8_ASAP7_75t_L g1285 ( 
.A(n_1208),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1223),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1116),
.A2(n_1198),
.B1(n_1217),
.B2(n_1176),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1208),
.Y(n_1288)
);

BUFx4_ASAP7_75t_R g1289 ( 
.A(n_1183),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1094),
.B2(n_1136),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1183),
.A2(n_1190),
.B1(n_1152),
.B2(n_1154),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1230),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1183),
.A2(n_1190),
.B1(n_1127),
.B2(n_1101),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_1165),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1148),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1163),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1118),
.A2(n_1145),
.B1(n_1215),
.B2(n_1099),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1190),
.A2(n_1155),
.B1(n_1141),
.B2(n_1137),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1158),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1161),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1200),
.A2(n_1137),
.B1(n_1139),
.B2(n_1151),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1163),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1142),
.Y(n_1303)
);

INVx4_ASAP7_75t_SL g1304 ( 
.A(n_1142),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1137),
.A2(n_1126),
.B1(n_1113),
.B2(n_1095),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1091),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1108),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1103),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1108),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1140),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1096),
.A2(n_1106),
.B1(n_1181),
.B2(n_1192),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1091),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1140),
.B(n_1129),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1117),
.A2(n_1129),
.B1(n_1091),
.B2(n_1172),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1171),
.A2(n_1224),
.B1(n_1117),
.B2(n_1195),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1221),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1195),
.A2(n_1202),
.B1(n_1203),
.B2(n_1221),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1195),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1202),
.A2(n_593),
.B1(n_1210),
.B2(n_1220),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1203),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1221),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1130),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_593),
.B2(n_1219),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1228),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1228),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1130),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1110),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1228),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1110),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1162),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1130),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1104),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1189),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1130),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1110),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_593),
.B2(n_1219),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_L g1337 ( 
.A(n_1104),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1177),
.A2(n_593),
.B1(n_707),
.B2(n_585),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1130),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1110),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1189),
.Y(n_1341)
);

OAI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1175),
.A2(n_593),
.B(n_1220),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1210),
.A2(n_593),
.B1(n_1220),
.B2(n_707),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1180),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_593),
.B2(n_1219),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1130),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_593),
.B2(n_1219),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1104),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_593),
.B2(n_1219),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1104),
.Y(n_1350)
);

BUFx8_ASAP7_75t_L g1351 ( 
.A(n_1228),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1110),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1177),
.A2(n_593),
.B1(n_707),
.B2(n_585),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1090),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1211),
.A2(n_593),
.B1(n_1210),
.B2(n_1175),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1323),
.A2(n_1347),
.B1(n_1345),
.B2(n_1349),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1274),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1294),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1295),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1323),
.A2(n_1349),
.B1(n_1347),
.B2(n_1345),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1336),
.A2(n_1355),
.B1(n_1342),
.B2(n_1338),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1336),
.A2(n_1353),
.B1(n_1239),
.B2(n_1244),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1242),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1241),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1287),
.A2(n_1298),
.B(n_1313),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1302),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1316),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1278),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1270),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1312),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1245),
.B(n_1291),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1247),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1244),
.B(n_1253),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1234),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1294),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1311),
.A2(n_1315),
.B(n_1287),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1294),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1249),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1301),
.A2(n_1314),
.B(n_1319),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1321),
.A2(n_1266),
.B(n_1318),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1298),
.A2(n_1290),
.B(n_1293),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1322),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1232),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1308),
.A2(n_1290),
.B(n_1282),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1245),
.B(n_1291),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1311),
.A2(n_1315),
.B(n_1296),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1296),
.A2(n_1330),
.B(n_1257),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1273),
.A2(n_1339),
.B(n_1326),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1306),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1317),
.B(n_1306),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1331),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1317),
.B(n_1253),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1297),
.A2(n_1259),
.B(n_1343),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1232),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1334),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1237),
.B(n_1269),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1307),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1232),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1299),
.A2(n_1346),
.B(n_1283),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1304),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1344),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1239),
.A2(n_1289),
.B1(n_1243),
.B2(n_1320),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1293),
.A2(n_1262),
.B(n_1255),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1261),
.A2(n_1276),
.B(n_1262),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1243),
.A2(n_1255),
.B(n_1248),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1275),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1286),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1246),
.A2(n_1233),
.B(n_1352),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1303),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1265),
.A2(n_1271),
.B(n_1327),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1250),
.A2(n_1280),
.B(n_1329),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1307),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1246),
.A2(n_1280),
.B(n_1340),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1252),
.A2(n_1248),
.B1(n_1300),
.B2(n_1258),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1281),
.B(n_1340),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1327),
.B(n_1335),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1309),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1310),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1289),
.A2(n_1235),
.B1(n_1354),
.B2(n_1292),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1254),
.A2(n_1305),
.B(n_1268),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1341),
.B(n_1279),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1272),
.B(n_1333),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1272),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1285),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1251),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1251),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1260),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1325),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1260),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1325),
.A2(n_1328),
.B1(n_1351),
.B2(n_1337),
.Y(n_1434)
);

INVx4_ASAP7_75t_SL g1435 ( 
.A(n_1238),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1288),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1324),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1377),
.A2(n_1324),
.B(n_1351),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1420),
.B(n_1256),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1361),
.A2(n_1256),
.B(n_1236),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1419),
.B(n_1337),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1420),
.B(n_1277),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1361),
.A2(n_1350),
.B1(n_1325),
.B2(n_1328),
.Y(n_1443)
);

OAI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1407),
.A2(n_1267),
.B(n_1332),
.C(n_1348),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1356),
.A2(n_1328),
.B(n_1351),
.C(n_1267),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1419),
.B(n_1414),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1368),
.B(n_1364),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1421),
.B(n_1398),
.Y(n_1448)
);

AOI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1362),
.A2(n_1356),
.B(n_1360),
.C(n_1404),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1372),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1421),
.B(n_1403),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1426),
.B(n_1399),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1360),
.A2(n_1362),
.B1(n_1404),
.B2(n_1395),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1423),
.A2(n_1373),
.B1(n_1394),
.B2(n_1386),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1363),
.B(n_1428),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1375),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1386),
.A2(n_1395),
.B(n_1381),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1428),
.B(n_1436),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1376),
.A2(n_1373),
.B(n_1378),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_SL g1460 ( 
.A(n_1395),
.B(n_1390),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1416),
.A2(n_1423),
.B(n_1394),
.C(n_1437),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1429),
.A2(n_1431),
.B(n_1430),
.C(n_1433),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1382),
.B(n_1358),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1395),
.A2(n_1381),
.B1(n_1387),
.B2(n_1371),
.Y(n_1464)
);

AO32x2_ASAP7_75t_L g1465 ( 
.A1(n_1358),
.A2(n_1378),
.A3(n_1368),
.B1(n_1385),
.B2(n_1396),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1428),
.B(n_1436),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1379),
.Y(n_1467)
);

AO32x1_ASAP7_75t_L g1468 ( 
.A1(n_1366),
.A2(n_1367),
.A3(n_1370),
.B1(n_1374),
.B2(n_1391),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1371),
.A2(n_1387),
.B1(n_1381),
.B2(n_1376),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1429),
.B(n_1437),
.C(n_1430),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1417),
.B(n_1418),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1388),
.A2(n_1406),
.B(n_1389),
.Y(n_1472)
);

AO32x2_ASAP7_75t_L g1473 ( 
.A1(n_1385),
.A2(n_1400),
.A3(n_1396),
.B1(n_1369),
.B2(n_1381),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1405),
.A2(n_1406),
.B(n_1425),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1418),
.B(n_1380),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1392),
.B(n_1369),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1418),
.B(n_1380),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1392),
.B(n_1384),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1480)
);

AO32x2_ASAP7_75t_L g1481 ( 
.A1(n_1383),
.A2(n_1365),
.A3(n_1415),
.B1(n_1410),
.B2(n_1412),
.Y(n_1481)
);

AO32x1_ASAP7_75t_L g1482 ( 
.A1(n_1366),
.A2(n_1367),
.A3(n_1374),
.B1(n_1370),
.B2(n_1391),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1405),
.A2(n_1425),
.B(n_1413),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1408),
.B(n_1409),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1376),
.A2(n_1432),
.B1(n_1431),
.B2(n_1433),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1453),
.A2(n_1405),
.B1(n_1383),
.B2(n_1432),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1470),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1464),
.B(n_1401),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1475),
.B(n_1365),
.Y(n_1489)
);

AOI222xp33_ASAP7_75t_L g1490 ( 
.A1(n_1440),
.A2(n_1432),
.B1(n_1435),
.B2(n_1408),
.C1(n_1409),
.C2(n_1397),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1456),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1475),
.B(n_1391),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1470),
.B(n_1397),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1473),
.B(n_1383),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1481),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1453),
.B(n_1405),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1402),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1467),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1443),
.A2(n_1434),
.B(n_1427),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1468),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1447),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1473),
.B(n_1383),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1481),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1401),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1440),
.A2(n_1427),
.B1(n_1393),
.B2(n_1415),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1359),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_1357),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.B(n_1359),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1460),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1483),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1465),
.B(n_1411),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1446),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1477),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1455),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1493),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1515),
.B(n_1471),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1487),
.A2(n_1449),
.B1(n_1443),
.B2(n_1454),
.C(n_1512),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1501),
.B(n_1450),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1514),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1515),
.B(n_1474),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1497),
.B(n_1463),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1497),
.B(n_1513),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1488),
.B(n_1449),
.C(n_1461),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1510),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1463),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1484),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1491),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1493),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1510),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1499),
.B(n_1444),
.C(n_1469),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1509),
.B(n_1484),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1496),
.A2(n_1448),
.B1(n_1451),
.B2(n_1458),
.Y(n_1538)
);

INVx5_ASAP7_75t_SL g1539 ( 
.A(n_1497),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_SL g1540 ( 
.A(n_1499),
.B(n_1462),
.C(n_1516),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1492),
.B(n_1465),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1491),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1512),
.B(n_1452),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1496),
.B(n_1514),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

OAI211xp5_ASAP7_75t_L g1548 ( 
.A1(n_1486),
.A2(n_1445),
.B(n_1485),
.C(n_1459),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1466),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1534),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1531),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1547),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1519),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1530),
.B(n_1537),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1522),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1547),
.B(n_1495),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1547),
.B(n_1495),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1537),
.B(n_1495),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1527),
.B(n_1495),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.B(n_1541),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1533),
.B(n_1502),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1549),
.B(n_1521),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1532),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1522),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1480),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1519),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1489),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1546),
.B(n_1528),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1539),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1539),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1539),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1550),
.B(n_1539),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1559),
.B(n_1518),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1553),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1578),
.B(n_1518),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1575),
.A2(n_1526),
.B1(n_1520),
.B2(n_1496),
.Y(n_1588)
);

AND2x4_ASAP7_75t_SL g1589 ( 
.A(n_1552),
.B(n_1540),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1555),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1592)
);

INVx5_ASAP7_75t_L g1593 ( 
.A(n_1555),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

AOI33xp33_ASAP7_75t_L g1595 ( 
.A1(n_1568),
.A2(n_1538),
.A3(n_1486),
.B1(n_1505),
.B2(n_1489),
.B3(n_1577),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1579),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1539),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1566),
.B(n_1503),
.Y(n_1601)
);

NOR2x1p5_ASAP7_75t_SL g1602 ( 
.A(n_1561),
.B(n_1500),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1578),
.B(n_1526),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1572),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1570),
.B(n_1442),
.Y(n_1606)
);

OAI21xp33_ASAP7_75t_L g1607 ( 
.A1(n_1558),
.A2(n_1496),
.B(n_1548),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1557),
.B(n_1529),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1551),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1551),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1563),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1563),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1556),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1563),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1558),
.A2(n_1508),
.B1(n_1500),
.B2(n_1506),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1567),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1557),
.B(n_1529),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1605),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1618),
.B(n_1568),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1593),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1605),
.Y(n_1623)
);

NAND4xp25_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1576),
.C(n_1490),
.D(n_1505),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1606),
.B(n_1441),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1609),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1568),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1609),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1593),
.B(n_1560),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1603),
.B(n_1564),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1603),
.B(n_1441),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1566),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1610),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1579),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.B(n_1579),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1595),
.B(n_1523),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1590),
.Y(n_1639)
);

XNOR2xp5_ASAP7_75t_L g1640 ( 
.A(n_1589),
.B(n_1439),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1589),
.B(n_1544),
.Y(n_1641)
);

AOI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1607),
.A2(n_1615),
.B(n_1590),
.C(n_1597),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1569),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1607),
.B(n_1594),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1589),
.B(n_1544),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1593),
.A2(n_1490),
.B1(n_1489),
.B2(n_1438),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1585),
.B(n_1545),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1600),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1599),
.B(n_1569),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1593),
.B(n_1569),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1594),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1615),
.A2(n_1511),
.B(n_1560),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1581),
.B(n_1562),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1599),
.B(n_1571),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1639),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1635),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1644),
.A2(n_1580),
.B1(n_1598),
.B2(n_1582),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1648),
.B(n_1580),
.Y(n_1658)
);

OAI321xp33_ASAP7_75t_L g1659 ( 
.A1(n_1642),
.A2(n_1596),
.A3(n_1586),
.B1(n_1580),
.B2(n_1583),
.C(n_1582),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1640),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1648),
.B(n_1582),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1651),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_SL g1663 ( 
.A(n_1646),
.B(n_1583),
.C(n_1598),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1635),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1583),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1621),
.B(n_1581),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1643),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1640),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1631),
.B(n_1587),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1630),
.B(n_1587),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1627),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1627),
.B(n_1653),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1625),
.B(n_1584),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_R g1675 ( 
.A1(n_1643),
.A2(n_1592),
.B(n_1584),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1619),
.Y(n_1676)
);

AOI31xp33_ASAP7_75t_L g1677 ( 
.A1(n_1629),
.A2(n_1598),
.A3(n_1586),
.B(n_1596),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1644),
.B(n_1608),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1626),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1624),
.B(n_1584),
.Y(n_1680)
);

AOI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1659),
.A2(n_1644),
.B(n_1623),
.Y(n_1681)
);

OAI31xp33_ASAP7_75t_L g1682 ( 
.A1(n_1660),
.A2(n_1629),
.A3(n_1641),
.B(n_1645),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1644),
.B1(n_1669),
.B2(n_1657),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1663),
.A2(n_1680),
.B1(n_1677),
.B2(n_1662),
.C(n_1655),
.Y(n_1684)
);

XNOR2x1_ASAP7_75t_L g1685 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1676),
.Y(n_1687)
);

OAI222xp33_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1629),
.B1(n_1643),
.B2(n_1650),
.C1(n_1653),
.C2(n_1637),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1662),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1667),
.Y(n_1690)
);

AOI211xp5_ASAP7_75t_L g1691 ( 
.A1(n_1665),
.A2(n_1652),
.B(n_1620),
.C(n_1623),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1666),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1656),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1666),
.B(n_1620),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1668),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1668),
.B(n_1650),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1658),
.B(n_1650),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1699)
);

AO22x2_ASAP7_75t_L g1700 ( 
.A1(n_1686),
.A2(n_1679),
.B1(n_1664),
.B2(n_1628),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1684),
.B(n_1682),
.C(n_1683),
.D(n_1681),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1698),
.Y(n_1702)
);

OAI222xp33_ASAP7_75t_L g1703 ( 
.A1(n_1692),
.A2(n_1658),
.B1(n_1661),
.B2(n_1690),
.C1(n_1687),
.C2(n_1695),
.Y(n_1703)
);

INVxp33_ASAP7_75t_L g1704 ( 
.A(n_1685),
.Y(n_1704)
);

XNOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1698),
.B(n_1697),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1697),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1696),
.Y(n_1707)
);

XNOR2xp5_ASAP7_75t_L g1708 ( 
.A(n_1691),
.B(n_1661),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1700),
.Y(n_1709)
);

NOR3xp33_ASAP7_75t_L g1710 ( 
.A(n_1701),
.B(n_1689),
.C(n_1688),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1704),
.B(n_1671),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1700),
.Y(n_1712)
);

NAND2x1_ASAP7_75t_L g1713 ( 
.A(n_1707),
.B(n_1696),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1707),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1708),
.A2(n_1674),
.B(n_1671),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1705),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1703),
.A2(n_1691),
.B(n_1694),
.C(n_1622),
.Y(n_1717)
);

NAND4xp25_ASAP7_75t_L g1718 ( 
.A(n_1710),
.B(n_1699),
.C(n_1702),
.D(n_1706),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1713),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1709),
.A2(n_1712),
.B1(n_1717),
.B2(n_1715),
.C(n_1711),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1716),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1714),
.A2(n_1622),
.B1(n_1632),
.B2(n_1637),
.C(n_1636),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1720),
.A2(n_1632),
.B(n_1628),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_SL g1724 ( 
.A(n_1721),
.B(n_1636),
.C(n_1633),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_SL g1725 ( 
.A(n_1719),
.B(n_1649),
.C(n_1654),
.D(n_1633),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1718),
.A2(n_1634),
.B1(n_1649),
.B2(n_1654),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1722),
.A2(n_1647),
.B1(n_1591),
.B2(n_1604),
.C(n_1617),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1634),
.B(n_1604),
.C(n_1617),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1724),
.B(n_1591),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_L g1730 ( 
.A(n_1725),
.B(n_1634),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1726),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1727),
.Y(n_1732)
);

OAI211xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1728),
.A2(n_1611),
.B(n_1617),
.C(n_1591),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1730),
.A2(n_1723),
.B(n_1602),
.C(n_1604),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1729),
.Y(n_1735)
);

AND3x1_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1614),
.C(n_1611),
.Y(n_1736)
);

AND3x4_ASAP7_75t_L g1737 ( 
.A(n_1736),
.B(n_1732),
.C(n_1733),
.Y(n_1737)
);

OAI22x1_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1735),
.B1(n_1734),
.B2(n_1584),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1738),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1739),
.A2(n_1574),
.B1(n_1612),
.B2(n_1614),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1614),
.B1(n_1611),
.B2(n_1612),
.Y(n_1741)
);

AND2x2_ASAP7_75t_SL g1742 ( 
.A(n_1741),
.B(n_1435),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1742),
.B(n_1602),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1612),
.B(n_1616),
.Y(n_1744)
);

XNOR2xp5_ASAP7_75t_L g1745 ( 
.A(n_1743),
.B(n_1435),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_R g1746 ( 
.A1(n_1745),
.A2(n_1744),
.B1(n_1435),
.B2(n_1601),
.C(n_1613),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1610),
.B(n_1616),
.C(n_1613),
.Y(n_1747)
);


endmodule