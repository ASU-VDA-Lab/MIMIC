module fake_netlist_6_4840_n_1107 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1107);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1107;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_698;
wire n_617;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_544;
wire n_468;
wire n_372;
wire n_923;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_645;
wire n_321;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_689;
wire n_345;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_861;
wire n_296;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_SL g280 ( 
.A(n_134),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_211),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_203),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_102),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_171),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_222),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_23),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_41),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_81),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_83),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_219),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_240),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_144),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_114),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_181),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_97),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_187),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_197),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_162),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_104),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_25),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_66),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_122),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_250),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_272),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_101),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_32),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_3),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_73),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_100),
.B(n_51),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_129),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_36),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_193),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_237),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_146),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_93),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_238),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_205),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_186),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_184),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_142),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_199),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_1),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_18),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_108),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_208),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_248),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_15),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_13),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_127),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_264),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_245),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_63),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_92),
.Y(n_354)
);

BUFx8_ASAP7_75t_SL g355 ( 
.A(n_226),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_22),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_221),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_77),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_16),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_30),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_161),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_262),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_133),
.Y(n_363)
);

BUFx8_ASAP7_75t_SL g364 ( 
.A(n_31),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_271),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_46),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_132),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_15),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_53),
.Y(n_369)
);

BUFx10_ASAP7_75t_L g370 ( 
.A(n_54),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_98),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_176),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_166),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_140),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_124),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_168),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_35),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_256),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_267),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_174),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_94),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_202),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_258),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_210),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_20),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_52),
.B(n_16),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_249),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_110),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_59),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_204),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_218),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_106),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_215),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_42),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_154),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_68),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_57),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_96),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_207),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_149),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_115),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_27),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_137),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_239),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_21),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_69),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_153),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_175),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_201),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_232),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_120),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_123),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_227),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_190),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_88),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_139),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_19),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_13),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_91),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_103),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_138),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_269),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_21),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_20),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_6),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_50),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_37),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_130),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_164),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_85),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_89),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_74),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_217),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_1),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_241),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_229),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_178),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_276),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_180),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_113),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_71),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_223),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_56),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_247),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_198),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_246),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_150),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_255),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_278),
.B(n_244),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_251),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_34),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_147),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_275),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_159),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_5),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_352),
.B(n_0),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_310),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_298),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_343),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_356),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_312),
.B(n_2),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_4),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_348),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_310),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_314),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_310),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_359),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

BUFx8_ASAP7_75t_L g471 ( 
.A(n_316),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_324),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_330),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_366),
.B(n_7),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_414),
.B(n_8),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_324),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_330),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_376),
.B(n_8),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

BUFx8_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_330),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_9),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_286),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_351),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_396),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_351),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_351),
.Y(n_489)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_304),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_10),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_285),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_315),
.B(n_11),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_282),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_290),
.Y(n_497)
);

OAI22x1_ASAP7_75t_SL g498 ( 
.A1(n_288),
.A2(n_12),
.B1(n_14),
.B2(n_17),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_296),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_386),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_300),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_306),
.A2(n_19),
.B(n_22),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_304),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_431),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_295),
.B(n_23),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_305),
.B(n_26),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_323),
.A2(n_28),
.B(n_29),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_308),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_342),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_349),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_355),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_318),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g517 ( 
.A(n_327),
.B(n_33),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_334),
.B(n_38),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_325),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_370),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_346),
.B(n_39),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_326),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_364),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_328),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_329),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_370),
.Y(n_527)
);

OA21x2_ASAP7_75t_L g528 ( 
.A1(n_331),
.A2(n_43),
.B(n_44),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_369),
.B(n_45),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_377),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_335),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_341),
.B(n_47),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_336),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_350),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_358),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_360),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_386),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_385),
.A2(n_442),
.B(n_451),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_407),
.B(n_58),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_362),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_367),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_375),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_381),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_399),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_397),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_400),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_399),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_339),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_411),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_283),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_284),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_368),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_496),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_494),
.B(n_280),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_552),
.B(n_554),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_462),
.A2(n_387),
.B1(n_384),
.B2(n_341),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_550),
.B(n_412),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_521),
.Y(n_562)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_509),
.A2(n_423),
.B(n_417),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_485),
.B(n_384),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_466),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_489),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_466),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_468),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_505),
.B(n_555),
.Y(n_570)
);

CKINVDCx6p67_ASAP7_75t_R g571 ( 
.A(n_527),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_468),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_517),
.B(n_309),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_496),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_474),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_507),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_474),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_527),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_428),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_513),
.B(n_394),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_492),
.B(n_281),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_527),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_432),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_492),
.B(n_287),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_544),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_463),
.B(n_337),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_553),
.B(n_289),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_544),
.B(n_433),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_548),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_497),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_464),
.B(n_292),
.C(n_291),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_500),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_293),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_500),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_479),
.B(n_353),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_506),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_506),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_506),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_548),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_530),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

NOR2x1_ASAP7_75t_L g623 ( 
.A(n_505),
.B(n_435),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_405),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_549),
.B(n_405),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

INVx8_ASAP7_75t_L g629 ( 
.A(n_490),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_535),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_472),
.B(n_438),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_548),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_542),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_547),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_484),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_609),
.B(n_514),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_624),
.B(n_519),
.Y(n_638)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_564),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_556),
.B(n_518),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_607),
.B(n_599),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_620),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_597),
.B(n_539),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_620),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_524),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_627),
.B(n_476),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_557),
.B(n_472),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_459),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_564),
.B(n_477),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_621),
.B(n_459),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_626),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_570),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_459),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_585),
.B(n_477),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_582),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_582),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_574),
.B(n_483),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_587),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_610),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_599),
.B(n_497),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_495),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_562),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_518),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_593),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_559),
.A2(n_495),
.B1(n_522),
.B2(n_475),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_577),
.B(n_522),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_568),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_577),
.B(n_532),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_598),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_619),
.B(n_499),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_603),
.B(n_458),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_561),
.B(n_471),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_588),
.B(n_511),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_616),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_559),
.B(n_471),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_603),
.B(n_458),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_614),
.C(n_592),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_616),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_618),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_584),
.B(n_525),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_595),
.B(n_481),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_619),
.B(n_499),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_526),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_590),
.B(n_481),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_583),
.B(n_531),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_566),
.B(n_533),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_566),
.B(n_534),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_614),
.B(n_475),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_618),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_580),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_632),
.B(n_508),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_563),
.B(n_361),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_567),
.B(n_573),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_586),
.B(n_502),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_586),
.B(n_409),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_592),
.B(n_418),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_623),
.B(n_294),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_612),
.B(n_538),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_594),
.B(n_297),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_502),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_602),
.B(n_299),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_629),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_560),
.B(n_543),
.Y(n_709)
);

OAI22xp33_ASAP7_75t_L g710 ( 
.A1(n_622),
.A2(n_467),
.B1(n_487),
.B2(n_501),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_565),
.B(n_543),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_596),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_569),
.B(n_546),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_572),
.B(n_546),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_633),
.B(n_301),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_575),
.B(n_551),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_596),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_639),
.B(n_576),
.Y(n_718)
);

O2A1O1Ixp5_ASAP7_75t_L g719 ( 
.A1(n_663),
.A2(n_529),
.B(n_551),
.C(n_444),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_636),
.B(n_567),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_704),
.A2(n_528),
.B(n_628),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_643),
.A2(n_528),
.B(n_628),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_646),
.B(n_573),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_675),
.A2(n_630),
.B(n_625),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_649),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_668),
.A2(n_439),
.B1(n_450),
.B2(n_453),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_671),
.A2(n_510),
.B(n_503),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_680),
.A2(n_630),
.B(n_631),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_701),
.B(n_702),
.C(n_679),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_638),
.B(n_576),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_699),
.A2(n_537),
.B(n_635),
.C(n_634),
.Y(n_732)
);

AOI21x1_ASAP7_75t_L g733 ( 
.A1(n_684),
.A2(n_591),
.B(n_578),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_658),
.A2(n_581),
.B(n_579),
.C(n_480),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_640),
.A2(n_581),
.B(n_579),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_640),
.A2(n_606),
.B(n_604),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_666),
.A2(n_611),
.B(n_608),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_681),
.A2(n_503),
.B1(n_545),
.B2(n_540),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_696),
.B(n_613),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_617),
.B(n_615),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_692),
.A2(n_605),
.B(n_600),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_648),
.A2(n_605),
.B(n_600),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_684),
.B(n_540),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_706),
.B(n_645),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_661),
.B(n_695),
.Y(n_745)
);

INVx6_ASAP7_75t_L g746 ( 
.A(n_708),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_698),
.A2(n_303),
.B(n_302),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_642),
.B(n_540),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_647),
.A2(n_461),
.B(n_465),
.C(n_460),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_670),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_652),
.A2(n_311),
.B(n_307),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_644),
.B(n_541),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_656),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_650),
.A2(n_473),
.B(n_469),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_676),
.A2(n_469),
.B(n_473),
.C(n_480),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_657),
.Y(n_756)
);

AOI222xp33_ASAP7_75t_L g757 ( 
.A1(n_710),
.A2(n_498),
.B1(n_685),
.B2(n_655),
.C1(n_637),
.C2(n_688),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_677),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_659),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_690),
.A2(n_691),
.B(n_654),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_641),
.A2(n_317),
.B(n_313),
.Y(n_761)
);

BUFx8_ASAP7_75t_L g762 ( 
.A(n_665),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_664),
.Y(n_763)
);

AOI21x1_ASAP7_75t_L g764 ( 
.A1(n_672),
.A2(n_470),
.B(n_320),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_660),
.B(n_541),
.Y(n_765)
);

CKINVDCx8_ASAP7_75t_R g766 ( 
.A(n_708),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_653),
.A2(n_402),
.B1(n_321),
.B2(n_322),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_697),
.B(n_319),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_687),
.B(n_332),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_674),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_689),
.B(n_629),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_705),
.B(n_629),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_700),
.B(n_333),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_690),
.A2(n_340),
.B(n_338),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_703),
.A2(n_408),
.B1(n_345),
.B2(n_456),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_682),
.Y(n_776)
);

O2A1O1Ixp5_ASAP7_75t_L g777 ( 
.A1(n_712),
.A2(n_545),
.B(n_541),
.C(n_455),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_691),
.A2(n_347),
.B(n_344),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_708),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_683),
.A2(n_678),
.B(n_667),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_707),
.B(n_354),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_651),
.A2(n_363),
.B(n_357),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_709),
.A2(n_371),
.B(n_365),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_694),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_711),
.A2(n_373),
.B(n_372),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_713),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_714),
.A2(n_416),
.B(n_454),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_662),
.B(n_374),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_716),
.A2(n_421),
.B(n_452),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_673),
.B(n_686),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_670),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_715),
.A2(n_712),
.B(n_717),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_721),
.A2(n_693),
.B(n_670),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_SL g794 ( 
.A(n_757),
.B(n_415),
.C(n_379),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_744),
.B(n_693),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_722),
.A2(n_693),
.B(n_61),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_753),
.Y(n_797)
);

AOI21x1_ASAP7_75t_L g798 ( 
.A1(n_733),
.A2(n_735),
.B(n_760),
.Y(n_798)
);

AO21x2_ASAP7_75t_L g799 ( 
.A1(n_728),
.A2(n_730),
.B(n_792),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_750),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_545),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_756),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_780),
.A2(n_60),
.B(n_62),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_725),
.B(n_378),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_736),
.A2(n_64),
.B(n_65),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_737),
.A2(n_67),
.B(n_70),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_740),
.A2(n_72),
.B(n_75),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_790),
.A2(n_449),
.B(n_448),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_723),
.B(n_380),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_719),
.A2(n_447),
.B(n_446),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_758),
.B(n_731),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_759),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_786),
.B(n_743),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_720),
.B(n_383),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_738),
.A2(n_445),
.B(n_443),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_718),
.B(n_388),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_739),
.B(n_390),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_750),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_724),
.B(n_391),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_729),
.B(n_392),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_750),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_727),
.A2(n_441),
.B(n_440),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_763),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_741),
.A2(n_76),
.B(n_78),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_770),
.Y(n_825)
);

INVx3_ASAP7_75t_SL g826 ( 
.A(n_746),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_771),
.B(n_395),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_776),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_732),
.B(n_398),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_784),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_781),
.A2(n_745),
.B1(n_768),
.B2(n_773),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_742),
.A2(n_437),
.B(n_434),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_734),
.B(n_403),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_791),
.B(n_745),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_748),
.A2(n_430),
.B(n_429),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_767),
.B(n_406),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_769),
.B(n_410),
.Y(n_837)
);

BUFx12f_ASAP7_75t_L g838 ( 
.A(n_762),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_754),
.A2(n_785),
.B(n_782),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_765),
.A2(n_422),
.B(n_413),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_797),
.Y(n_842)
);

AO21x2_ASAP7_75t_L g843 ( 
.A1(n_799),
.A2(n_764),
.B(n_789),
.Y(n_843)
);

AO21x2_ASAP7_75t_L g844 ( 
.A1(n_799),
.A2(n_761),
.B(n_752),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_826),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_834),
.Y(n_846)
);

NAND2x1p5_ASAP7_75t_L g847 ( 
.A(n_824),
.B(n_779),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_796),
.A2(n_777),
.B(n_749),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_812),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_800),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_811),
.B(n_773),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_806),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_813),
.A2(n_747),
.B(n_774),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_794),
.A2(n_829),
.B(n_813),
.C(n_836),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_798),
.A2(n_751),
.B(n_778),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_839),
.A2(n_788),
.B(n_787),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_804),
.B(n_772),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_807),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_803),
.A2(n_783),
.B(n_775),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_805),
.A2(n_755),
.B(n_80),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_841),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_841),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_802),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_838),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_817),
.B(n_766),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_800),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_823),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_793),
.A2(n_79),
.B(n_82),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_809),
.A2(n_84),
.B(n_86),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_825),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_810),
.A2(n_87),
.B(n_90),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_818),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_801),
.A2(n_795),
.B(n_819),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_810),
.A2(n_95),
.B(n_99),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_863),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_849),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_870),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_863),
.B(n_801),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_854),
.A2(n_809),
.B(n_814),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_867),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_867),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_842),
.Y(n_882)
);

AO21x1_ASAP7_75t_SL g883 ( 
.A1(n_869),
.A2(n_829),
.B(n_831),
.Y(n_883)
);

AO21x2_ASAP7_75t_L g884 ( 
.A1(n_853),
.A2(n_819),
.B(n_815),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_842),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_861),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_872),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_860),
.A2(n_833),
.B(n_820),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_851),
.B(n_814),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_873),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_860),
.A2(n_833),
.B(n_830),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_857),
.A2(n_828),
.B1(n_815),
.B2(n_837),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_872),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_845),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_850),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_861),
.B(n_841),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_873),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_866),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_846),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_865),
.B(n_816),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_862),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_868),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_868),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_884),
.A2(n_844),
.B(n_852),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_899),
.B(n_827),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_892),
.A2(n_874),
.B1(n_871),
.B2(n_822),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_882),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_900),
.A2(n_822),
.B1(n_861),
.B2(n_821),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_876),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_886),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_901),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_845),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_880),
.B(n_874),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_881),
.B(n_874),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_886),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_843),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_887),
.B(n_871),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_877),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_882),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_875),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_889),
.B(n_808),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_885),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_893),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_875),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_878),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_878),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_890),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_898),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_886),
.B(n_871),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_893),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_890),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_894),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_883),
.A2(n_843),
.B1(n_844),
.B2(n_859),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_897),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_895),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_886),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_926),
.B(n_927),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_924),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_894),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_918),
.B(n_926),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_928),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_879),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_912),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_924),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_931),
.B(n_884),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_911),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_928),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_932),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_917),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_910),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_906),
.A2(n_884),
.B1(n_843),
.B2(n_844),
.Y(n_952)
);

AND3x1_ASAP7_75t_L g953 ( 
.A(n_905),
.B(n_864),
.C(n_762),
.Y(n_953)
);

CKINVDCx14_ASAP7_75t_R g954 ( 
.A(n_933),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_922),
.B(n_896),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_930),
.Y(n_956)
);

BUFx2_ASAP7_75t_SL g957 ( 
.A(n_910),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_915),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_913),
.B(n_897),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_932),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_936),
.B(n_891),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_906),
.A2(n_864),
.B1(n_896),
.B2(n_859),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_909),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_929),
.B(n_896),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_915),
.B(n_902),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_919),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_923),
.B(n_891),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_907),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_907),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_933),
.A2(n_847),
.B1(n_903),
.B2(n_902),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_913),
.B(n_903),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_915),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_920),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_908),
.B(n_847),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_942),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_941),
.B(n_914),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_941),
.B(n_914),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_942),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_940),
.B(n_914),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_946),
.B(n_934),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_939),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_955),
.B(n_947),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_944),
.B(n_930),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_943),
.B(n_938),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_943),
.B(n_938),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_938),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_950),
.B(n_937),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_963),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_966),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_945),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_961),
.B(n_934),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_956),
.B(n_935),
.Y(n_992)
);

AND2x2_ASAP7_75t_SL g993 ( 
.A(n_962),
.B(n_930),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_948),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_959),
.B(n_935),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_956),
.B(n_904),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_956),
.B(n_920),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_959),
.B(n_921),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_951),
.B(n_921),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_971),
.B(n_967),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_971),
.B(n_925),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_949),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_949),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_988),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_1001),
.B(n_952),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_990),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_981),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_981),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_994),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_975),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_995),
.B(n_974),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1003),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1004),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_996),
.B(n_974),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_984),
.B(n_954),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_SL g1018 ( 
.A(n_991),
.B(n_957),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_975),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_978),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_978),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_996),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_1000),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_982),
.B(n_985),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_997),
.B(n_970),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1016),
.B(n_980),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_982),
.Y(n_1027)
);

AOI322xp5_ASAP7_75t_L g1028 ( 
.A1(n_1010),
.A2(n_993),
.A3(n_962),
.B1(n_952),
.B2(n_954),
.C1(n_987),
.C2(n_983),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1005),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1013),
.B(n_976),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_958),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1007),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1011),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1022),
.B(n_986),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1012),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1006),
.A2(n_986),
.B1(n_964),
.B2(n_999),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1014),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_1009),
.B(n_987),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1015),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1013),
.B(n_977),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1019),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1021),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_1023),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_1025),
.B(n_972),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1028),
.A2(n_993),
.B1(n_1017),
.B2(n_979),
.Y(n_1045)
);

OAI31xp33_ASAP7_75t_L g1046 ( 
.A1(n_1036),
.A2(n_1008),
.A3(n_1024),
.B(n_1002),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_1020),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_1043),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1026),
.B(n_1025),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1031),
.A2(n_953),
.B1(n_965),
.B2(n_998),
.Y(n_1050)
);

XOR2x2_ASAP7_75t_L g1051 ( 
.A(n_1027),
.B(n_992),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1030),
.B(n_968),
.Y(n_1052)
);

OAI31xp33_ASAP7_75t_L g1053 ( 
.A1(n_1029),
.A2(n_973),
.A3(n_969),
.B(n_847),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1031),
.A2(n_925),
.B1(n_960),
.B2(n_858),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1044),
.A2(n_852),
.B1(n_858),
.B2(n_888),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1044),
.A2(n_960),
.B1(n_852),
.B2(n_858),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1040),
.B(n_888),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_1033),
.A2(n_1039),
.B1(n_1037),
.B2(n_1032),
.C(n_1041),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1042),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1035),
.B(n_832),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1034),
.B(n_856),
.Y(n_1061)
);

OAI31xp33_ASAP7_75t_L g1062 ( 
.A1(n_1036),
.A2(n_840),
.A3(n_835),
.B(n_109),
.Y(n_1062)
);

AOI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_1045),
.A2(n_105),
.B1(n_107),
.B2(n_111),
.C(n_112),
.Y(n_1063)
);

AOI322xp5_ASAP7_75t_L g1064 ( 
.A1(n_1058),
.A2(n_116),
.A3(n_117),
.B1(n_118),
.B2(n_119),
.C1(n_121),
.C2(n_126),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1059),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1049),
.A2(n_1062),
.B1(n_1046),
.B2(n_1050),
.Y(n_1066)
);

AOI322xp5_ASAP7_75t_L g1067 ( 
.A1(n_1052),
.A2(n_128),
.A3(n_131),
.B1(n_135),
.B2(n_136),
.C1(n_141),
.C2(n_143),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_1057),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.C(n_152),
.Y(n_1068)
);

XOR2xp5_ASAP7_75t_L g1069 ( 
.A(n_1051),
.B(n_1054),
.Y(n_1069)
);

AO22x2_ASAP7_75t_L g1070 ( 
.A1(n_1048),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1053),
.A2(n_160),
.B1(n_163),
.B2(n_165),
.C(n_167),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1060),
.A2(n_1061),
.B1(n_1055),
.B2(n_1056),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1047),
.B(n_856),
.Y(n_1073)
);

OAI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1045),
.A2(n_848),
.B(n_855),
.C(n_172),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1045),
.A2(n_855),
.B(n_848),
.C(n_173),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_SL g1076 ( 
.A1(n_1045),
.A2(n_169),
.B(n_170),
.Y(n_1076)
);

AOI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1046),
.A2(n_177),
.B(n_179),
.C(n_182),
.Y(n_1077)
);

NAND4xp25_ASAP7_75t_L g1078 ( 
.A(n_1045),
.B(n_183),
.C(n_188),
.D(n_189),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1048),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1059),
.Y(n_1080)
);

NOR4xp25_ASAP7_75t_L g1081 ( 
.A(n_1078),
.B(n_192),
.C(n_195),
.D(n_200),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1079),
.B(n_206),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_1076),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_SL g1084 ( 
.A(n_1071),
.B(n_220),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1065),
.Y(n_1085)
);

NAND4xp25_ASAP7_75t_L g1086 ( 
.A(n_1084),
.B(n_1063),
.C(n_1077),
.D(n_1066),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1085),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_1081),
.B(n_1075),
.C(n_1074),
.Y(n_1088)
);

NOR2x1_ASAP7_75t_L g1089 ( 
.A(n_1082),
.B(n_1069),
.Y(n_1089)
);

NOR3x1_ASAP7_75t_L g1090 ( 
.A(n_1083),
.B(n_1080),
.C(n_1073),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_1090),
.B(n_1064),
.C(n_1067),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1089),
.B(n_1072),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1087),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1086),
.B(n_1068),
.C(n_1070),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.Y(n_1095)
);

NAND4xp75_ASAP7_75t_L g1096 ( 
.A(n_1092),
.B(n_1088),
.C(n_1070),
.D(n_228),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_1094),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1097),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1098),
.Y(n_1099)
);

AO22x2_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_1096),
.B1(n_1091),
.B2(n_230),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1100),
.A2(n_224),
.B(n_225),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_SL g1103 ( 
.A1(n_1102),
.A2(n_231),
.B(n_234),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1101),
.B(n_236),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_1104),
.A2(n_235),
.B(n_242),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_243),
.B(n_252),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1106),
.A2(n_259),
.B1(n_260),
.B2(n_266),
.Y(n_1107)
);


endmodule