module real_jpeg_26476_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_17),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_0),
.B(n_75),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_0),
.B(n_29),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_0),
.B(n_25),
.Y(n_332)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_17),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_2),
.B(n_57),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_2),
.B(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_29),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_2),
.B(n_25),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_2),
.B(n_269),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_103),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_75),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_33),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_4),
.B(n_29),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_5),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_17),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_5),
.B(n_75),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_5),
.B(n_57),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_5),
.B(n_33),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_57),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_29),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_8),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_9),
.B(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_9),
.B(n_57),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_33),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_9),
.B(n_29),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_9),
.B(n_25),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_9),
.B(n_251),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_11),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_75),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_57),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_33),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_11),
.B(n_29),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_11),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_11),
.B(n_251),
.Y(n_339)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_33),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_13),
.B(n_103),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_13),
.B(n_75),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_13),
.B(n_57),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_75),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_14),
.B(n_57),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_14),
.B(n_33),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_14),
.B(n_29),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_14),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_14),
.B(n_251),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_17),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.C(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_52),
.C(n_55),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_49),
.B1(n_55),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_39),
.B(n_118),
.Y(n_211)
);

INVx11_ASAP7_75t_L g251 ( 
.A(n_39),
.Y(n_251)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_43),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_43),
.B(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_44),
.B(n_124),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_44),
.B(n_247),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_53),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_72),
.C(n_74),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_55),
.A2(n_74),
.B1(n_79),
.B2(n_326),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_56),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_56),
.B(n_73),
.Y(n_259)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_81),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_60),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.C(n_77),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_61),
.B(n_370),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_62),
.B(n_81),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.CI(n_65),
.CON(n_62),
.SN(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_69),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_66),
.B(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_71),
.B(n_77),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_72),
.B(n_351),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_74),
.A2(n_297),
.B1(n_298),
.B2(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_74),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_SL g355 ( 
.A(n_74),
.B(n_297),
.C(n_324),
.Y(n_355)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_374),
.C(n_375),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_365),
.C(n_366),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_343),
.C(n_344),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_319),
.C(n_320),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_287),
.C(n_288),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_253),
.C(n_254),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_217),
.C(n_218),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_187),
.C(n_188),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_165),
.C(n_166),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_147),
.C(n_148),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_125),
.C(n_126),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.C(n_115),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_107),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_108),
.C(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_105),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_103),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_124),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.C(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_146),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.C(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_181),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_182),
.C(n_186),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_176),
.C(n_177),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_175),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_177),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.CI(n_180),
.CON(n_177),
.SN(n_177)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.CI(n_185),
.CON(n_182),
.SN(n_182)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_203),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_192),
.C(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_199),
.C(n_202),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_194),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.CI(n_197),
.CON(n_194),
.SN(n_194)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_210),
.C(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_206),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_209),
.B(n_242),
.C(n_243),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_213),
.C(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_238),
.B2(n_252),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_239),
.C(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_223),
.C(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_227),
.C(n_230),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_229),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_235),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_283),
.C(n_284),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.CI(n_250),
.CON(n_244),
.SN(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_285),
.B2(n_286),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_277),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_277),
.C(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_266),
.C(n_267),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_261),
.C(n_263),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_270),
.B1(n_271),
.B2(n_276),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_273),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_294),
.C(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_280),
.C(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_291),
.C(n_318),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_305),
.B2(n_318),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_300),
.C(n_301),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_301),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.CI(n_304),
.CON(n_301),
.SN(n_301)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_303),
.C(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_308),
.C(n_309),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_317),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_313),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_314),
.A2(n_315),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_340),
.C(n_341),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_342),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_333),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_333),
.C(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_328),
.C(n_329),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_329),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.CI(n_332),
.CON(n_329),
.SN(n_329)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_331),
.C(n_332),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_336),
.C(n_337),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_347),
.C(n_357),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_356),
.B2(n_357),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_354),
.C(n_355),
.Y(n_368)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_360),
.C(n_363),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_371),
.B1(n_372),
.B2(n_373),
.Y(n_366)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_367),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_369),
.C(n_373),
.Y(n_374)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);


endmodule