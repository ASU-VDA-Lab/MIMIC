module real_jpeg_11667_n_17 (n_248, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_248;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_213;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_56),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_11),
.B(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_12),
.B(n_53),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_26),
.C(n_40),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_12),
.B(n_61),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_12),
.A2(n_97),
.B(n_153),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_49),
.B(n_62),
.C(n_180),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_12),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_13),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_67),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_188)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_102),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.C(n_59),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_22),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_23),
.B(n_33),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_24),
.A2(n_28),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_24),
.A2(n_28),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_24),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_25),
.B(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_28),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_31),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_34),
.Y(n_224)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_36),
.B(n_142),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_37),
.A2(n_63),
.B(n_138),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_38),
.A2(n_45),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_38),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_38),
.B(n_140),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_38),
.A2(n_45),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_42),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_42),
.B(n_138),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_42),
.A2(n_150),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_45),
.B(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_46),
.B(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_57),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_47),
.A2(n_54),
.B(n_138),
.C(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_48),
.A2(n_55),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_49),
.A2(n_51),
.A3(n_54),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_64),
.B(n_65),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_64),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_60),
.A2(n_65),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_60),
.A2(n_88),
.B1(n_115),
.B2(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_66),
.Y(n_116)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_83),
.B2(n_84),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_82),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_94),
.B2(n_101),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_88),
.A2(n_116),
.B(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_92),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_98),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_97),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_97),
.A2(n_98),
.B1(n_123),
.B2(n_182),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_159),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_98),
.A2(n_167),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_107),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_103),
.B(n_105),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_107),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_117),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_235)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_117),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_122),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_231),
.A3(n_240),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_213),
.B(n_230),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_192),
.B(n_212),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_175),
.B(n_191),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_155),
.B(n_174),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_133),
.B(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_136),
.A2(n_139),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_163),
.B(n_173),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_161),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_172),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_186),
.C(n_190),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_194),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_205),
.B2(n_206),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_208),
.C(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_200),
.C(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_227),
.C(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_225),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_222),
.C(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_234),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_237),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule