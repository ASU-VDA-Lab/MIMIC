module fake_jpeg_26291_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_16),
.B1(n_15),
.B2(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_18),
.B1(n_11),
.B2(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_0),
.Y(n_24)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_33)
);

OR2x4_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_9),
.B(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_13),
.B1(n_26),
.B2(n_4),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.C(n_19),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_32),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_11),
.B1(n_13),
.B2(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_42),
.B1(n_33),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_1),
.B1(n_3),
.B2(n_8),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.C(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_36),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_47),
.C(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_51),
.C(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_53),
.Y(n_54)
);

NOR2xp67_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_30),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_57),
.C(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_1),
.B1(n_3),
.B2(n_50),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_55),
.C(n_58),
.Y(n_61)
);


endmodule