module fake_netlist_5_2166_n_1529 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1529);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1529;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_56),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_89),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_106),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_105),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_87),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_9),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_83),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_42),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_15),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_74),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_32),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_41),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_32),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_134),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_22),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_2),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_84),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_57),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_42),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_43),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_63),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_41),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_31),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_102),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_9),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_92),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_140),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_123),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_26),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_19),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_45),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_40),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_1),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_54),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_103),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_30),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_100),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_132),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_68),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_12),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_20),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_37),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_66),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_80),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_28),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_21),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_8),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_137),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_22),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_34),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_47),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_70),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_27),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_23),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_23),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_33),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_25),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_53),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_64),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_19),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_96),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_85),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_125),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_73),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_98),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_51),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_101),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_59),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_61),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_82),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_46),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_4),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_44),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_28),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_16),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_24),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_48),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_38),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_130),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_157),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_179),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_180),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_181),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_186),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_191),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_176),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_202),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_194),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_219),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_176),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_176),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_195),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_176),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_176),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_238),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_276),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_175),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_165),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_288),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_170),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_201),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_206),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_217),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_188),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_302),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_229),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_204),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_231),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_231),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_223),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_188),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_178),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_210),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_232),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_284),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_210),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_237),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_239),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_240),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_243),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_170),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_172),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_172),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_254),
.Y(n_375)
);

BUFx2_ASAP7_75t_SL g376 ( 
.A(n_211),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_294),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_214),
.B(n_187),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_364),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_310),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_254),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_330),
.B(n_211),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_331),
.B(n_167),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_235),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_299),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_319),
.A2(n_207),
.B1(n_248),
.B2(n_255),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_167),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

CKINVDCx8_ASAP7_75t_R g415 ( 
.A(n_361),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_235),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_352),
.A2(n_275),
.B1(n_258),
.B2(n_251),
.Y(n_423)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_313),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_351),
.B(n_355),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_306),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_340),
.B(n_306),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_307),
.A2(n_174),
.B1(n_303),
.B2(n_267),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_355),
.B(n_199),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_309),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_315),
.B(n_317),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_315),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_366),
.A2(n_174),
.B1(n_303),
.B2(n_267),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_154),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_324),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_318),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_318),
.B(n_154),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_320),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_320),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_314),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_436),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_316),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

CKINVDCx6p67_ASAP7_75t_R g447 ( 
.A(n_408),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_386),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_345),
.B1(n_343),
.B2(n_329),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_325),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_435),
.B(n_347),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_407),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_435),
.B(n_357),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_377),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_360),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_394),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_415),
.Y(n_464)
);

BUFx6f_ASAP7_75t_SL g465 ( 
.A(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_425),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_382),
.A2(n_299),
.B1(n_374),
.B2(n_372),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_406),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_367),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_424),
.B(n_365),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_416),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

INVx8_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_406),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_368),
.Y(n_480)
);

AO21x2_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_171),
.B(n_160),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_369),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_406),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_434),
.B(n_371),
.C(n_370),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_408),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_377),
.B(n_199),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_434),
.B(n_156),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_321),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_388),
.B(n_161),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_396),
.B(n_363),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_SL g501 ( 
.A(n_416),
.B(n_269),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_388),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_415),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_440),
.Y(n_506)
);

AND3x2_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_266),
.C(n_159),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_428),
.B(n_373),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_428),
.B(n_339),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_407),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_401),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_411),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_423),
.A2(n_333),
.B1(n_326),
.B2(n_353),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_440),
.B(n_274),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_378),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_382),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_389),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_378),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_423),
.B(n_356),
.C(n_375),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_380),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_415),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_409),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_383),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_383),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_387),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_392),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_392),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_390),
.A2(n_322),
.B(n_224),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_395),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_411),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_430),
.B(n_363),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_430),
.B(n_156),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_390),
.B(n_269),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_400),
.A2(n_271),
.B1(n_190),
.B2(n_183),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_398),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_430),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_382),
.A2(n_268),
.B1(n_236),
.B2(n_242),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_430),
.B(n_158),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_393),
.B(n_322),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_400),
.B(n_158),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_382),
.B(n_356),
.C(n_375),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_393),
.B(n_250),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_393),
.B(n_403),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_393),
.B(n_403),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_382),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_410),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_410),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_397),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_412),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_412),
.B(n_256),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_409),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_413),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_409),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_418),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_420),
.B(n_162),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_420),
.Y(n_574)
);

AND2x2_ASAP7_75t_SL g575 ( 
.A(n_397),
.B(n_215),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_414),
.B(n_337),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_422),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_414),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_460),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_574),
.B(n_419),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_455),
.B(n_162),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_575),
.B(n_274),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_476),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_419),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_575),
.B(n_421),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_493),
.A2(n_341),
.B1(n_155),
.B2(n_265),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_463),
.B(n_421),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_463),
.B(n_422),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_200),
.C(n_218),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_456),
.B(n_270),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_457),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_492),
.B(n_270),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_526),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_502),
.B(n_188),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_510),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_561),
.A2(n_252),
.B1(n_292),
.B2(n_260),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_466),
.B(n_418),
.Y(n_599)
);

OAI221xp5_ASAP7_75t_L g600 ( 
.A1(n_509),
.A2(n_297),
.B1(n_301),
.B2(n_216),
.C(n_212),
.Y(n_600)
);

AO221x1_ASAP7_75t_L g601 ( 
.A1(n_544),
.A2(n_274),
.B1(n_287),
.B2(n_177),
.C(n_304),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_561),
.A2(n_230),
.B(n_264),
.C(n_205),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_493),
.B(n_281),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_442),
.B(n_502),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_513),
.B(n_164),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_264),
.Y(n_606)
);

AND2x4_ASAP7_75t_SL g607 ( 
.A(n_494),
.B(n_184),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_189),
.C(n_197),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_466),
.B(n_418),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_470),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_468),
.B(n_418),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_468),
.B(n_384),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_471),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_513),
.B(n_358),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_469),
.B(n_384),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_445),
.B(n_164),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_469),
.B(n_384),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

BUFx8_ASAP7_75t_L g619 ( 
.A(n_465),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_477),
.B(n_391),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_483),
.B(n_391),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_391),
.Y(n_622)
);

NAND3x1_ASAP7_75t_L g623 ( 
.A(n_449),
.B(n_259),
.C(n_198),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_500),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_503),
.B(n_185),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_505),
.B(n_208),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_486),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_514),
.B(n_220),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_500),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_489),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_446),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_474),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_450),
.B(n_166),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_454),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_547),
.B(n_166),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_493),
.B(n_282),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_499),
.B(n_221),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_458),
.B(n_168),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_518),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_454),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_518),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_493),
.A2(n_289),
.B1(n_283),
.B2(n_285),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_527),
.B(n_257),
.C(n_182),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_577),
.B(n_169),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_474),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_552),
.A2(n_274),
.B1(n_287),
.B2(n_286),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_478),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_451),
.B(n_169),
.Y(n_649)
);

NAND2x1p5_ASAP7_75t_L g650 ( 
.A(n_540),
.B(n_234),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_576),
.B(n_358),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_493),
.B(n_249),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_493),
.B(n_262),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_461),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_453),
.B(n_173),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_452),
.A2(n_279),
.B1(n_300),
.B2(n_298),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_525),
.B(n_290),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_495),
.B(n_173),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_554),
.B(n_291),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_475),
.B(n_273),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_559),
.B(n_295),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_566),
.B(n_273),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_539),
.B(n_278),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_461),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_560),
.B(n_287),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_539),
.B(n_280),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_443),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_573),
.A2(n_359),
.B(n_280),
.C(n_279),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_496),
.B(n_287),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g672 ( 
.A(n_448),
.B(n_49),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_494),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_522),
.A2(n_287),
.B1(n_300),
.B2(n_296),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_548),
.B(n_241),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_462),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_563),
.B(n_572),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_551),
.A2(n_263),
.B(n_261),
.C(n_253),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_501),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_247),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_481),
.A2(n_246),
.B1(n_245),
.B2(n_244),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_538),
.B(n_233),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_541),
.B(n_227),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_499),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_539),
.B(n_213),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_209),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_478),
.B(n_203),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_462),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_540),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_545),
.B(n_196),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_549),
.B(n_193),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_501),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_521),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_481),
.B(n_192),
.Y(n_695)
);

O2A1O1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_520),
.A2(n_3),
.B(n_6),
.C(n_7),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_481),
.B(n_65),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_546),
.B(n_58),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_546),
.B(n_69),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_546),
.B(n_564),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_528),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_528),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_473),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_531),
.Y(n_704)
);

AOI221xp5_ASAP7_75t_L g705 ( 
.A1(n_542),
.A2(n_3),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_564),
.B(n_75),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_564),
.B(n_76),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_542),
.B(n_11),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_443),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_473),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_459),
.B(n_13),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_464),
.B(n_14),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_478),
.A2(n_556),
.B(n_567),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_567),
.B(n_86),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_497),
.A2(n_78),
.B(n_148),
.Y(n_715)
);

NAND2x1_ASAP7_75t_L g716 ( 
.A(n_567),
.B(n_52),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_459),
.B(n_17),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_534),
.B(n_90),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_464),
.B(n_18),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_504),
.B(n_18),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_535),
.B(n_93),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_535),
.B(n_50),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_L g723 ( 
.A(n_645),
.B(n_659),
.C(n_656),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_651),
.B(n_504),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_688),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_604),
.B(n_578),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_595),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_604),
.B(n_497),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_498),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_648),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_596),
.B(n_529),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_653),
.B(n_498),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_671),
.B(n_569),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_690),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_610),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_690),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_668),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_613),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_529),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_633),
.B(n_507),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_597),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_618),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_587),
.B(n_519),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_447),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_708),
.A2(n_452),
.B1(n_512),
.B2(n_465),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_663),
.A2(n_616),
.B1(n_634),
.B2(n_594),
.Y(n_748)
);

NAND2x1_ASAP7_75t_L g749 ( 
.A(n_648),
.B(n_487),
.Y(n_749)
);

AOI21x1_ASAP7_75t_L g750 ( 
.A1(n_582),
.A2(n_558),
.B(n_557),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_645),
.B(n_447),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_624),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_628),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_543),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_553),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_648),
.B(n_506),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_648),
.B(n_478),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_597),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_636),
.B(n_512),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_592),
.B(n_562),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_565),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_630),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_598),
.B(n_562),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_598),
.B(n_565),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_636),
.B(n_517),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_701),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_709),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_663),
.B(n_465),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_593),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_597),
.B(n_482),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_640),
.B(n_515),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_704),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_642),
.B(n_479),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_583),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_672),
.B(n_506),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_634),
.B(n_506),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_580),
.B(n_584),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_591),
.B(n_550),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_681),
.A2(n_511),
.B1(n_517),
.B2(n_516),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_615),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_617),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_620),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_585),
.B(n_588),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_627),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_679),
.B(n_693),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_621),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_716),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_700),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_589),
.B(n_490),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_605),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_622),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_608),
.B(n_467),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_605),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_619),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_677),
.B(n_695),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_684),
.B(n_568),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_703),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_619),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_659),
.B(n_520),
.C(n_511),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_608),
.B(n_488),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_581),
.Y(n_804)
);

BUFx5_ASAP7_75t_L g805 ( 
.A(n_720),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_673),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_710),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_627),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_649),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_649),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_647),
.A2(n_536),
.B1(n_484),
.B2(n_487),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_661),
.A2(n_444),
.B1(n_484),
.B2(n_487),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_607),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_632),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_712),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_656),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_627),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_661),
.A2(n_444),
.B1(n_484),
.B2(n_555),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_SL g819 ( 
.A(n_657),
.B(n_24),
.C(n_25),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_586),
.B(n_467),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_635),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_641),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_683),
.B(n_467),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_655),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_639),
.Y(n_825)
);

BUFx4f_ASAP7_75t_L g826 ( 
.A(n_638),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_582),
.B(n_444),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_698),
.B(n_467),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_665),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_SL g830 ( 
.A(n_600),
.B(n_705),
.C(n_708),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_676),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_683),
.A2(n_571),
.B(n_488),
.C(n_508),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_698),
.B(n_488),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_689),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_680),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_684),
.B(n_570),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_682),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_606),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_599),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_SL g840 ( 
.A1(n_692),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_609),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_611),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_714),
.B(n_488),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_686),
.B(n_691),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_670),
.A2(n_530),
.B(n_570),
.C(n_555),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_606),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_625),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_662),
.B(n_488),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_638),
.B(n_555),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_644),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_571),
.Y(n_851)
);

BUFx8_ASAP7_75t_L g852 ( 
.A(n_623),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_606),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_626),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_647),
.B(n_571),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_697),
.B(n_571),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_658),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_629),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_650),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_36),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_638),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_861)
);

BUFx4f_ASAP7_75t_L g862 ( 
.A(n_650),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_666),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_718),
.Y(n_864)
);

NOR2x2_ASAP7_75t_L g865 ( 
.A(n_590),
.B(n_40),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_660),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_696),
.A2(n_43),
.B(n_571),
.C(n_537),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_699),
.B(n_537),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_706),
.B(n_537),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_685),
.B(n_530),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_707),
.A2(n_530),
.B(n_523),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_719),
.B(n_523),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_652),
.Y(n_873)
);

NOR2x2_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_94),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_654),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_674),
.B(n_523),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_674),
.B(n_508),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_868),
.A2(n_713),
.B(n_603),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_723),
.B(n_678),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_748),
.A2(n_669),
.B(n_715),
.C(n_675),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_739),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_731),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_726),
.B(n_601),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_724),
.B(n_667),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_809),
.B(n_664),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_793),
.A2(n_602),
.B(n_687),
.C(n_643),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_793),
.B(n_717),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_761),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_796),
.B(n_722),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_830),
.A2(n_637),
.B(n_721),
.C(n_119),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_777),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_868),
.A2(n_508),
.B(n_524),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_770),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_869),
.A2(n_508),
.B(n_524),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_725),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_761),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_869),
.A2(n_524),
.B(n_118),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_796),
.A2(n_524),
.B(n_121),
.C(n_124),
.Y(n_898)
);

AOI22x1_ASAP7_75t_L g899 ( 
.A1(n_863),
.A2(n_112),
.B1(n_126),
.B2(n_145),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_810),
.A2(n_524),
.B1(n_146),
.B2(n_151),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_816),
.B(n_741),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_786),
.B(n_780),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_779),
.A2(n_823),
.B(n_856),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_805),
.B(n_837),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_856),
.A2(n_791),
.B(n_786),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_830),
.A2(n_745),
.B(n_835),
.C(n_788),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_798),
.B(n_835),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_798),
.B(n_847),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_766),
.B(n_854),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_799),
.B(n_838),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_759),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_732),
.B(n_804),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_731),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_871),
.A2(n_731),
.B(n_828),
.Y(n_914)
);

OR2x6_ASAP7_75t_SL g915 ( 
.A(n_768),
.B(n_801),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_731),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_727),
.B(n_813),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_866),
.B(n_734),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_825),
.B(n_758),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_858),
.B(n_857),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_747),
.B(n_746),
.C(n_840),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_805),
.B(n_862),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_728),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_729),
.B(n_776),
.Y(n_924)
);

INVx5_ASAP7_75t_L g925 ( 
.A(n_728),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_728),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_805),
.B(n_862),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_871),
.A2(n_833),
.B(n_828),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_758),
.B(n_859),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_850),
.A2(n_844),
.B(n_769),
.C(n_867),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_805),
.B(n_747),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_743),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_867),
.A2(n_781),
.B(n_755),
.C(n_754),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_729),
.B(n_783),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_833),
.A2(n_843),
.B(n_778),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_870),
.A2(n_875),
.B(n_873),
.C(n_860),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_797),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_742),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_736),
.B(n_738),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_799),
.B(n_838),
.Y(n_940)
);

CKINVDCx14_ASAP7_75t_R g941 ( 
.A(n_826),
.Y(n_941)
);

CKINVDCx11_ASAP7_75t_R g942 ( 
.A(n_846),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_787),
.B(n_846),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_805),
.B(n_754),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_775),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_805),
.A2(n_872),
.B1(n_859),
.B2(n_836),
.Y(n_946)
);

AO22x1_ASAP7_75t_L g947 ( 
.A1(n_852),
.A2(n_742),
.B1(n_815),
.B2(n_808),
.Y(n_947)
);

BUFx12f_ASAP7_75t_L g948 ( 
.A(n_846),
.Y(n_948)
);

AND3x1_ASAP7_75t_SL g949 ( 
.A(n_874),
.B(n_865),
.C(n_861),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_836),
.B(n_743),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_819),
.B(n_753),
.C(n_762),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_843),
.A2(n_757),
.B(n_851),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_784),
.B(n_785),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_853),
.A2(n_806),
.B1(n_817),
.B2(n_808),
.Y(n_954)
);

BUFx2_ASAP7_75t_SL g955 ( 
.A(n_743),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_817),
.B(n_808),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_849),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_792),
.A2(n_855),
.B(n_827),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_817),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_789),
.B(n_794),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_826),
.B(n_787),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_763),
.A2(n_765),
.B1(n_876),
.B2(n_755),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_827),
.A2(n_756),
.B(n_820),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_839),
.B(n_841),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_842),
.B(n_752),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_876),
.A2(n_763),
.B(n_765),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_740),
.B(n_744),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_SL g968 ( 
.A1(n_795),
.A2(n_803),
.B(n_737),
.C(n_782),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_775),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_756),
.A2(n_848),
.B(n_771),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_845),
.B(n_730),
.Y(n_971)
);

INVx3_ASAP7_75t_SL g972 ( 
.A(n_787),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_SL g973 ( 
.A1(n_735),
.A2(n_760),
.B(n_877),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_808),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_735),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_849),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_845),
.A2(n_730),
.B(n_733),
.Y(n_977)
);

INVx8_ASAP7_75t_L g978 ( 
.A(n_790),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_800),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_733),
.A2(n_811),
.B(n_864),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_764),
.A2(n_767),
.B(n_774),
.C(n_773),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_811),
.A2(n_772),
.B(n_750),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_R g983 ( 
.A(n_807),
.B(n_834),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_864),
.A2(n_790),
.B(n_802),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_749),
.B(n_790),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_812),
.A2(n_818),
.B(n_814),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_821),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_824),
.B(n_864),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_822),
.A2(n_829),
.B(n_831),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_852),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_726),
.B(n_786),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_724),
.B(n_596),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_761),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_726),
.A2(n_723),
.B1(n_810),
.B2(n_809),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_728),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_723),
.A2(n_748),
.B(n_604),
.C(n_726),
.Y(n_996)
);

CKINVDCx11_ASAP7_75t_R g997 ( 
.A(n_797),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_777),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_731),
.B(n_728),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_911),
.B(n_992),
.Y(n_1000)
);

NAND2x1_ASAP7_75t_L g1001 ( 
.A(n_916),
.B(n_957),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_987),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_SL g1003 ( 
.A1(n_880),
.A2(n_968),
.B(n_996),
.C(n_936),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_882),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_902),
.B(n_907),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_905),
.A2(n_878),
.B(n_902),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_977),
.A2(n_971),
.B(n_973),
.Y(n_1008)
);

NAND3x1_ASAP7_75t_L g1009 ( 
.A(n_921),
.B(n_887),
.C(n_912),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_908),
.B(n_991),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_939),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_991),
.B(n_909),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_994),
.A2(n_931),
.B1(n_951),
.B2(n_901),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_994),
.A2(n_885),
.B1(n_884),
.B2(n_944),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_906),
.B(n_983),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_952),
.A2(n_935),
.B(n_989),
.Y(n_1016)
);

AOI31xp67_ASAP7_75t_L g1017 ( 
.A1(n_879),
.A2(n_883),
.A3(n_904),
.B(n_946),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_953),
.B(n_960),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_930),
.A2(n_889),
.B(n_890),
.C(n_933),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_998),
.Y(n_1020)
);

AOI221xp5_ASAP7_75t_SL g1021 ( 
.A1(n_962),
.A2(n_924),
.B1(n_934),
.B2(n_966),
.C(n_883),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_958),
.A2(n_963),
.A3(n_886),
.B(n_897),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_943),
.B(n_978),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_970),
.A2(n_903),
.B(n_986),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_965),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_892),
.A2(n_894),
.B(n_966),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_918),
.B(n_881),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_SL g1028 ( 
.A(n_957),
.B(n_916),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_997),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_915),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_891),
.B(n_953),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_938),
.B(n_895),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_919),
.Y(n_1033)
);

AO21x1_ASAP7_75t_L g1034 ( 
.A1(n_924),
.A2(n_934),
.B(n_900),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_985),
.A2(n_922),
.B(n_927),
.Y(n_1035)
);

BUFx10_ASAP7_75t_L g1036 ( 
.A(n_956),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_920),
.B(n_893),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_923),
.Y(n_1038)
);

AOI211x1_ASAP7_75t_L g1039 ( 
.A1(n_964),
.A2(n_975),
.B(n_969),
.C(n_945),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_898),
.A2(n_981),
.A3(n_900),
.B(n_967),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_888),
.B(n_896),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_899),
.A2(n_999),
.B(n_950),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_882),
.A2(n_913),
.B(n_978),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_932),
.A2(n_979),
.B(n_974),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_913),
.A2(n_978),
.B(n_925),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_976),
.A2(n_993),
.B1(n_910),
.B2(n_940),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_995),
.A2(n_956),
.B(n_959),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_917),
.A2(n_910),
.B(n_940),
.C(n_941),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_SL g1049 ( 
.A1(n_988),
.A2(n_949),
.B(n_929),
.C(n_925),
.Y(n_1049)
);

AO21x1_ASAP7_75t_L g1050 ( 
.A1(n_925),
.A2(n_955),
.B(n_923),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_925),
.A2(n_923),
.B(n_926),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_948),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_926),
.A2(n_943),
.B(n_947),
.Y(n_1053)
);

AO31x2_ASAP7_75t_L g1054 ( 
.A1(n_926),
.A2(n_943),
.A3(n_961),
.B(n_942),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_990),
.A2(n_509),
.B1(n_510),
.B2(n_830),
.C(n_810),
.Y(n_1055)
);

AO32x2_ASAP7_75t_L g1056 ( 
.A1(n_972),
.A2(n_962),
.A3(n_994),
.B1(n_840),
.B2(n_861),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_937),
.B(n_902),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_SL g1058 ( 
.A1(n_902),
.A2(n_648),
.B(n_936),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_973),
.A2(n_980),
.B(n_723),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_910),
.B(n_940),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_971),
.A2(n_977),
.B(n_928),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_880),
.A2(n_968),
.B(n_996),
.C(n_936),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_902),
.Y(n_1063)
);

AOI211x1_ASAP7_75t_L g1064 ( 
.A1(n_991),
.A2(n_830),
.B(n_908),
.C(n_953),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_907),
.B(n_809),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_902),
.A2(n_723),
.B1(n_810),
.B2(n_809),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_921),
.A2(n_509),
.B1(n_510),
.B2(n_830),
.C(n_810),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_939),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_939),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_982),
.A2(n_971),
.A3(n_936),
.B(n_977),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_907),
.B(n_809),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_905),
.A2(n_878),
.B(n_902),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_906),
.A2(n_723),
.B(n_996),
.C(n_880),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_910),
.B(n_940),
.Y(n_1077)
);

NAND3x1_ASAP7_75t_L g1078 ( 
.A(n_921),
.B(n_705),
.C(n_509),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_902),
.B(n_907),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_994),
.B(n_596),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_973),
.A2(n_980),
.B(n_723),
.Y(n_1081)
);

AOI211x1_ASAP7_75t_L g1082 ( 
.A1(n_991),
.A2(n_830),
.B(n_908),
.C(n_953),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_905),
.A2(n_878),
.B(n_902),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_902),
.A2(n_648),
.B(n_936),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_939),
.Y(n_1085)
);

CKINVDCx11_ASAP7_75t_R g1086 ( 
.A(n_997),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_923),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_L g1088 ( 
.A(n_902),
.B(n_809),
.Y(n_1088)
);

INVx3_ASAP7_75t_SL g1089 ( 
.A(n_881),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_939),
.Y(n_1090)
);

AO32x2_ASAP7_75t_L g1091 ( 
.A1(n_962),
.A2(n_994),
.A3(n_840),
.B1(n_861),
.B2(n_954),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_902),
.B(n_907),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1093)
);

OA22x2_ASAP7_75t_L g1094 ( 
.A1(n_994),
.A2(n_407),
.B1(n_840),
.B2(n_861),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_902),
.B(n_907),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_984),
.A2(n_914),
.B(n_928),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_887),
.A2(n_809),
.B1(n_816),
.B2(n_810),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_939),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_994),
.B(n_596),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_907),
.B(n_809),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_982),
.A2(n_971),
.A3(n_936),
.B(n_977),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_SL g1102 ( 
.A1(n_902),
.A2(n_648),
.B(n_936),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_911),
.B(n_724),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_902),
.B(n_907),
.Y(n_1104)
);

INVx6_ASAP7_75t_L g1105 ( 
.A(n_948),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_996),
.A2(n_723),
.B(n_906),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_982),
.A2(n_971),
.A3(n_936),
.B(n_977),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_996),
.A2(n_723),
.B(n_906),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_882),
.B(n_723),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_939),
.Y(n_1110)
);

BUFx12f_ASAP7_75t_L g1111 ( 
.A(n_997),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_906),
.A2(n_723),
.B(n_596),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_905),
.A2(n_878),
.B(n_902),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_SL g1114 ( 
.A1(n_902),
.A2(n_648),
.B(n_936),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_902),
.A2(n_723),
.B1(n_810),
.B2(n_809),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1023),
.B(n_1060),
.Y(n_1116)
);

NOR2x1_ASAP7_75t_SL g1117 ( 
.A(n_1015),
.B(n_1023),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_1111),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1005),
.B(n_1079),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1006),
.Y(n_1120)
);

BUFx4f_ASAP7_75t_L g1121 ( 
.A(n_1089),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_1032),
.Y(n_1122)
);

INVx3_ASAP7_75t_SL g1123 ( 
.A(n_1105),
.Y(n_1123)
);

AOI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1097),
.A2(n_1106),
.B1(n_1108),
.B2(n_1063),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1065),
.A2(n_1072),
.B(n_1071),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_1008),
.A2(n_1059),
.B(n_1081),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1078),
.A2(n_1068),
.B1(n_1010),
.B2(n_1009),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1128)
);

OAI221xp5_ASAP7_75t_L g1129 ( 
.A1(n_1055),
.A2(n_1099),
.B1(n_1080),
.B2(n_1076),
.C(n_1112),
.Y(n_1129)
);

BUFx4_ASAP7_75t_R g1130 ( 
.A(n_1036),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1036),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1067),
.A2(n_1115),
.B1(n_1003),
.B2(n_1062),
.C(n_1031),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_1020),
.B(n_1057),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_1105),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1088),
.A2(n_1103),
.B1(n_1100),
.B2(n_1074),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1011),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1093),
.A2(n_1096),
.B(n_1026),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1069),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1034),
.A2(n_1083),
.A3(n_1075),
.B(n_1113),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1058),
.A2(n_1114),
.B(n_1084),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1070),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1023),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1102),
.A2(n_1014),
.B(n_1013),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1018),
.A2(n_1104),
.B(n_1013),
.C(n_1012),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1042),
.A2(n_1035),
.B(n_1061),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1041),
.B(n_1110),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1094),
.A2(n_1030),
.B1(n_1033),
.B2(n_1056),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_1021),
.A2(n_1044),
.B(n_1014),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1085),
.B(n_1098),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1066),
.A2(n_1017),
.B(n_1109),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_1027),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1025),
.A2(n_1037),
.B1(n_1048),
.B2(n_1090),
.Y(n_1152)
);

OR3x4_ASAP7_75t_SL g1153 ( 
.A(n_1056),
.B(n_1091),
.C(n_1049),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1054),
.Y(n_1154)
);

INVx3_ASAP7_75t_SL g1155 ( 
.A(n_1029),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1046),
.A2(n_1043),
.B(n_1047),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1039),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1051),
.A2(n_1045),
.B(n_1047),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1001),
.A2(n_1053),
.B(n_1050),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1028),
.A2(n_1004),
.B(n_1022),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_R g1161 ( 
.A(n_1086),
.B(n_1052),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1073),
.A2(n_1107),
.B(n_1101),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1056),
.B(n_1077),
.Y(n_1163)
);

AOI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_1028),
.A2(n_1053),
.B(n_1077),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1064),
.A2(n_1082),
.B1(n_1004),
.B2(n_1091),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1091),
.A2(n_1064),
.B1(n_1082),
.B2(n_1087),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1040),
.A2(n_1054),
.B(n_1038),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1087),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1005),
.B(n_1079),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1036),
.Y(n_1170)
);

AND2x2_ASAP7_75t_SL g1171 ( 
.A(n_1068),
.B(n_921),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1010),
.A2(n_902),
.B(n_991),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1019),
.A2(n_723),
.B(n_1076),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1068),
.A2(n_723),
.B(n_906),
.C(n_1076),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1068),
.A2(n_830),
.B1(n_921),
.B2(n_723),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1006),
.Y(n_1176)
);

CKINVDCx6p67_ASAP7_75t_R g1177 ( 
.A(n_1089),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1005),
.B(n_1079),
.Y(n_1178)
);

OAI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1068),
.A2(n_723),
.B1(n_1055),
.B2(n_816),
.C(n_810),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1006),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1006),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1078),
.A2(n_810),
.B1(n_816),
.B2(n_809),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1068),
.A2(n_830),
.B1(n_921),
.B2(n_723),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1105),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1002),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1005),
.B(n_907),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1105),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1005),
.B(n_907),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1068),
.A2(n_723),
.B(n_906),
.C(n_1076),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1068),
.A2(n_509),
.B1(n_1055),
.B2(n_809),
.C(n_816),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1008),
.A2(n_1034),
.A3(n_982),
.B(n_1007),
.Y(n_1191)
);

BUFx2_ASAP7_75t_R g1192 ( 
.A(n_1089),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1068),
.A2(n_810),
.B1(n_816),
.B2(n_809),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1078),
.A2(n_810),
.B1(n_816),
.B2(n_809),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1080),
.B(n_596),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1068),
.A2(n_1019),
.B(n_1015),
.C(n_723),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1000),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1002),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1020),
.B(n_881),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1019),
.A2(n_723),
.B(n_1076),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1024),
.A2(n_1016),
.B(n_1006),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1002),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1008),
.A2(n_1021),
.B(n_1007),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1002),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1002),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1119),
.B(n_1128),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_1135),
.B(n_1131),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1140),
.A2(n_1143),
.B(n_1144),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1169),
.B(n_1178),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1175),
.B(n_1183),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1193),
.A2(n_1190),
.B1(n_1183),
.B2(n_1175),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1168),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1144),
.A2(n_1200),
.B(n_1173),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1171),
.A2(n_1179),
.B1(n_1129),
.B2(n_1182),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1196),
.A2(n_1189),
.B(n_1174),
.C(n_1127),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1126),
.Y(n_1216)
);

AOI221x1_ASAP7_75t_SL g1217 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1133),
.B2(n_1152),
.C(n_1165),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1146),
.B(n_1163),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1171),
.B(n_1147),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1186),
.B(n_1188),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1126),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1149),
.B(n_1195),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1136),
.B(n_1138),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1151),
.A2(n_1174),
.B1(n_1189),
.B2(n_1132),
.Y(n_1224)
);

BUFx4_ASAP7_75t_R g1225 ( 
.A(n_1117),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1166),
.B(n_1157),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1172),
.B(n_1124),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1185),
.B(n_1205),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1130),
.Y(n_1229)
);

AOI211xp5_ASAP7_75t_L g1230 ( 
.A1(n_1150),
.A2(n_1199),
.B(n_1164),
.C(n_1123),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1204),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1168),
.Y(n_1232)
);

AOI31xp33_ASAP7_75t_L g1233 ( 
.A1(n_1161),
.A2(n_1166),
.A3(n_1184),
.B(n_1187),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1134),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1141),
.A2(n_1123),
.B(n_1202),
.C(n_1198),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1134),
.A2(n_1154),
.B1(n_1142),
.B2(n_1121),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1142),
.B(n_1158),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1170),
.B(n_1121),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1148),
.B(n_1162),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1177),
.B(n_1155),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1148),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1155),
.A2(n_1203),
.B(n_1153),
.C(n_1130),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1145),
.A2(n_1137),
.B(n_1125),
.Y(n_1245)
);

CKINVDCx6p67_ASAP7_75t_R g1246 ( 
.A(n_1118),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1192),
.B(n_1156),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1162),
.B(n_1191),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1191),
.B(n_1139),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_1201),
.B(n_1180),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1201),
.A2(n_1181),
.B(n_1176),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1193),
.A2(n_810),
.B1(n_816),
.B2(n_809),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1129),
.A2(n_1179),
.B(n_1196),
.C(n_1189),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1140),
.A2(n_1143),
.B(n_1144),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1129),
.A2(n_1179),
.B(n_1196),
.C(n_1189),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1142),
.B(n_1116),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1129),
.A2(n_1179),
.B(n_1196),
.C(n_1189),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1197),
.B(n_1122),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1177),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1129),
.A2(n_1179),
.B(n_1196),
.C(n_1189),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1129),
.A2(n_1179),
.B(n_1196),
.C(n_1189),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1248),
.B(n_1249),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1238),
.B(n_1242),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1227),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1216),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1242),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1216),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1225),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1240),
.B(n_1221),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1225),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1235),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1214),
.B(n_1253),
.Y(n_1272)
);

BUFx8_ASAP7_75t_L g1273 ( 
.A(n_1212),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1243),
.A2(n_1213),
.B(n_1254),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1223),
.Y(n_1275)
);

INVx5_ASAP7_75t_L g1276 ( 
.A(n_1238),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1208),
.B(n_1254),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1250),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1213),
.A2(n_1208),
.B(n_1244),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1215),
.A2(n_1211),
.B(n_1261),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1226),
.A2(n_1231),
.B(n_1228),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_1206),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1262),
.B(n_1218),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1262),
.B(n_1245),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1265),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1271),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1262),
.B(n_1245),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1269),
.B(n_1245),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1263),
.B(n_1251),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1277),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1265),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1276),
.B(n_1256),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1279),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1267),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1273),
.B(n_1259),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1267),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1282),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1276),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1263),
.B(n_1266),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1282),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1278),
.A2(n_1260),
.B(n_1219),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1266),
.B(n_1222),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1285),
.B(n_1282),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1286),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1286),
.Y(n_1306)
);

AOI222xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1298),
.A2(n_1224),
.B1(n_1252),
.B2(n_1264),
.C1(n_1278),
.C2(n_1283),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1292),
.Y(n_1308)
);

NOR2x1_ASAP7_75t_L g1309 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1302),
.A2(n_1277),
.B(n_1281),
.Y(n_1310)
);

NAND2xp33_ASAP7_75t_R g1311 ( 
.A(n_1296),
.B(n_1259),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1302),
.B(n_1272),
.C(n_1210),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1292),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1298),
.A2(n_1272),
.B1(n_1210),
.B2(n_1281),
.C(n_1217),
.Y(n_1314)
);

NOR4xp25_ASAP7_75t_L g1315 ( 
.A(n_1301),
.B(n_1236),
.C(n_1264),
.D(n_1233),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1295),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1294),
.Y(n_1317)
);

OAI211xp5_ASAP7_75t_L g1318 ( 
.A1(n_1301),
.A2(n_1230),
.B(n_1209),
.C(n_1281),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1284),
.A2(n_1277),
.B1(n_1229),
.B2(n_1283),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1284),
.A2(n_1277),
.B1(n_1229),
.B2(n_1268),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1291),
.A2(n_1277),
.B1(n_1281),
.B2(n_1280),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1291),
.A2(n_1277),
.B1(n_1281),
.B2(n_1280),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1300),
.B(n_1303),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1295),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1291),
.A2(n_1280),
.B1(n_1247),
.B2(n_1274),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1303),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1297),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1291),
.A2(n_1280),
.B1(n_1274),
.B2(n_1270),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1303),
.B(n_1285),
.Y(n_1329)
);

INVx5_ASAP7_75t_SL g1330 ( 
.A(n_1287),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_SL g1331 ( 
.A(n_1296),
.B(n_1212),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1297),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1291),
.B(n_1299),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1284),
.A2(n_1229),
.B1(n_1270),
.B2(n_1268),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1299),
.B(n_1293),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.B(n_1288),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1305),
.Y(n_1337)
);

AND4x1_ASAP7_75t_L g1338 ( 
.A(n_1315),
.B(n_1241),
.C(n_1239),
.D(n_1246),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_SL g1339 ( 
.A(n_1307),
.B(n_1220),
.C(n_1258),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1313),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1330),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1313),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1306),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1336),
.B(n_1290),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1316),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1308),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1330),
.Y(n_1347)
);

AND2x6_ASAP7_75t_SL g1348 ( 
.A(n_1333),
.B(n_1246),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1327),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1304),
.B(n_1289),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1332),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1332),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1336),
.B(n_1290),
.Y(n_1353)
);

NOR2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1312),
.B(n_1232),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1324),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1317),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1309),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1330),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1340),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1355),
.B(n_1314),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1341),
.B(n_1299),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1355),
.B(n_1326),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1340),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1337),
.B(n_1343),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1339),
.B(n_1314),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1340),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1337),
.B(n_1275),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1344),
.B(n_1335),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1343),
.B(n_1275),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1356),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1344),
.B(n_1323),
.Y(n_1371)
);

NAND4xp25_ASAP7_75t_L g1372 ( 
.A(n_1339),
.B(n_1312),
.C(n_1310),
.D(n_1318),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1341),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1338),
.B(n_1318),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1346),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1344),
.B(n_1335),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_SL g1377 ( 
.A(n_1338),
.B(n_1311),
.C(n_1331),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1342),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1345),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1346),
.B(n_1315),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1345),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1350),
.B(n_1319),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1350),
.B(n_1319),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1345),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1349),
.B(n_1329),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1354),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1350),
.B(n_1329),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1307),
.C(n_1207),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1341),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1357),
.A2(n_1310),
.B(n_1280),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1353),
.B(n_1330),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1356),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1348),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1351),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1370),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1384),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1364),
.B(n_1360),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1393),
.B(n_1357),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1384),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1370),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1375),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1375),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1361),
.B(n_1341),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1341),
.Y(n_1404)
);

AOI32xp33_ASAP7_75t_L g1405 ( 
.A1(n_1365),
.A2(n_1325),
.A3(n_1322),
.B1(n_1321),
.B2(n_1328),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1392),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1388),
.B(n_1354),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1388),
.B(n_1349),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1374),
.B(n_1347),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1373),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1359),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1367),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1368),
.B(n_1347),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1373),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1380),
.B(n_1351),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1391),
.B(n_1347),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1374),
.A2(n_1274),
.B1(n_1320),
.B2(n_1334),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_L g1418 ( 
.A(n_1372),
.B(n_1347),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1362),
.B(n_1351),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1391),
.B(n_1347),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1369),
.B(n_1352),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1392),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1363),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1386),
.B(n_1232),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1389),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1385),
.B(n_1352),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1382),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1418),
.B(n_1268),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1402),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1425),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1398),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1398),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1399),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1416),
.B(n_1376),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1429),
.B(n_1371),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1412),
.B(n_1389),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1399),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1399),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_1397),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1409),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1409),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1397),
.B(n_1387),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1401),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1418),
.A2(n_1291),
.B1(n_1390),
.B2(n_1274),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1401),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1396),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1410),
.Y(n_1449)
);

INVx3_ASAP7_75t_SL g1450 ( 
.A(n_1410),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1414),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1409),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1403),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1433),
.B(n_1212),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1449),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1415),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1435),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1433),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1435),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1454),
.A2(n_1377),
.B1(n_1417),
.B2(n_1405),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1441),
.A2(n_1377),
.B1(n_1417),
.B2(n_1405),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1449),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1449),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1444),
.B(n_1421),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1443),
.B(n_1212),
.Y(n_1466)
);

AOI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1430),
.A2(n_1427),
.B(n_1414),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1446),
.A2(n_1413),
.B1(n_1383),
.B2(n_1416),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1450),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1442),
.A2(n_1404),
.B(n_1403),
.C(n_1396),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1439),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1431),
.B(n_1420),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1436),
.B(n_1420),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1469),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1469),
.B(n_1453),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1459),
.B(n_1450),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1456),
.B(n_1451),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1473),
.B(n_1472),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1455),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1465),
.B(n_1437),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1436),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1470),
.B(n_1451),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1461),
.A2(n_1452),
.B(n_1432),
.Y(n_1484)
);

NAND4xp25_ASAP7_75t_L g1485 ( 
.A(n_1484),
.B(n_1462),
.C(n_1457),
.D(n_1467),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1474),
.A2(n_1432),
.B1(n_1468),
.B2(n_1455),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1474),
.B(n_1438),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1483),
.A2(n_1466),
.B(n_1443),
.Y(n_1488)
);

AND3x1_ASAP7_75t_L g1489 ( 
.A(n_1476),
.B(n_1445),
.C(n_1471),
.Y(n_1489)
);

NOR3xp33_ASAP7_75t_L g1490 ( 
.A(n_1475),
.B(n_1447),
.C(n_1448),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1482),
.A2(n_1466),
.B1(n_1404),
.B2(n_1413),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1478),
.A2(n_1447),
.B(n_1460),
.C(n_1458),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_SL g1493 ( 
.A(n_1481),
.B(n_1444),
.C(n_1440),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1477),
.B(n_1449),
.C(n_1466),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1479),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1487),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1486),
.A2(n_1480),
.B(n_1449),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1493),
.A2(n_1411),
.B(n_1424),
.C(n_1419),
.Y(n_1498)
);

OAI22x1_ASAP7_75t_L g1499 ( 
.A1(n_1491),
.A2(n_1413),
.B1(n_1411),
.B2(n_1424),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1494),
.Y(n_1500)
);

OAI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1497),
.A2(n_1485),
.B1(n_1489),
.B2(n_1490),
.C(n_1488),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1500),
.B(n_1495),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1496),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1498),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1499),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1499),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1501),
.A2(n_1413),
.B1(n_1419),
.B2(n_1492),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1506),
.B(n_1423),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1505),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1502),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1503),
.B(n_1423),
.Y(n_1511)
);

AND3x4_ASAP7_75t_L g1512 ( 
.A(n_1508),
.B(n_1234),
.C(n_1504),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1509),
.A2(n_1395),
.B1(n_1422),
.B2(n_1406),
.C(n_1400),
.Y(n_1513)
);

AND3x4_ASAP7_75t_L g1514 ( 
.A(n_1508),
.B(n_1234),
.C(n_1395),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1514),
.B(n_1511),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1515),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1516),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1517),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1518),
.B(n_1510),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1519),
.A2(n_1507),
.B(n_1513),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1519),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1521),
.A2(n_1512),
.B1(n_1400),
.B2(n_1406),
.Y(n_1522)
);

XNOR2xp5_ASAP7_75t_L g1523 ( 
.A(n_1520),
.B(n_1426),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1523),
.A2(n_1522),
.B(n_1426),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1523),
.A2(n_1406),
.B(n_1400),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1524),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1525),
.A2(n_1422),
.B1(n_1379),
.B2(n_1378),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1526),
.A2(n_1422),
.B1(n_1394),
.B2(n_1366),
.C(n_1381),
.Y(n_1528)
);

AOI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1528),
.A2(n_1527),
.B(n_1428),
.C(n_1237),
.Y(n_1529)
);


endmodule