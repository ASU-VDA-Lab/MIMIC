module fake_jpeg_24663_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_47),
.Y(n_78)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_28),
.B1(n_49),
.B2(n_44),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_23),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_54),
.B(n_62),
.Y(n_108)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_21),
.B1(n_34),
.B2(n_36),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_21),
.B1(n_34),
.B2(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_73),
.B1(n_25),
.B2(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_26),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_36),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_101),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_96),
.B1(n_19),
.B2(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_110),
.Y(n_137)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_38),
.C(n_37),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_19),
.C(n_37),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_0),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_20),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_113),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_23),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_17),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_17),
.B1(n_27),
.B2(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_19),
.B1(n_18),
.B2(n_29),
.Y(n_138)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_20),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_124),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_80),
.B1(n_79),
.B2(n_77),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_138),
.B1(n_154),
.B2(n_29),
.Y(n_164)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_128),
.Y(n_174)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_132),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_17),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_20),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_149),
.C(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_68),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_157),
.Y(n_187)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_20),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_52),
.B1(n_56),
.B2(n_30),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_52),
.B1(n_71),
.B2(n_35),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_121),
.B1(n_92),
.B2(n_93),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_20),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_104),
.B(n_119),
.C(n_23),
.D(n_98),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_189),
.B(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_172),
.B1(n_181),
.B2(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_168),
.B(n_171),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_107),
.C(n_93),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_177),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_179),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_107),
.C(n_98),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_129),
.B(n_23),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_120),
.C(n_114),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_23),
.B1(n_31),
.B2(n_2),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_123),
.B1(n_116),
.B2(n_24),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_97),
.B1(n_122),
.B2(n_31),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_193),
.B1(n_164),
.B2(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_136),
.A2(n_97),
.B1(n_101),
.B2(n_87),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_186),
.B1(n_161),
.B2(n_192),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_136),
.B(n_148),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_218),
.B(n_177),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_213),
.B1(n_190),
.B2(n_162),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_149),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_210),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_140),
.A3(n_157),
.B1(n_131),
.B2(n_132),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_131),
.B1(n_150),
.B2(n_143),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_153),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_139),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_201),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_190),
.B1(n_178),
.B2(n_168),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_243),
.B1(n_0),
.B2(n_1),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_248),
.B1(n_205),
.B2(n_239),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_176),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_230),
.B(n_234),
.Y(n_253)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_241),
.B(n_224),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_170),
.B1(n_166),
.B2(n_194),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_245),
.B1(n_203),
.B2(n_211),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_170),
.B1(n_159),
.B2(n_126),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_194),
.B1(n_27),
.B2(n_26),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_124),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_199),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_236),
.C(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_264),
.C(n_267),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_258),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_254),
.B(n_263),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_206),
.B(n_220),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_246),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_204),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_200),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_261),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_227),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_210),
.C(n_200),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_202),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_16),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_16),
.C(n_1),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_248),
.B1(n_232),
.B2(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_231),
.B(n_3),
.Y(n_300)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_284),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_228),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_229),
.C(n_230),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_286),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_231),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_241),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_259),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_250),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_291),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_300),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_268),
.B(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_275),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_228),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_298),
.C(n_300),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_235),
.B(n_233),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_278),
.C(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_0),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_310),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_278),
.C(n_277),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_290),
.B1(n_287),
.B2(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_301),
.B(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_315),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_289),
.B(n_3),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_318),
.B1(n_308),
.B2(n_5),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_310),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_317),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_313),
.B(n_309),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_326),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_319),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_322),
.C(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_328),
.C(n_5),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_4),
.C(n_7),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_7),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule