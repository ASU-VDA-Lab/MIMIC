module fake_netlist_5_2221_n_1082 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_267, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1082);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1082;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_523;
wire n_315;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_643;
wire n_367;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_443;
wire n_677;
wire n_372;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_516;
wire n_498;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_556;
wire n_1063;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_341;
wire n_394;
wire n_992;
wire n_1049;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_519;
wire n_406;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_962;
wire n_400;
wire n_930;
wire n_436;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_866;
wire n_796;
wire n_573;
wire n_969;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_571;
wire n_338;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_630;
wire n_420;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_513;
wire n_425;
wire n_647;
wire n_527;
wire n_407;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_754;
wire n_712;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_639;
wire n_914;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_985;
wire n_904;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_9),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_241),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_85),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_134),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_65),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_102),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_8),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_174),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_137),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_124),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_167),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_116),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_138),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_77),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_57),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_155),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_51),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_75),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_74),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_122),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_98),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_207),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_33),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_5),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_199),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_48),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_158),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_61),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_147),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_243),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_113),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_108),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_179),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_15),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_17),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_231),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_259),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_42),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_27),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_112),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_183),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_72),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_56),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_110),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_44),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_162),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_126),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_32),
.B(n_220),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_213),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_120),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_168),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_232),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_188),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_2),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_187),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_0),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_269),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_18),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_210),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_36),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_256),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_152),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_240),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_88),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_52),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_215),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_139),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_200),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_236),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_257),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_90),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_251),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_193),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_148),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_169),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_93),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_212),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_222),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_192),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_87),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_185),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_58),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_265),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_62),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_23),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_181),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_141),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_83),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_247),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_35),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_173),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_25),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_234),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_67),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_94),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_178),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_190),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_219),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_160),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_76),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_23),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_157),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_14),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_2),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_238),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_130),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_154),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_252),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_196),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_239),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_28),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_45),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_235),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_60),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_159),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_145),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_225),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_264),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_202),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_31),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_184),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_171),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_151),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_254),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_86),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_99),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_204),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_14),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_244),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_89),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_47),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_253),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_136),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_55),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_248),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_258),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_164),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_211),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_263),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_29),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_5),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_209),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_4),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_223),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_337),
.B(n_0),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_270),
.B(n_287),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_337),
.B(n_1),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_332),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_285),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_339),
.B(n_1),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_332),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_343),
.B(n_3),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_3),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_318),
.B(n_4),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_321),
.B(n_6),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_354),
.B(n_6),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_332),
.B(n_37),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_332),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_325),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_366),
.A2(n_402),
.B1(n_350),
.B2(n_331),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_431),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_281),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_329),
.Y(n_464)
);

BUFx12f_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_288),
.B(n_7),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_397),
.B(n_7),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_324),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_9),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_351),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_278),
.B(n_10),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_10),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_388),
.B(n_424),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_359),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_272),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_359),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_433),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_298),
.B(n_11),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_433),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_433),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_303),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_273),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_319),
.B(n_11),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_397),
.B(n_282),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_271),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_276),
.A2(n_12),
.B(n_13),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_277),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_280),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_291),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_348),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_284),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_275),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_289),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_374),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_292),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_295),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_299),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_347),
.A2(n_400),
.B1(n_294),
.B2(n_320),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_282),
.A2(n_296),
.B1(n_387),
.B2(n_357),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_279),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_296),
.B(n_12),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_300),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_302),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_304),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_307),
.Y(n_514)
);

CKINVDCx6p67_ASAP7_75t_R g515 ( 
.A(n_301),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_283),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_308),
.A2(n_13),
.B(n_16),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_309),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_310),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_316),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_322),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_286),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_323),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_290),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_357),
.B(n_16),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_333),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_387),
.B(n_17),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_334),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_410),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_335),
.B(n_38),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_336),
.B(n_19),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_297),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_305),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_516),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_449),
.B(n_362),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g537 ( 
.A1(n_530),
.A2(n_274),
.B1(n_384),
.B2(n_428),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_444),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_342),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_461),
.B(n_391),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_345),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_492),
.A2(n_274),
.B1(n_384),
.B2(n_428),
.Y(n_547)
);

AO21x2_ASAP7_75t_L g548 ( 
.A1(n_476),
.A2(n_340),
.B(n_346),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_441),
.B(n_412),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_450),
.B(n_416),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_353),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_497),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_446),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_448),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_457),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_484),
.B(n_419),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_457),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_459),
.B(n_306),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_490),
.B(n_364),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_490),
.B(n_365),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_507),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_484),
.B(n_432),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_464),
.B(n_20),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_518),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

BUFx8_ASAP7_75t_SL g574 ( 
.A(n_480),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_462),
.B(n_312),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_443),
.B(n_313),
.Y(n_578)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_508),
.B(n_526),
.C(n_471),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_442),
.A2(n_440),
.B1(n_438),
.B2(n_314),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_456),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_523),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_456),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_479),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_315),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_369),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_456),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_479),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_493),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_481),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_481),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_525),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_466),
.B(n_317),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_522),
.B(n_370),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_511),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_482),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_519),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_460),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_482),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_498),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_532),
.B(n_326),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_477),
.B(n_371),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_610),
.B(n_445),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_549),
.B(n_489),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_L g615 ( 
.A1(n_547),
.A2(n_453),
.B(n_454),
.C(n_451),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_592),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_556),
.B(n_548),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_549),
.B(n_465),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_539),
.B(n_510),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_551),
.B(n_489),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_578),
.B(n_528),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_578),
.B(n_515),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_547),
.B(n_532),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_536),
.B(n_489),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_564),
.B(n_327),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_536),
.B(n_445),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_543),
.B(n_445),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_608),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_548),
.B(n_473),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_605),
.B(n_328),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_610),
.B(n_527),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_586),
.B(n_546),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_559),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g635 ( 
.A(n_580),
.B(n_473),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_478),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_575),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_531),
.B(n_491),
.Y(n_638)
);

BUFx8_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_553),
.B(n_473),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_585),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_595),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_558),
.B(n_495),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_560),
.B(n_483),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_561),
.B(n_483),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_585),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_612),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_600),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_579),
.A2(n_611),
.B(n_612),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_556),
.B(n_502),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_502),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_562),
.B(n_568),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_535),
.B(n_330),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_483),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_554),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_590),
.B(n_494),
.Y(n_656)
);

OAI221xp5_ASAP7_75t_L g657 ( 
.A1(n_598),
.A2(n_503),
.B1(n_495),
.B2(n_496),
.C(n_501),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_555),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_535),
.B(n_338),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_550),
.A2(n_467),
.B1(n_531),
.B2(n_411),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_604),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_488),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_488),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_593),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_583),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_542),
.B(n_496),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_544),
.B(n_341),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_611),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_537),
.B(n_467),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_598),
.A2(n_503),
.B(n_501),
.C(n_463),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_565),
.B(n_513),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_566),
.B(n_513),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_583),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_544),
.B(n_352),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_606),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_554),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_612),
.A2(n_531),
.B1(n_494),
.B2(n_517),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_588),
.B(n_488),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_537),
.B(n_355),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_L g683 ( 
.A(n_550),
.B(n_378),
.C(n_377),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_606),
.Y(n_684)
);

NOR2x1p5_ASAP7_75t_L g685 ( 
.A(n_589),
.B(n_485),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_612),
.A2(n_531),
.B1(n_517),
.B2(n_520),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_599),
.B(n_513),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_597),
.B(n_504),
.Y(n_688)
);

O2A1O1Ixp5_ASAP7_75t_L g689 ( 
.A1(n_576),
.A2(n_520),
.B(n_468),
.C(n_474),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_609),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_602),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_612),
.B(n_504),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_562),
.A2(n_529),
.B1(n_504),
.B2(n_475),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_619),
.B(n_568),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_621),
.B(n_557),
.C(n_552),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_633),
.A2(n_590),
.B(n_581),
.Y(n_696)
);

OA22x2_ASAP7_75t_L g697 ( 
.A1(n_623),
.A2(n_485),
.B1(n_486),
.B2(n_470),
.Y(n_697)
);

CKINVDCx14_ASAP7_75t_R g698 ( 
.A(n_630),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_643),
.B(n_596),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_617),
.A2(n_590),
.B(n_581),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_636),
.B(n_569),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_632),
.B(n_572),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_671),
.B(n_574),
.Y(n_703)
);

BUFx4f_ASAP7_75t_L g704 ( 
.A(n_652),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_674),
.B(n_576),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_649),
.A2(n_584),
.B1(n_379),
.B2(n_381),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_658),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_617),
.A2(n_590),
.B(n_584),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_414),
.B1(n_382),
.B2(n_383),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_618),
.B(n_573),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_634),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_555),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_638),
.A2(n_392),
.B(n_385),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_587),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_638),
.A2(n_417),
.B1(n_415),
.B2(n_394),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

O2A1O1Ixp5_ASAP7_75t_L g717 ( 
.A1(n_689),
.A2(n_418),
.B(n_395),
.C(n_396),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_655),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_686),
.A2(n_421),
.B1(n_406),
.B2(n_408),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_661),
.B(n_587),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_639),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_615),
.A2(n_423),
.B(n_436),
.C(n_413),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_628),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_685),
.B(n_582),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_642),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_639),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_692),
.A2(n_607),
.B(n_603),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_680),
.A2(n_425),
.B(n_420),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_669),
.A2(n_426),
.B1(n_427),
.B2(n_429),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_692),
.A2(n_603),
.B(n_545),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_687),
.B(n_434),
.Y(n_731)
);

BUFx2_ASAP7_75t_R g732 ( 
.A(n_682),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_670),
.B(n_356),
.Y(n_733)
);

OR2x6_ASAP7_75t_SL g734 ( 
.A(n_672),
.B(n_358),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_683),
.A2(n_398),
.B1(n_361),
.B2(n_363),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_629),
.A2(n_591),
.B(n_585),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_622),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_656),
.A2(n_541),
.B(n_540),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_679),
.B(n_486),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_691),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_647),
.A2(n_591),
.B(n_585),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_614),
.B(n_470),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_656),
.A2(n_390),
.B(n_367),
.Y(n_744)
);

OAI321xp33_ASAP7_75t_L g745 ( 
.A1(n_657),
.A2(n_529),
.A3(n_594),
.B1(n_591),
.B2(n_25),
.C(n_26),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_648),
.Y(n_746)
);

INVx6_ASAP7_75t_L g747 ( 
.A(n_641),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_647),
.A2(n_594),
.B(n_591),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_659),
.B(n_662),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_677),
.B(n_360),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_625),
.A2(n_393),
.B1(n_372),
.B2(n_373),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_673),
.A2(n_407),
.B(n_375),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_647),
.A2(n_594),
.B(n_401),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_672),
.A2(n_409),
.B1(n_376),
.B2(n_386),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_626),
.A2(n_594),
.B(n_435),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_664),
.B(n_529),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_651),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_693),
.B(n_567),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_650),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_624),
.A2(n_430),
.B1(n_389),
.B2(n_368),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_641),
.Y(n_762)
);

OAI22x1_ASAP7_75t_L g763 ( 
.A1(n_653),
.A2(n_567),
.B1(n_660),
.B2(n_631),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_650),
.A2(n_132),
.B(n_266),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_690),
.B(n_39),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_688),
.A2(n_133),
.B(n_262),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_635),
.A2(n_131),
.B1(n_255),
.B2(n_250),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_627),
.A2(n_128),
.B(n_249),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_716),
.B(n_676),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_707),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_762),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_762),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_713),
.A2(n_667),
.B(n_620),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_725),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_694),
.A2(n_715),
.B1(n_709),
.B2(n_719),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_739),
.A2(n_654),
.B(n_681),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_746),
.B(n_668),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_699),
.B(n_678),
.Y(n_778)
);

AOI21x1_ASAP7_75t_L g779 ( 
.A1(n_700),
.A2(n_645),
.B(n_666),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_708),
.A2(n_684),
.B(n_665),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_752),
.B(n_613),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_722),
.A2(n_644),
.B(n_640),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_738),
.A2(n_704),
.B1(n_744),
.B2(n_728),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_759),
.A2(n_641),
.B1(n_646),
.B2(n_24),
.C(n_26),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_701),
.B(n_646),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_711),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_717),
.A2(n_646),
.B(n_129),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_742),
.A2(n_267),
.B(n_127),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_706),
.A2(n_125),
.B(n_245),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_765),
.B(n_40),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_726),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_729),
.A2(n_21),
.A3(n_22),
.B(n_24),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_704),
.B(n_22),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_760),
.A2(n_705),
.B1(n_755),
.B2(n_758),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_698),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_710),
.B(n_41),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_696),
.A2(n_714),
.B(n_749),
.Y(n_797)
);

BUFx12f_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

OAI21x1_ASAP7_75t_SL g799 ( 
.A1(n_768),
.A2(n_142),
.B(n_43),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_737),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_740),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_736),
.A2(n_143),
.B(n_46),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_703),
.B(n_27),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_740),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_49),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_697),
.Y(n_806)
);

AND2x4_ASAP7_75t_SL g807 ( 
.A(n_724),
.B(n_50),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_748),
.A2(n_246),
.B(n_54),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_727),
.A2(n_242),
.B(n_59),
.Y(n_809)
);

AOI221x1_ASAP7_75t_L g810 ( 
.A1(n_763),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_743),
.B(n_68),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_730),
.A2(n_69),
.B(n_70),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_754),
.A2(n_741),
.B(n_723),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_731),
.B(n_71),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_723),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_741),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_762),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_774),
.Y(n_818)
);

AO21x2_ASAP7_75t_L g819 ( 
.A1(n_787),
.A2(n_789),
.B(n_782),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_778),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_806),
.B(n_734),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_780),
.A2(n_764),
.B(n_766),
.Y(n_822)
);

NOR2x1_ASAP7_75t_SL g823 ( 
.A(n_817),
.B(n_720),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_791),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_779),
.A2(n_756),
.B(n_757),
.Y(n_825)
);

INVx6_ASAP7_75t_L g826 ( 
.A(n_817),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_785),
.B(n_733),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_776),
.A2(n_695),
.B(n_765),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_812),
.A2(n_753),
.B(n_767),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_804),
.Y(n_830)
);

AOI22x1_ASAP7_75t_L g831 ( 
.A1(n_797),
.A2(n_718),
.B1(n_745),
.B2(n_750),
.Y(n_831)
);

OAI21x1_ASAP7_75t_L g832 ( 
.A1(n_809),
.A2(n_761),
.B(n_751),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_786),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_788),
.A2(n_735),
.B(n_747),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_800),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_808),
.A2(n_747),
.B(n_712),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_783),
.A2(n_732),
.A3(n_78),
.B(n_79),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_815),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_770),
.Y(n_839)
);

AOI21x1_ASAP7_75t_L g840 ( 
.A1(n_794),
.A2(n_73),
.B(n_80),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_777),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_813),
.A2(n_81),
.B(n_82),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_801),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_795),
.Y(n_844)
);

AO21x2_ASAP7_75t_L g845 ( 
.A1(n_787),
.A2(n_84),
.B(n_92),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_798),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_775),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_782),
.A2(n_100),
.B(n_101),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_814),
.A2(n_103),
.B(n_105),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_816),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_825),
.A2(n_842),
.B(n_836),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_818),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_818),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_838),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_838),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_833),
.Y(n_856)
);

AO21x2_ASAP7_75t_L g857 ( 
.A1(n_819),
.A2(n_773),
.B(n_775),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_820),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_826),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_850),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_850),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_821),
.B(n_790),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_835),
.Y(n_863)
);

BUFx6f_ASAP7_75t_SL g864 ( 
.A(n_841),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_830),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_843),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_848),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_848),
.Y(n_868)
);

AO21x2_ASAP7_75t_L g869 ( 
.A1(n_819),
.A2(n_773),
.B(n_805),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_828),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_823),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_842),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_827),
.B(n_801),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_821),
.B(n_793),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_834),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_847),
.B(n_817),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_847),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_839),
.B(n_781),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_SL g879 ( 
.A1(n_829),
.A2(n_784),
.B(n_811),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_852),
.B(n_837),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_866),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_863),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_852),
.B(n_837),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_859),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_859),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_873),
.B(n_803),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_863),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_874),
.B(n_837),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_853),
.B(n_837),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_878),
.A2(n_831),
.B1(n_807),
.B2(n_844),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_853),
.B(n_792),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_865),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_865),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_854),
.B(n_792),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_858),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_878),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_877),
.A2(n_819),
.B1(n_845),
.B2(n_796),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_871),
.B(n_771),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_854),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_862),
.B(n_777),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_856),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_860),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_855),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_859),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_862),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_855),
.B(n_861),
.Y(n_906)
);

AND2x2_ASAP7_75t_SL g907 ( 
.A(n_877),
.B(n_802),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_861),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_860),
.B(n_792),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_857),
.B(n_876),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_857),
.B(n_845),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_870),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_876),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_912),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_912),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_910),
.B(n_909),
.Y(n_916)
);

AND2x4_ASAP7_75t_SL g917 ( 
.A(n_913),
.B(n_876),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_910),
.B(n_857),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_899),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_909),
.B(n_869),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_891),
.B(n_869),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_899),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_886),
.B(n_810),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_896),
.B(n_870),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_881),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_895),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_891),
.B(n_869),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_884),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_901),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_903),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_888),
.B(n_867),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_906),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_905),
.B(n_824),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_902),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_911),
.B(n_867),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_913),
.B(n_867),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_913),
.B(n_876),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_913),
.B(n_875),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_882),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_906),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_903),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_884),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_894),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_908),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_908),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_887),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_894),
.B(n_880),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_900),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_880),
.B(n_868),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_892),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_946),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_916),
.B(n_911),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_916),
.B(n_883),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_918),
.B(n_883),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_934),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_926),
.B(n_893),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_948),
.B(n_889),
.Y(n_957)
);

AND3x2_ASAP7_75t_L g958 ( 
.A(n_950),
.B(n_889),
.C(n_898),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_946),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_914),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_939),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_924),
.B(n_890),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_917),
.B(n_937),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_947),
.B(n_898),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_943),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_943),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_940),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_914),
.Y(n_969)
);

NAND2x1_ASAP7_75t_L g970 ( 
.A(n_937),
.B(n_885),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_938),
.B(n_937),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_915),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_935),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_925),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_925),
.B(n_907),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_947),
.B(n_868),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_918),
.B(n_898),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_915),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_931),
.B(n_868),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_919),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_974),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_955),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_SL g983 ( 
.A(n_958),
.B(n_917),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_963),
.A2(n_933),
.B1(n_923),
.B2(n_845),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_960),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_974),
.Y(n_986)
);

AND2x4_ASAP7_75t_SL g987 ( 
.A(n_965),
.B(n_942),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_951),
.Y(n_988)
);

NOR2x1p5_ASAP7_75t_SL g989 ( 
.A(n_979),
.B(n_840),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_956),
.B(n_932),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_957),
.B(n_920),
.Y(n_991)
);

NAND3x2_ASAP7_75t_L g992 ( 
.A(n_976),
.B(n_846),
.C(n_931),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_977),
.B(n_949),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_962),
.Y(n_994)
);

NOR4xp25_ASAP7_75t_L g995 ( 
.A(n_975),
.B(n_879),
.C(n_897),
.D(n_944),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_952),
.B(n_935),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_953),
.B(n_949),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_951),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_968),
.B(n_920),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_959),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_970),
.B(n_936),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_983),
.A2(n_966),
.B1(n_967),
.B2(n_942),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_995),
.A2(n_954),
.B(n_973),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_990),
.B(n_973),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_982),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_959),
.Y(n_1006)
);

OAI32xp33_ASAP7_75t_L g1007 ( 
.A1(n_981),
.A2(n_954),
.A3(n_980),
.B1(n_928),
.B2(n_936),
.Y(n_1007)
);

AOI211x1_ASAP7_75t_L g1008 ( 
.A1(n_999),
.A2(n_927),
.B(n_921),
.C(n_849),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_991),
.B(n_971),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_992),
.A2(n_995),
.B(n_984),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_983),
.A2(n_984),
.B1(n_1001),
.B2(n_996),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_985),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_1001),
.A2(n_964),
.B1(n_971),
.B2(n_864),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_1001),
.B(n_958),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_997),
.B(n_971),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1000),
.B(n_921),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_994),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_993),
.B(n_964),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_986),
.B(n_927),
.Y(n_1019)
);

AOI222xp33_ASAP7_75t_L g1020 ( 
.A1(n_989),
.A2(n_864),
.B1(n_897),
.B2(n_769),
.C1(n_907),
.C2(n_945),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_1005),
.B(n_988),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_1010),
.A2(n_928),
.B(n_987),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1012),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1013),
.A2(n_938),
.B1(n_942),
.B2(n_969),
.Y(n_1024)
);

AOI222xp33_ASAP7_75t_L g1025 ( 
.A1(n_1003),
.A2(n_1011),
.B1(n_1014),
.B2(n_1004),
.C1(n_1002),
.C2(n_1007),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_1014),
.B(n_942),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_1019),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_1020),
.A2(n_978),
.B(n_972),
.Y(n_1028)
);

AOI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1017),
.A2(n_942),
.B(n_972),
.C(n_969),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1009),
.A2(n_938),
.B(n_885),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1015),
.A2(n_978),
.B1(n_961),
.B2(n_944),
.Y(n_1031)
);

AOI211xp5_ASAP7_75t_L g1032 ( 
.A1(n_1006),
.A2(n_961),
.B(n_884),
.C(n_904),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1016),
.B(n_919),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1008),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1010),
.A2(n_832),
.B(n_930),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_1010),
.A2(n_799),
.B(n_941),
.Y(n_1036)
);

OAI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_1014),
.A2(n_941),
.B1(n_930),
.B2(n_922),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_1004),
.B(n_922),
.Y(n_1038)
);

AOI211xp5_ASAP7_75t_L g1039 ( 
.A1(n_1035),
.A2(n_1022),
.B(n_1034),
.C(n_1026),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1027),
.B(n_824),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1025),
.A2(n_844),
.B(n_832),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1030),
.A2(n_829),
.B(n_836),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_1038),
.B(n_864),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_L g1044 ( 
.A(n_1036),
.B(n_904),
.C(n_884),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1023),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1024),
.A2(n_904),
.B1(n_872),
.B2(n_802),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1021),
.B(n_1033),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1032),
.B(n_872),
.C(n_904),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_1028),
.A2(n_822),
.B(n_834),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1037),
.A2(n_822),
.B(n_825),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1031),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_1029),
.A2(n_769),
.B1(n_875),
.B2(n_771),
.C(n_772),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1034),
.A2(n_875),
.B1(n_826),
.B2(n_851),
.Y(n_1053)
);

AOI31xp33_ASAP7_75t_L g1054 ( 
.A1(n_1025),
.A2(n_106),
.A3(n_107),
.B(n_109),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_1034),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.C(n_117),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1025),
.A2(n_851),
.B(n_119),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_1054),
.B(n_118),
.Y(n_1057)
);

NAND4xp25_ASAP7_75t_L g1058 ( 
.A(n_1041),
.B(n_121),
.C(n_135),
.D(n_140),
.Y(n_1058)
);

NAND5xp2_ASAP7_75t_L g1059 ( 
.A(n_1039),
.B(n_1052),
.C(n_1055),
.D(n_1051),
.E(n_1040),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1056),
.B(n_144),
.C(n_146),
.Y(n_1060)
);

AND3x2_ASAP7_75t_L g1061 ( 
.A(n_1043),
.B(n_149),
.C(n_150),
.Y(n_1061)
);

AND5x1_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_1049),
.C(n_1046),
.D(n_1044),
.E(n_1048),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_L g1063 ( 
.A(n_1058),
.B(n_1057),
.C(n_1060),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1061),
.B(n_1047),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_L g1065 ( 
.A(n_1059),
.B(n_1053),
.C(n_1045),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_L g1066 ( 
.A(n_1059),
.B(n_1042),
.C(n_1050),
.Y(n_1066)
);

NAND4xp75_ASAP7_75t_L g1067 ( 
.A(n_1064),
.B(n_1047),
.C(n_156),
.D(n_163),
.Y(n_1067)
);

NOR2x1p5_ASAP7_75t_L g1068 ( 
.A(n_1062),
.B(n_153),
.Y(n_1068)
);

NAND4xp75_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_1065),
.C(n_1063),
.D(n_170),
.Y(n_1069)
);

OAI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1066),
.A2(n_165),
.B(n_166),
.C(n_176),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_1067),
.Y(n_1071)
);

AND3x4_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_826),
.C(n_180),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1068),
.Y(n_1073)
);

OAI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_177),
.B(n_182),
.C(n_186),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_191),
.B1(n_195),
.B2(n_197),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1071),
.Y(n_1076)
);

XNOR2x1_ASAP7_75t_L g1077 ( 
.A(n_1076),
.B(n_1073),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1077),
.B(n_1075),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_1074),
.B(n_201),
.Y(n_1079)
);

XNOR2xp5_ASAP7_75t_L g1080 ( 
.A(n_1079),
.B(n_198),
.Y(n_1080)
);

OA22x2_ASAP7_75t_L g1081 ( 
.A1(n_1080),
.A2(n_203),
.B1(n_205),
.B2(n_214),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1081),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_1082)
);


endmodule