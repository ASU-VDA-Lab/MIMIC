module fake_jpeg_21219_n_345 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_19),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_47),
.B1(n_31),
.B2(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_85),
.Y(n_104)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_75),
.Y(n_109)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_93),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_50),
.C(n_51),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_50),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_23),
.B1(n_31),
.B2(n_51),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_33),
.Y(n_118)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_103),
.B1(n_65),
.B2(n_44),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_73),
.B1(n_99),
.B2(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI211xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_22),
.B(n_25),
.C(n_26),
.Y(n_101)
);

HB1xp67_ASAP7_75t_SL g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_19),
.Y(n_129)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_34),
.B(n_26),
.Y(n_106)
);

OR2x2_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_27),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_68),
.B1(n_61),
.B2(n_51),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_135),
.B1(n_113),
.B2(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_132),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_94),
.B1(n_86),
.B2(n_84),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_50),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_126),
.C(n_130),
.Y(n_149)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_121),
.B1(n_103),
.B2(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_27),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_44),
.B1(n_45),
.B2(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_21),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_18),
.B(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_46),
.C(n_63),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_132),
.B1(n_127),
.B2(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_76),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_151),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_74),
.A3(n_29),
.B1(n_45),
.B2(n_22),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_145),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_75),
.B1(n_45),
.B2(n_55),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_58),
.B1(n_63),
.B2(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_153),
.B1(n_116),
.B2(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_88),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_83),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_122),
.B1(n_109),
.B2(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_91),
.B1(n_29),
.B2(n_21),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_38),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_114),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_46),
.C(n_120),
.Y(n_175)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_112),
.B1(n_107),
.B2(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_137),
.B1(n_138),
.B2(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_163),
.B(n_115),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_130),
.B1(n_126),
.B2(n_113),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_170),
.B(n_176),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_185),
.B1(n_161),
.B2(n_158),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_119),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_175),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_25),
.B(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_172),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_150),
.B1(n_143),
.B2(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_174),
.A2(n_39),
.B1(n_35),
.B2(n_41),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_122),
.B(n_20),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_131),
.C(n_46),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_181),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_138),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_39),
.B(n_139),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_114),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_110),
.B1(n_20),
.B2(n_115),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_136),
.B(n_20),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_37),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_24),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_144),
.C(n_139),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_192),
.B(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_170),
.B1(n_167),
.B2(n_164),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_206),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_157),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_100),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_212),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_30),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_167),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_162),
.A2(n_35),
.B1(n_39),
.B2(n_32),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_30),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_0),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_221),
.B(n_219),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_169),
.C(n_176),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_230),
.C(n_237),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_246),
.B(n_195),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_187),
.C(n_185),
.Y(n_230)
);

INVx6_ASAP7_75t_SL g232 ( 
.A(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_196),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_162),
.B(n_37),
.C(n_39),
.D(n_11),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_207),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_204),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_204),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_37),
.C(n_10),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_37),
.C(n_10),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_218),
.C(n_198),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_8),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_0),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_230),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_202),
.B1(n_203),
.B2(n_212),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_256),
.B1(n_231),
.B2(n_229),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_255),
.B1(n_257),
.B2(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_202),
.B1(n_197),
.B2(n_198),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_224),
.A2(n_203),
.B1(n_220),
.B2(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_211),
.C(n_209),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_264),
.C(n_266),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_206),
.C(n_216),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_215),
.C(n_8),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_232),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_231),
.C(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_277),
.C(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_242),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_240),
.C(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_237),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_239),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_238),
.B(n_226),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_244),
.C(n_236),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_246),
.B(n_233),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_246),
.B(n_250),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_262),
.B1(n_255),
.B2(n_260),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_299),
.B1(n_0),
.B2(n_2),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_0),
.Y(n_314)
);

HAxp5_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_257),
.CON(n_295),
.SN(n_295)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_296),
.B(n_273),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_271),
.A2(n_266),
.B1(n_1),
.B2(n_2),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_11),
.C(n_16),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_295),
.B1(n_302),
.B2(n_301),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_275),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_305),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_275),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_276),
.B(n_279),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_309),
.B(n_299),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_282),
.B(n_12),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_314),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_6),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_300),
.C(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_323),
.C(n_12),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_321),
.B1(n_12),
.B2(n_15),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_292),
.B1(n_298),
.B2(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_2),
.C(n_3),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_6),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_303),
.B(n_306),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_333),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_321),
.B(n_14),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_316),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_336),
.B1(n_329),
.B2(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_339),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_330),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_339),
.B(n_328),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_323),
.B(n_332),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_4),
.B(n_5),
.C(n_15),
.Y(n_343)
);

AOI31xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_4),
.A3(n_5),
.B(n_2),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_3),
.B(n_141),
.Y(n_345)
);


endmodule