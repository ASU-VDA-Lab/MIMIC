module real_jpeg_20293_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_2),
.A2(n_3),
.B1(n_39),
.B2(n_58),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_39),
.B1(n_61),
.B2(n_62),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_8),
.B1(n_41),
.B2(n_58),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_41),
.B(n_63),
.C(n_87),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_8),
.A2(n_41),
.B1(n_61),
.B2(n_62),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_9),
.B(n_62),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_10),
.B(n_23),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_35),
.B(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_59),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_37)
);

BUFx3_ASAP7_75t_SL g35 ( 
.A(n_11),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_108),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_107),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_95),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_16),
.B(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_80),
.B2(n_94),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B1(n_31),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_21),
.A2(n_22),
.B1(n_48),
.B2(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_21),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_22),
.A2(n_25),
.B(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_22),
.B(n_41),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_24),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_30),
.A2(n_31),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_30),
.A2(n_31),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_31),
.B(n_88),
.C(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_31),
.B(n_159),
.C(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_32),
.B(n_37),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_34),
.A2(n_35),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_35),
.A2(n_36),
.B(n_41),
.C(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_37),
.B(n_41),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_41),
.B(n_74),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_41),
.A2(n_62),
.B(n_76),
.C(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_45),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_47),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_48),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_50),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_49),
.A2(n_50),
.B1(n_102),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_50),
.B(n_122),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_50),
.B(n_102),
.C(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_53),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_55),
.A2(n_56),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_102),
.C(n_104),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B(n_64),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_59),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_60),
.B(n_67),
.C(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_74),
.B(n_75),
.C(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_75),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_74),
.B1(n_78),
.B2(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_93),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_139),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_130),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_90),
.A2(n_91),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_91),
.B(n_128),
.C(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.C(n_101),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_96),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_99),
.B(n_101),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_102),
.A2(n_104),
.B1(n_154),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_104),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_185),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_181),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_168),
.B(n_180),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_156),
.B(n_167),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_142),
.B(n_155),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_133),
.B(n_141),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_124),
.B(n_132),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_120),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_128),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B(n_131),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_158),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_170),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);


endmodule