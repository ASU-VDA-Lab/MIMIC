module real_jpeg_12794_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_52),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_52),
.B1(n_63),
.B2(n_65),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_142),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_142),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_4),
.A2(n_63),
.B1(n_65),
.B2(n_142),
.Y(n_268)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_6),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_36),
.B1(n_63),
.B2(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_184),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_7),
.A2(n_63),
.B1(n_65),
.B2(n_184),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_163),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_163),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_11),
.B(n_28),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_61),
.C(n_63),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_177),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_11),
.A2(n_85),
.B1(n_88),
.B2(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_11),
.B(n_82),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_14),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_14),
.A2(n_24),
.B1(n_63),
.B2(n_65),
.Y(n_174)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_99),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_99),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_83),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_20),
.A2(n_21),
.B1(n_72),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_41),
.C(n_56),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_22),
.A2(n_70),
.B1(n_103),
.B2(n_113),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_23),
.A2(n_28),
.B1(n_96),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g176 ( 
.A(n_25),
.B(n_177),
.CON(n_176),
.SN(n_176)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_25),
.B(n_31),
.C(n_33),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_97),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_28),
.A2(n_96),
.B1(n_176),
.B2(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_29),
.A2(n_37),
.B1(n_141),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_29),
.A2(n_37),
.B1(n_162),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_30),
.A2(n_32),
.B(n_176),
.C(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g235 ( 
.A(n_32),
.B(n_177),
.CON(n_235),
.SN(n_235)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_32),
.B(n_46),
.C(n_49),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_37),
.A2(n_141),
.B(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_69),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_50),
.B(n_53),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_42),
.A2(n_109),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_42),
.A2(n_47),
.B1(n_180),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_42),
.A2(n_47),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_51),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_43),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_43),
.A2(n_54),
.B(n_110),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_43),
.A2(n_82),
.B1(n_212),
.B2(n_235),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_45),
.A2(n_48),
.B(n_235),
.C(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_47),
.A2(n_81),
.B(n_111),
.Y(n_139)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_49),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_48),
.B(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_69),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_66),
.B(n_67),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_57),
.A2(n_66),
.B1(n_93),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_57),
.A2(n_67),
.B(n_94),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_57),
.A2(n_74),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_57),
.A2(n_66),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_57),
.A2(n_66),
.B1(n_240),
.B2(n_263),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_SL g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_62),
.A2(n_78),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_63),
.Y(n_65)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_65),
.B(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_66),
.A2(n_76),
.B(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_66),
.B(n_177),
.Y(n_276)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_73),
.B(n_79),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_145),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B(n_95),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_95),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_84),
.A2(n_92),
.B1(n_125),
.B2(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_85),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_85),
.A2(n_88),
.B1(n_266),
.B2(n_274),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_85),
.A2(n_136),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_86),
.A2(n_87),
.B1(n_155),
.B2(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_86),
.A2(n_90),
.B(n_157),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_86),
.A2(n_87),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_135),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_88),
.A2(n_133),
.B(n_174),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_88),
.B(n_177),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_92),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_114),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_147),
.B(n_316),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_144),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_120),
.B(n_144),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_127),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_126),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_127),
.A2(n_128),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_140),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_129),
.A2(n_130),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_140),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_309),
.B(n_315),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_195),
.B(n_308),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_185),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_150),
.B(n_185),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_166),
.C(n_168),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_151),
.B(n_166),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_160),
.C(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_158),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_168),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.C(n_181),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_170),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_181),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_187),
.B(n_192),
.C(n_194),
.Y(n_314)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_223),
.B(n_303),
.C(n_307),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_216),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.C(n_209),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_198),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_201),
.C(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_217),
.B(n_221),
.C(n_222),
.Y(n_304)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_297),
.B(n_302),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_252),
.B(n_296),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_242),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_242),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.C(n_238),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_229),
.A2(n_230),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_238),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_248),
.C(n_250),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_290),
.B(n_295),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_280),
.B(n_289),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_269),
.B(n_279),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_264),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_264),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B(n_278),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_287),
.C(n_288),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_314),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);


endmodule