module real_jpeg_13004_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_18),
.B(n_19),
.C(n_25),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_46)
);

NAND2x1_ASAP7_75t_SL g68 ( 
.A(n_7),
.B(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_7),
.B(n_32),
.C(n_55),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_70),
.B(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_59),
.Y(n_71)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_74),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_73),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_63),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_63),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_40),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_27),
.Y(n_16)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_18),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g45 ( 
.A1(n_18),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_21),
.B(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_28),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_22),
.A2(n_23),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_23),
.B(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B(n_36),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_28),
.A2(n_36),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_29),
.B(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_29),
.A2(n_37),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_31),
.B(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2x1_ASAP7_75t_R g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_58),
.B2(n_60),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_57),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_66),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.C(n_69),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_87),
.B(n_105),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B(n_104),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_93),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_99),
.B(n_103),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);


endmodule