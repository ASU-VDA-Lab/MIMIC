module fake_jpeg_29054_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_27),
.B(n_9),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_64),
.Y(n_111)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_9),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_27),
.A2(n_18),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_24),
.Y(n_133)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_27),
.Y(n_68)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_73),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_9),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_25),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_35),
.Y(n_107)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_10),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_100),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_32),
.B1(n_50),
.B2(n_35),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_154),
.B1(n_157),
.B2(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_50),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_124),
.B(n_134),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_40),
.B(n_33),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_73),
.B(n_47),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_47),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_137),
.B(n_143),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_73),
.B(n_32),
.Y(n_143)
);

BUFx12f_ASAP7_75t_SL g145 ( 
.A(n_78),
.Y(n_145)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_24),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_88),
.A2(n_38),
.B1(n_19),
.B2(n_49),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_38),
.A3(n_39),
.B1(n_30),
.B2(n_19),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_69),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_30),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_77),
.A2(n_51),
.B1(n_23),
.B2(n_30),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_81),
.A2(n_51),
.B1(n_23),
.B2(n_30),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_52),
.B(n_43),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_49),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_84),
.A2(n_51),
.B1(n_30),
.B2(n_39),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_102),
.C(n_101),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_174),
.B(n_219),
.C(n_226),
.Y(n_264)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_175),
.Y(n_252)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_176),
.Y(n_259)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_181),
.Y(n_233)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_111),
.A2(n_33),
.B1(n_43),
.B2(n_40),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_218),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_63),
.B1(n_156),
.B2(n_135),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_185),
.A2(n_200),
.B1(n_216),
.B2(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_186),
.B(n_224),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_189),
.Y(n_238)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_197),
.Y(n_255)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_199),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_201),
.B(n_202),
.Y(n_261)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_203),
.B(n_204),
.Y(n_266)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_206),
.Y(n_272)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_106),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_209),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_150),
.B1(n_26),
.B2(n_135),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_26),
.Y(n_209)
);

INVx5_ASAP7_75t_SL g210 ( 
.A(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_211),
.Y(n_275)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_98),
.B1(n_97),
.B2(n_93),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_215),
.B1(n_221),
.B2(n_120),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_26),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_214),
.B(n_120),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_89),
.B1(n_86),
.B2(n_103),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_39),
.B1(n_75),
.B2(n_38),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_217),
.Y(n_277)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_151),
.B(n_79),
.C(n_76),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_222),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_127),
.A2(n_67),
.B1(n_46),
.B2(n_38),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_225),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_150),
.B(n_39),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_157),
.A2(n_26),
.B1(n_39),
.B2(n_34),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx12_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_229),
.A2(n_109),
.B1(n_163),
.B2(n_34),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_232),
.A2(n_237),
.B1(n_243),
.B2(n_251),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_165),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_241),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_187),
.A2(n_165),
.B1(n_117),
.B2(n_148),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_117),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_249),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_208),
.B1(n_171),
.B2(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_246),
.B(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_191),
.B(n_141),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_192),
.B(n_139),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_253),
.B(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_179),
.B(n_123),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_267),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_184),
.B(n_141),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_213),
.B(n_123),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_170),
.B(n_195),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_4),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_226),
.A2(n_163),
.B1(n_131),
.B2(n_46),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_269),
.A2(n_276),
.B1(n_248),
.B2(n_271),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_188),
.A2(n_140),
.B1(n_109),
.B2(n_131),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_202),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_279),
.B1(n_18),
.B2(n_6),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_216),
.A2(n_34),
.B1(n_0),
.B2(n_2),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_188),
.A2(n_210),
.B1(n_223),
.B2(n_211),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_185),
.A2(n_10),
.B(n_1),
.C(n_2),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_280),
.A2(n_4),
.B(n_6),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_205),
.B(n_169),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_308),
.B(n_326),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_222),
.B1(n_218),
.B2(n_197),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_183),
.C(n_198),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_290),
.C(n_300),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g288 ( 
.A(n_240),
.Y(n_288)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_288),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_293),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_229),
.C(n_200),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_251),
.A2(n_190),
.B1(n_180),
.B2(n_221),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_291),
.A2(n_305),
.B1(n_317),
.B2(n_244),
.Y(n_348)
);

INVx11_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_294),
.B(n_302),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_299),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_11),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_11),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_238),
.B(n_0),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_301),
.A2(n_307),
.B(n_310),
.Y(n_364)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_274),
.B(n_11),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_306),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_239),
.A2(n_251),
.B1(n_232),
.B2(n_269),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g308 ( 
.A(n_263),
.B(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_309),
.B(n_311),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_266),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_4),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_314),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_277),
.B1(n_231),
.B2(n_258),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_249),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_316),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_242),
.B(n_7),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_246),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_270),
.B1(n_245),
.B2(n_252),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_13),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_321),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_238),
.B(n_13),
.C(n_15),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_244),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_261),
.B(n_13),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_323),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_272),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_15),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_325),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_15),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_239),
.A2(n_17),
.B(n_18),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_R g327 ( 
.A1(n_280),
.A2(n_17),
.B1(n_18),
.B2(n_250),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_327),
.A2(n_17),
.B1(n_278),
.B2(n_301),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_297),
.A2(n_250),
.B1(n_276),
.B2(n_233),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_329),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_331),
.A2(n_343),
.B(n_281),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_297),
.A2(n_233),
.B1(n_259),
.B2(n_277),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_307),
.A2(n_303),
.B1(n_282),
.B2(n_292),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_303),
.A2(n_259),
.B1(n_272),
.B2(n_255),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_288),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_282),
.A2(n_292),
.B1(n_289),
.B2(n_287),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_337),
.A2(n_340),
.B1(n_342),
.B2(n_355),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_338),
.B(n_316),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_317),
.A2(n_255),
.B1(n_256),
.B2(n_270),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_348),
.B1(n_296),
.B2(n_314),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_290),
.A2(n_256),
.B1(n_230),
.B2(n_260),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_283),
.A2(n_230),
.B1(n_260),
.B2(n_258),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_247),
.B1(n_236),
.B2(n_252),
.Y(n_343)
);

AOI22x1_ASAP7_75t_L g353 ( 
.A1(n_288),
.A2(n_298),
.B1(n_284),
.B2(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_323),
.A2(n_254),
.B1(n_257),
.B2(n_245),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_300),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_306),
.A2(n_254),
.B1(n_257),
.B2(n_247),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_358),
.A2(n_360),
.B1(n_338),
.B2(n_332),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_244),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_363),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_295),
.A2(n_278),
.B1(n_236),
.B2(n_17),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_361),
.A2(n_315),
.B(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_311),
.B(n_295),
.Y(n_363)
);

OAI22x1_ASAP7_75t_SL g369 ( 
.A1(n_353),
.A2(n_298),
.B1(n_308),
.B2(n_301),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_369),
.A2(n_381),
.B1(n_395),
.B2(n_361),
.Y(n_416)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_365),
.Y(n_372)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_365),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_378),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_396),
.B1(n_397),
.B2(n_357),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_377),
.A2(n_391),
.B1(n_392),
.B2(n_399),
.Y(n_421)
);

AOI32xp33_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_326),
.A3(n_299),
.B1(n_312),
.B2(n_320),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_320),
.C(n_309),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_398),
.C(n_374),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_362),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_382),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

AOI32xp33_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_324),
.A3(n_304),
.B1(n_294),
.B2(n_305),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_390),
.B(n_361),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_278),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_359),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_364),
.A2(n_293),
.B(n_302),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_386),
.A2(n_389),
.B(n_366),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_285),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_393),
.B1(n_394),
.B2(n_400),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_364),
.A2(n_293),
.B(n_286),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_281),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_330),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_348),
.A2(n_339),
.B1(n_343),
.B2(n_329),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_352),
.A2(n_333),
.B1(n_345),
.B2(n_328),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_340),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_402),
.B1(n_350),
.B2(n_366),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_349),
.B(n_334),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_407),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_404),
.A2(n_422),
.B1(n_429),
.B2(n_381),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_405),
.B(n_409),
.C(n_411),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_347),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_413),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_342),
.C(n_345),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_347),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_346),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_417),
.C(n_419),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_346),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_341),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_418),
.A2(n_421),
.B(n_428),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_371),
.B(n_349),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_370),
.B(n_341),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_424),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_396),
.A2(n_356),
.B1(n_353),
.B2(n_360),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_370),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_368),
.A2(n_331),
.B1(n_353),
.B2(n_335),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_426),
.A2(n_390),
.B1(n_372),
.B2(n_395),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_431),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_368),
.A2(n_358),
.B1(n_355),
.B2(n_336),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_350),
.C(n_336),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_432),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_399),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_386),
.C(n_391),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_400),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_426),
.A2(n_369),
.B(n_393),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_448),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_436),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_455),
.B1(n_411),
.B2(n_408),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_443),
.B(n_449),
.Y(n_461)
);

BUFx12f_ASAP7_75t_SL g444 ( 
.A(n_415),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_444),
.A2(n_409),
.B(n_432),
.Y(n_467)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_431),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_453),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_414),
.B(n_401),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_451),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_420),
.B(n_392),
.Y(n_453)
);

INVx13_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_454),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_422),
.A2(n_404),
.B1(n_429),
.B2(n_430),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_419),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_457),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_424),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_459),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_417),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_405),
.C(n_412),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_474),
.C(n_481),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_444),
.B(n_407),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_466),
.Y(n_498)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_468),
.A2(n_473),
.B1(n_459),
.B2(n_456),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_403),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_476),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_451),
.B(n_447),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_472),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_458),
.B(n_439),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_437),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_442),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_435),
.B(n_437),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_476),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_450),
.Y(n_480)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_457),
.C(n_455),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_486),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_470),
.A2(n_446),
.B1(n_438),
.B2(n_453),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_485),
.A2(n_468),
.B1(n_464),
.B2(n_465),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_471),
.B(n_439),
.CI(n_440),
.CON(n_486),
.SN(n_486)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_443),
.C(n_445),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_489),
.C(n_493),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_436),
.C(n_448),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_477),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_491),
.B(n_494),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_434),
.C(n_454),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_434),
.C(n_454),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_475),
.C(n_461),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_462),
.A2(n_434),
.B1(n_470),
.B2(n_460),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_496),
.A2(n_464),
.B1(n_460),
.B2(n_478),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_479),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_500),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_461),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_502),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_490),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_505),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_483),
.A2(n_480),
.B(n_465),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_509),
.C(n_510),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_475),
.C(n_471),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_467),
.C(n_497),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_490),
.B(n_498),
.Y(n_511)
);

OAI321xp33_ASAP7_75t_L g512 ( 
.A1(n_486),
.A2(n_492),
.A3(n_491),
.B1(n_494),
.B2(n_485),
.C(n_493),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_486),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_515),
.A2(n_503),
.B1(n_514),
.B2(n_516),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_507),
.Y(n_516)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_510),
.C(n_488),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_521),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_495),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_482),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_506),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_524),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_515),
.B(n_492),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_528),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_513),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_517),
.C(n_519),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_530),
.B(n_531),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_524),
.B(n_509),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_532),
.B(n_505),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_527),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_535),
.B(n_533),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_529),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_499),
.B(n_520),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_534),
.C(n_520),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_500),
.C(n_483),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_502),
.C(n_482),
.Y(n_541)
);


endmodule