module fake_jpeg_4359_n_78 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_24),
.A2(n_14),
.B1(n_5),
.B2(n_7),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_4),
.B1(n_5),
.B2(n_26),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_51),
.B(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR4xp25_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_4),
.C(n_52),
.D(n_27),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_31),
.B(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_59),
.C(n_31),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_53),
.C(n_60),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_30),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_74),
.B1(n_67),
.B2(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_32),
.B1(n_48),
.B2(n_44),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_32),
.Y(n_78)
);


endmodule