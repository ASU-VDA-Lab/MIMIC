module real_jpeg_30308_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_1),
.Y(n_543)
);

CKINVDCx11_ASAP7_75t_R g545 ( 
.A(n_1),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_2),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_2),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_2),
.A2(n_289),
.B1(n_360),
.B2(n_363),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_2),
.A2(n_289),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_2),
.A2(n_289),
.B1(n_496),
.B2(n_498),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_30),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_5),
.A2(n_30),
.B1(n_248),
.B2(n_251),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_5),
.A2(n_30),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_6),
.Y(n_273)
);

OAI22x1_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_7),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_95),
.B1(n_119),
.B2(n_122),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_7),
.A2(n_95),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_7),
.B(n_443),
.Y(n_442)
);

OAI32xp33_ASAP7_75t_L g475 ( 
.A1(n_7),
.A2(n_476),
.A3(n_478),
.B1(n_480),
.B2(n_485),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_7),
.B(n_105),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_8),
.B(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_13),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_13),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_13),
.A2(n_52),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_13),
.A2(n_52),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_13),
.A2(n_52),
.B1(n_270),
.B2(n_274),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_299),
.B(n_539),
.C(n_544),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_199),
.Y(n_16)
);

AOI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_191),
.B1(n_192),
.B2(n_195),
.C(n_198),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_163),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_152),
.B(n_162),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_20),
.B(n_152),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_20),
.B(n_153),
.C(n_159),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_20),
.A2(n_152),
.B(n_162),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.C(n_101),
.Y(n_20)
);

OA21x2_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_32),
.B(n_45),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_22),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_22),
.A2(n_32),
.B(n_45),
.Y(n_166)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_29),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_29),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_33),
.A2(n_55),
.B(n_184),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2x1p5_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_34),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_34),
.B(n_286),
.Y(n_314)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_37),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_37),
.Y(n_350)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_42),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_42),
.Y(n_366)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_46),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_55),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_47),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_51),
.Y(n_346)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_55),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_55),
.B(n_286),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_58),
.Y(n_293)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_63),
.A2(n_102),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_63),
.B(n_171),
.C(n_181),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_63),
.B(n_390),
.C(n_392),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_63),
.A2(n_168),
.B1(n_390),
.B2(n_402),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_76),
.B(n_90),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_64),
.B(n_90),
.Y(n_211)
);

NAND2x1_ASAP7_75t_L g254 ( 
.A(n_64),
.B(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_64),
.B(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_64),
.B(n_449),
.Y(n_463)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_R g516 ( 
.A(n_65),
.B(n_95),
.Y(n_516)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_68),
.Y(n_488)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_71),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_71),
.Y(n_322)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_75),
.Y(n_244)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_75),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_75),
.Y(n_484)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_75),
.Y(n_497)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_75),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_76),
.B(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_76),
.B(n_90),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_76),
.B(n_449),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_87),
.Y(n_445)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_87),
.Y(n_453)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_94),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_95),
.A2(n_185),
.B(n_188),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_95),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_95),
.B(n_158),
.Y(n_408)
);

AOI32xp33_ASAP7_75t_L g435 ( 
.A1(n_95),
.A2(n_436),
.A3(n_439),
.B1(n_441),
.B2(n_442),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_95),
.B(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_95),
.B(n_353),
.Y(n_523)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_127),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_104),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_104),
.B(n_358),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_116),
.Y(n_104)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_129),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_105),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_105),
.B(n_359),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_138),
.B(n_144),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_108),
.Y(n_250)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_114),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_137),
.B(n_161),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_117),
.B(n_137),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_R g264 ( 
.A1(n_127),
.A2(n_222),
.B(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_SL g209 ( 
.A(n_128),
.B(n_210),
.C(n_221),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_128),
.B(n_391),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_130),
.A2(n_348),
.B(n_351),
.Y(n_347)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_132),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_132),
.Y(n_362)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp67_ASAP7_75t_L g358 ( 
.A(n_136),
.B(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_138),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_147),
.Y(n_440)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_156),
.B(n_285),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_159),
.B(n_315),
.C(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_160),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.C(n_182),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_165),
.B(n_182),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_171),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_170),
.B(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B(n_179),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_179),
.B(n_358),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_180),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_183),
.B(n_314),
.Y(n_392)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_188),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_SL g199 ( 
.A(n_191),
.B(n_200),
.C(n_202),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_191),
.B(n_200),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_192),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_193),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_225),
.B(n_255),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_196),
.B(n_541),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_197),
.B(n_255),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_258),
.B(n_298),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_203),
.B(n_302),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_256),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_204),
.B(n_256),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_224),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_208),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_209),
.A2(n_210),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_211),
.B(n_448),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_212),
.B(n_267),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_212),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_214),
.B(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_217),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_220),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_225),
.A2(n_226),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_227),
.A2(n_245),
.B1(n_255),
.B2(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_227),
.B(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_227),
.A2(n_255),
.B1(n_434),
.B2(n_435),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_232),
.B(n_240),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_232),
.A2(n_319),
.B(n_326),
.Y(n_318)
);

NAND2x1_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_239),
.Y(n_325)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_241),
.B(n_277),
.Y(n_411)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_245),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_253),
.B(n_254),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_254),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_254),
.B(n_448),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_R g261 ( 
.A(n_262),
.B(n_265),
.C(n_294),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_262),
.A2(n_263),
.B1(n_295),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_265),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_281),
.C(n_284),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_266),
.B(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_268),
.B(n_368),
.Y(n_367)
);

AOI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_277),
.B(n_278),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_327),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_269),
.B(n_277),
.Y(n_354)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_273),
.Y(n_477)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_277),
.B(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_278),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_283),
.Y(n_467)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_295),
.Y(n_423)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_424),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_416),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_380),
.C(n_395),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g416 ( 
.A1(n_308),
.A2(n_417),
.B(n_418),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_369),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_309),
.B(n_369),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_330),
.C(n_367),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_311),
.B(n_367),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_313),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

XOR2x2_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_317),
.B(n_463),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_319),
.A2(n_353),
.B(n_354),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_322),
.Y(n_522)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_326),
.B(n_494),
.Y(n_517)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_328),
.Y(n_512)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_329),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_330),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_355),
.C(n_356),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_352),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_343),
.B(n_347),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_354),
.B(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_357),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_374),
.C(n_376),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_376),
.B1(n_377),
.B2(n_379),
.Y(n_373)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_374),
.Y(n_379)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_393),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_393),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.C(n_388),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_382),
.A2(n_383),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_389),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_390),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_467),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_396),
.B(n_537),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_413),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_398),
.B(n_413),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_406),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_455),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_406),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.C(n_409),
.Y(n_406)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR3xp33_ASAP7_75t_L g535 ( 
.A(n_417),
.B(n_418),
.C(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_419),
.B(n_420),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_535),
.B(n_538),
.Y(n_424)
);

OAI21x1_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_456),
.B(n_534),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_454),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_454),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.C(n_446),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_447),
.Y(n_459)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_447),
.Y(n_446)
);

INVx4_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_470),
.B(n_533),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_460),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.C(n_468),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_466),
.Y(n_531)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_469),
.B(n_531),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_527),
.B(n_532),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_507),
.B(n_526),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_491),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_491),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_489),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_474),
.A2(n_475),
.B1(n_489),
.B2(n_490),
.Y(n_513)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx2_ASAP7_75t_SL g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_502),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_492),
.Y(n_529)
);

AND2x4_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_511),
.Y(n_510)
);

BUFx4f_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_506),
.C(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_514),
.B(n_525),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_513),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_513),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_520),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_512),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_515),
.A2(n_518),
.B(n_524),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_517),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_530),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_SL g539 ( 
.A(n_540),
.B(n_542),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_542),
.B(n_545),
.Y(n_544)
);


endmodule