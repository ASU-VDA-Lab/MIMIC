module fake_aes_11656_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_0), .B(n_2), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
BUFx2_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_1), .Y(n_7) );
INVx1_ASAP7_75t_SL g8 ( .A(n_7), .Y(n_8) );
NAND3xp33_ASAP7_75t_SL g9 ( .A(n_8), .B(n_6), .C(n_5), .Y(n_9) );
NOR3xp33_ASAP7_75t_L g10 ( .A(n_9), .B(n_5), .C(n_2), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
endmodule