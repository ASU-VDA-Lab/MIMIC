module fake_netlist_5_1505_n_4902 (n_924, n_1263, n_977, n_611, n_1126, n_1166, n_469, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_667, n_790, n_1055, n_111, n_880, n_544, n_1007, n_155, n_552, n_1292, n_1198, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_1323, n_688, n_1353, n_800, n_1347, n_671, n_819, n_1022, n_915, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_292, n_625, n_854, n_674, n_417, n_516, n_933, n_1152, n_497, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_1285, n_373, n_307, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_191, n_1104, n_1294, n_659, n_51, n_1257, n_171, n_1182, n_579, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1314, n_709, n_317, n_1236, n_569, n_227, n_920, n_1289, n_94, n_335, n_370, n_976, n_343, n_308, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_1328, n_223, n_264, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_436, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_1267, n_496, n_958, n_1034, n_670, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_395, n_164, n_553, n_901, n_813, n_1284, n_214, n_675, n_888, n_1167, n_637, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_468, n_213, n_129, n_342, n_464, n_363, n_197, n_1069, n_1075, n_1322, n_460, n_889, n_973, n_477, n_571, n_461, n_1211, n_1197, n_907, n_190, n_989, n_1039, n_34, n_228, n_283, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_440, n_793, n_478, n_476, n_534, n_884, n_345, n_944, n_91, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_596, n_558, n_702, n_1276, n_822, n_728, n_266, n_1162, n_272, n_1199, n_352, n_53, n_1038, n_520, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_434, n_868, n_639, n_914, n_411, n_414, n_1293, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_64, n_759, n_28, n_806, n_324, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_367, n_452, n_525, n_1260, n_649, n_547, n_43, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_1308, n_254, n_1233, n_23, n_526, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1008, n_946, n_1001, n_498, n_689, n_738, n_640, n_252, n_624, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1195, n_610, n_936, n_568, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1306, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_456, n_959, n_535, n_152, n_940, n_9, n_592, n_1169, n_45, n_1017, n_123, n_978, n_1054, n_1269, n_1095, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_484, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_374, n_185, n_396, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_723, n_1065, n_1336, n_473, n_1309, n_1043, n_355, n_486, n_614, n_337, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_361, n_700, n_1237, n_573, n_69, n_1132, n_388, n_1300, n_1127, n_761, n_1006, n_329, n_274, n_1270, n_582, n_1332, n_73, n_19, n_309, n_30, n_512, n_84, n_130, n_322, n_1249, n_652, n_1111, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1304, n_1324, n_987, n_261, n_174, n_767, n_993, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_83, n_513, n_1094, n_1354, n_560, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_495, n_602, n_574, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_1327, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1037, n_1080, n_1274, n_1316, n_426, n_1082, n_589, n_716, n_562, n_62, n_952, n_1229, n_391, n_701, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_162, n_960, n_222, n_1290, n_1123, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1029, n_925, n_1206, n_424, n_1311, n_256, n_950, n_380, n_419, n_1346, n_444, n_1299, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_376, n_967, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1357, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_983, n_38, n_280, n_1305, n_873, n_378, n_1112, n_762, n_1283, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1288, n_212, n_385, n_507, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1301, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1329, n_1312, n_804, n_537, n_945, n_492, n_153, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_132, n_1214, n_1342, n_900, n_856, n_918, n_942, n_189, n_1147, n_13, n_1077, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1350, n_1096, n_234, n_833, n_5, n_225, n_1307, n_988, n_814, n_192, n_1201, n_1114, n_655, n_669, n_472, n_1176, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_734, n_638, n_866, n_107, n_969, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_338, n_149, n_693, n_14, n_836, n_990, n_975, n_1256, n_567, n_778, n_1122, n_151, n_306, n_458, n_770, n_1102, n_711, n_85, n_1187, n_1164, n_489, n_1174, n_617, n_1303, n_876, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_172, n_206, n_217, n_726, n_982, n_818, n_861, n_1183, n_899, n_1253, n_210, n_774, n_1335, n_1059, n_1345, n_176, n_1133, n_557, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_393, n_108, n_487, n_665, n_66, n_177, n_421, n_1356, n_910, n_768, n_1302, n_205, n_1136, n_1313, n_754, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_1310, n_202, n_427, n_791, n_732, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_541, n_538, n_1117, n_799, n_687, n_715, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1155, n_89, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_1352, n_626, n_1144, n_1137, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_194, n_855, n_1178, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_780, n_998, n_467, n_1227, n_840, n_1334, n_501, n_823, n_245, n_725, n_1295, n_672, n_581, n_382, n_554, n_898, n_1013, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_997, n_932, n_612, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_737, n_986, n_509, n_1317, n_147, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_733, n_941, n_981, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1108, n_782, n_1100, n_862, n_760, n_381, n_220, n_390, n_1330, n_31, n_481, n_769, n_42, n_1046, n_271, n_934, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_221, n_622, n_1087, n_386, n_994, n_848, n_1223, n_1272, n_104, n_682, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_432, n_839, n_1210, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_78, n_772, n_499, n_517, n_98, n_402, n_413, n_1086, n_796, n_236, n_1012, n_1, n_1348, n_903, n_740, n_203, n_384, n_80, n_35, n_1315, n_277, n_1061, n_92, n_333, n_1298, n_462, n_1193, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_40, n_1028, n_781, n_474, n_542, n_463, n_595, n_502, n_466, n_420, n_1337, n_632, n_699, n_979, n_1245, n_846, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_312, n_1076, n_1091, n_494, n_641, n_730, n_1325, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1220, n_37, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_863, n_805, n_1275, n_113, n_712, n_246, n_1042, n_269, n_285, n_412, n_657, n_644, n_1160, n_491, n_1258, n_1074, n_251, n_160, n_566, n_565, n_597, n_1181, n_1196, n_651, n_1340, n_334, n_811, n_807, n_835, n_175, n_666, n_262, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_166, n_1180, n_1271, n_533, n_1251, n_278, n_4902);

input n_924;
input n_1263;
input n_977;
input n_611;
input n_1126;
input n_1166;
input n_469;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_667;
input n_790;
input n_1055;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1292;
input n_1198;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_688;
input n_1353;
input n_800;
input n_1347;
input n_671;
input n_819;
input n_1022;
input n_915;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_292;
input n_625;
input n_854;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1314;
input n_709;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_1289;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_308;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1328;
input n_223;
input n_264;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_436;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_496;
input n_958;
input n_1034;
input n_670;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1284;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_637;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_197;
input n_1069;
input n_1075;
input n_1322;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_461;
input n_1211;
input n_1197;
input n_907;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_440;
input n_793;
input n_478;
input n_476;
input n_534;
input n_884;
input n_345;
input n_944;
input n_91;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_596;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_434;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1293;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_64;
input n_759;
input n_28;
input n_806;
input n_324;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_649;
input n_547;
input n_43;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_254;
input n_1233;
input n_23;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1008;
input n_946;
input n_1001;
input n_498;
input n_689;
input n_738;
input n_640;
input n_252;
input n_624;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1306;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_9;
input n_592;
input n_1169;
input n_45;
input n_1017;
input n_123;
input n_978;
input n_1054;
input n_1269;
input n_1095;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_484;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_374;
input n_185;
input n_396;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_723;
input n_1065;
input n_1336;
input n_473;
input n_1309;
input n_1043;
input n_355;
input n_486;
input n_614;
input n_337;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1132;
input n_388;
input n_1300;
input n_1127;
input n_761;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_582;
input n_1332;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_84;
input n_130;
input n_322;
input n_1249;
input n_652;
input n_1111;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1304;
input n_1324;
input n_987;
input n_261;
input n_174;
input n_767;
input n_993;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_495;
input n_602;
input n_574;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_426;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_256;
input n_950;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_376;
input n_967;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1357;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_983;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1301;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1329;
input n_1312;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_132;
input n_1214;
input n_1342;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_13;
input n_1077;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1350;
input n_1096;
input n_234;
input n_833;
input n_5;
input n_225;
input n_1307;
input n_988;
input n_814;
input n_192;
input n_1201;
input n_1114;
input n_655;
input n_669;
input n_472;
input n_1176;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_338;
input n_149;
input n_693;
input n_14;
input n_836;
input n_990;
input n_975;
input n_1256;
input n_567;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1102;
input n_711;
input n_85;
input n_1187;
input n_1164;
input n_489;
input n_1174;
input n_617;
input n_1303;
input n_876;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_1253;
input n_210;
input n_774;
input n_1335;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_557;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_393;
input n_108;
input n_487;
input n_665;
input n_66;
input n_177;
input n_421;
input n_1356;
input n_910;
input n_768;
input n_1302;
input n_205;
input n_1136;
input n_1313;
input n_754;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_202;
input n_427;
input n_791;
input n_732;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1155;
input n_89;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1352;
input n_626;
input n_1144;
input n_1137;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_194;
input n_855;
input n_1178;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_780;
input n_998;
input n_467;
input n_1227;
input n_840;
input n_1334;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1295;
input n_672;
input n_581;
input n_382;
input n_554;
input n_898;
input n_1013;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_997;
input n_932;
input n_612;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_737;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_733;
input n_941;
input n_981;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1108;
input n_782;
input n_1100;
input n_862;
input n_760;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_31;
input n_481;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_221;
input n_622;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_432;
input n_839;
input n_1210;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_78;
input n_772;
input n_499;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_236;
input n_1012;
input n_1;
input n_1348;
input n_903;
input n_740;
input n_203;
input n_384;
input n_80;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_1298;
input n_462;
input n_1193;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_40;
input n_1028;
input n_781;
input n_474;
input n_542;
input n_463;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_632;
input n_699;
input n_979;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_312;
input n_1076;
input n_1091;
input n_494;
input n_641;
input n_730;
input n_1325;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1220;
input n_37;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_863;
input n_805;
input n_1275;
input n_113;
input n_712;
input n_246;
input n_1042;
input n_269;
input n_285;
input n_412;
input n_657;
input n_644;
input n_1160;
input n_491;
input n_1258;
input n_1074;
input n_251;
input n_160;
input n_566;
input n_565;
input n_597;
input n_1181;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1251;
input n_278;

output n_4902;

wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_3912;
wire n_1423;
wire n_1729;
wire n_4706;
wire n_2739;
wire n_2380;
wire n_1751;
wire n_2771;
wire n_1508;
wire n_3241;
wire n_4129;
wire n_4604;
wire n_4871;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_4798;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_4419;
wire n_2746;
wire n_1677;
wire n_4477;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_2899;
wire n_2955;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4699;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_1370;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_4577;
wire n_4240;
wire n_4508;
wire n_4854;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_4639;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_3663;
wire n_2487;
wire n_1466;
wire n_1695;
wire n_3766;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4238;
wire n_1451;
wire n_4038;
wire n_2302;
wire n_4109;
wire n_2374;
wire n_1545;
wire n_3341;
wire n_1947;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_4412;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3599;
wire n_3571;
wire n_3785;
wire n_1462;
wire n_2396;
wire n_2069;
wire n_1799;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_4635;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_4013;
wire n_2011;
wire n_2096;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2538;
wire n_2105;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4780;
wire n_3163;
wire n_4425;
wire n_1686;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_2543;
wire n_1860;
wire n_4155;
wire n_1359;
wire n_3695;
wire n_1728;
wire n_2076;
wire n_3036;
wire n_2031;
wire n_2482;
wire n_3891;
wire n_4330;
wire n_4145;
wire n_2677;
wire n_4144;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1705;
wire n_2584;
wire n_4561;
wire n_2639;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_1698;
wire n_3880;
wire n_2329;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_4548;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_3283;
wire n_3048;
wire n_3258;
wire n_4501;
wire n_3937;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_4525;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_4499;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_4816;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_2091;
wire n_1517;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_4691;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_4829;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_4483;
wire n_2149;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_2643;
wire n_4715;
wire n_4793;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_4394;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_4350;
wire n_2384;
wire n_4485;
wire n_4626;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_4468;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_4135;
wire n_2439;
wire n_1931;
wire n_4811;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_1547;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_4615;
wire n_4760;
wire n_4652;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_4624;
wire n_4758;
wire n_3744;
wire n_4263;
wire n_2235;
wire n_1862;
wire n_3980;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_2551;
wire n_1796;
wire n_3291;
wire n_4255;
wire n_4716;
wire n_1473;
wire n_2682;
wire n_1587;
wire n_3755;
wire n_4484;
wire n_2432;
wire n_3668;
wire n_4258;
wire n_1521;
wire n_4498;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_4745;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_4569;
wire n_2506;
wire n_2699;
wire n_4064;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3436;
wire n_1626;
wire n_3542;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_2118;
wire n_2985;
wire n_2944;
wire n_4770;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_4629;
wire n_2932;
wire n_4901;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_3262;
wire n_3136;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_4857;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_4741;
wire n_4861;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_4752;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3837;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_4421;
wire n_2275;
wire n_2855;
wire n_4503;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_4310;
wire n_4836;
wire n_3367;
wire n_4464;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_3096;
wire n_2251;
wire n_1377;
wire n_3915;
wire n_4414;
wire n_2370;
wire n_3496;
wire n_4469;
wire n_3954;
wire n_4114;
wire n_2544;
wire n_4532;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_4067;
wire n_4674;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_4385;
wire n_3320;
wire n_4556;
wire n_3007;
wire n_2688;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_1667;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_4195;
wire n_4218;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4504;
wire n_4375;
wire n_2241;
wire n_4717;
wire n_4788;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_1385;
wire n_2590;
wire n_4815;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_4531;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_4609;
wire n_2987;
wire n_2042;
wire n_1527;
wire n_4567;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_3328;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4471;
wire n_4161;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_2305;
wire n_3392;
wire n_3430;
wire n_3975;
wire n_4444;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_4151;
wire n_4148;
wire n_1883;
wire n_1906;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_4415;
wire n_1387;
wire n_4466;
wire n_3649;
wire n_3528;
wire n_2262;
wire n_4702;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4806;
wire n_4252;
wire n_2322;
wire n_4457;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_4786;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_4160;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_3989;
wire n_4475;
wire n_2837;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_4846;
wire n_1393;
wire n_2319;
wire n_4844;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_4097;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2808;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2679;
wire n_2676;
wire n_1709;
wire n_3981;
wire n_4683;
wire n_2108;
wire n_3640;
wire n_4491;
wire n_4388;
wire n_1538;
wire n_2930;
wire n_4206;
wire n_1838;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_2434;
wire n_1884;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_2967;
wire n_1369;
wire n_3909;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_4886;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_4647;
wire n_3923;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_4696;
wire n_4837;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_2454;
wire n_4371;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_2801;
wire n_3120;
wire n_4473;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_4620;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_2763;
wire n_4613;
wire n_1479;
wire n_1810;
wire n_4480;
wire n_4649;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_4438;
wire n_4876;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_4278;
wire n_4795;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4623;
wire n_4142;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_4553;
wire n_3819;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3978;
wire n_4325;
wire n_4832;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4809;
wire n_4372;
wire n_3500;
wire n_2413;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_2491;
wire n_1788;
wire n_3747;
wire n_1537;
wire n_3833;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_2671;
wire n_4262;
wire n_4184;
wire n_4618;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_4841;
wire n_1798;
wire n_2022;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_4585;
wire n_2876;
wire n_4720;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_2592;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_3484;
wire n_3620;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4842;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_4685;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_4645;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_4490;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_4511;
wire n_2928;
wire n_3128;
wire n_4694;
wire n_1734;
wire n_4533;
wire n_3038;
wire n_4820;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_4757;
wire n_4603;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_4810;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_4648;
wire n_2469;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_4391;
wire n_4641;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_3855;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_2054;
wire n_1503;
wire n_3765;
wire n_1468;
wire n_4638;
wire n_4892;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_3816;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_3113;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_3760;
wire n_4108;
wire n_4486;
wire n_4557;
wire n_4707;
wire n_4078;
wire n_4451;
wire n_1760;
wire n_2875;
wire n_2960;
wire n_1500;
wire n_4527;
wire n_2796;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_4627;
wire n_1851;
wire n_4156;
wire n_3205;
wire n_4848;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_3095;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_4787;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_4541;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_3856;
wire n_2145;
wire n_1639;
wire n_3703;
wire n_4324;
wire n_3030;
wire n_3558;
wire n_4821;
wire n_2580;
wire n_1871;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_3271;
wire n_4771;
wire n_2039;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_4814;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_2084;
wire n_1781;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_4432;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_4855;
wire n_3969;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_2459;
wire n_3031;
wire n_4692;
wire n_4154;
wire n_4619;
wire n_4673;
wire n_3396;
wire n_3701;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_4822;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_4420;
wire n_1773;
wire n_3243;
wire n_1596;
wire n_2666;
wire n_1692;
wire n_2982;
wire n_3385;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_4801;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_4019;
wire n_4826;
wire n_2420;
wire n_2900;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_2339;
wire n_2320;
wire n_2473;
wire n_2038;
wire n_3287;
wire n_4637;
wire n_2137;
wire n_3378;
wire n_4640;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_3767;
wire n_4279;
wire n_4769;
wire n_4785;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_3820;
wire n_4367;
wire n_4589;
wire n_3741;
wire n_3410;
wire n_4578;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_2029;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_4232;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_4413;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_2346;
wire n_2457;
wire n_4387;
wire n_4790;
wire n_2312;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_3015;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_1920;
wire n_1592;
wire n_2536;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_2338;
wire n_1758;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_4847;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_4510;
wire n_4610;
wire n_2571;
wire n_3730;
wire n_3883;
wire n_4489;
wire n_3276;
wire n_2565;
wire n_4152;
wire n_3897;
wire n_3845;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_4570;
wire n_4542;
wire n_2261;
wire n_2156;
wire n_2729;
wire n_1820;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_4447;
wire n_4661;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_2111;
wire n_2521;
wire n_1724;
wire n_3301;
wire n_4285;
wire n_4651;
wire n_3466;
wire n_4534;
wire n_4500;
wire n_3458;
wire n_1420;
wire n_3185;
wire n_3330;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4606;
wire n_4800;
wire n_3960;
wire n_4774;
wire n_2595;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_4597;
wire n_3905;
wire n_4329;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_3586;
wire n_4672;
wire n_3519;
wire n_4433;
wire n_2231;
wire n_1390;
wire n_4682;
wire n_2017;
wire n_2879;
wire n_2474;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_2033;
wire n_1591;
wire n_4071;
wire n_4341;
wire n_4257;
wire n_4766;
wire n_3453;
wire n_1682;
wire n_2628;
wire n_2390;
wire n_1980;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_4460;
wire n_2400;
wire n_4633;
wire n_3645;
wire n_4614;
wire n_3838;
wire n_3223;
wire n_1909;
wire n_3929;
wire n_3077;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_4732;
wire n_2272;
wire n_3984;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_4665;
wire n_1913;
wire n_2878;
wire n_4693;
wire n_1823;
wire n_4434;
wire n_4662;
wire n_3679;
wire n_3779;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_2831;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_4882;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_4744;
wire n_4110;
wire n_2803;
wire n_2851;
wire n_3707;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_4545;
wire n_4868;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_3229;
wire n_4213;
wire n_4463;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_4687;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_4595;
wire n_1849;
wire n_3788;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_2410;
wire n_1961;
wire n_4313;
wire n_4037;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_4802;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_2240;
wire n_2696;
wire n_4063;
wire n_4428;
wire n_4863;
wire n_2436;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3618;
wire n_3592;
wire n_4031;
wire n_4650;
wire n_3525;
wire n_4888;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3995;
wire n_4669;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_4339;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4041;
wire n_2461;
wire n_2858;
wire n_2243;
wire n_4583;
wire n_4060;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_4763;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_4594;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_4666;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3890;
wire n_1611;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_2301;
wire n_3583;
wire n_4494;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_4714;
wire n_3465;
wire n_2419;
wire n_1708;
wire n_3215;
wire n_4796;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_4776;
wire n_4102;
wire n_4891;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_4799;
wire n_1437;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_4807;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_4775;
wire n_3993;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1424;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_4590;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1467;
wire n_4455;
wire n_2053;
wire n_2163;
wire n_4830;
wire n_2328;
wire n_1958;
wire n_4664;
wire n_2254;
wire n_3860;
wire n_1382;
wire n_3546;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3941;
wire n_4754;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_4443;
wire n_3847;
wire n_2664;
wire n_4507;
wire n_4554;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_4575;
wire n_4845;
wire n_3053;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_4663;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3569;
wire n_3548;
wire n_4348;
wire n_4452;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_3953;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_1632;
wire n_3110;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4003;
wire n_3800;
wire n_2402;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_4572;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_4608;
wire n_4840;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_4104;
wire n_4512;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_3749;
wire n_3178;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_4784;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1644;
wire n_4172;
wire n_2334;
wire n_2637;
wire n_4791;
wire n_4384;
wire n_4536;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_4521;
wire n_4488;
wire n_2086;
wire n_3537;
wire n_4423;
wire n_4773;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_2701;
wire n_2783;
wire n_4497;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_4611;
wire n_1763;
wire n_4755;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_4588;
wire n_2475;
wire n_2733;
wire n_2993;
wire n_1719;
wire n_4286;
wire n_3864;
wire n_4598;
wire n_4478;
wire n_2785;
wire n_4658;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_4519;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_4470;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_2499;
wire n_4422;
wire n_4890;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_3417;
wire n_2903;
wire n_3482;
wire n_3921;
wire n_1967;
wire n_3866;
wire n_2233;
wire n_1579;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1439;
wire n_4555;
wire n_4856;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_3326;
wire n_4689;
wire n_3956;
wire n_3572;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4721;
wire n_4047;
wire n_3734;
wire n_3237;
wire n_2082;
wire n_4778;
wire n_2429;
wire n_1992;
wire n_1643;
wire n_1983;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_4550;
wire n_1400;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_4441;
wire n_4496;
wire n_4761;
wire n_3529;
wire n_3854;
wire n_2169;
wire n_1804;
wire n_2468;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_4338;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_4727;
wire n_3952;
wire n_4568;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_4599;
wire n_3633;
wire n_3363;
wire n_4479;
wire n_1373;
wire n_4812;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_2318;
wire n_2393;
wire n_1697;
wire n_1735;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_1881;
wire n_4416;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_2751;
wire n_2707;
wire n_3372;
wire n_3451;
wire n_4539;
wire n_4873;
wire n_2971;
wire n_4657;
wire n_4893;
wire n_3442;
wire n_1549;
wire n_2311;
wire n_1934;
wire n_3950;
wire n_4000;
wire n_4458;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_2298;
wire n_1472;
wire n_2471;
wire n_1807;
wire n_4476;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_4860;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_3342;
wire n_4748;
wire n_2303;
wire n_1824;
wire n_2295;
wire n_1917;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_4667;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_4690;
wire n_1814;
wire n_2822;
wire n_4437;
wire n_4710;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_1848;
wire n_4607;
wire n_2126;
wire n_4547;
wire n_4117;
wire n_2893;
wire n_4573;
wire n_3636;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_4803;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_4668;
wire n_2600;
wire n_4487;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_2795;
wire n_4091;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2282;
wire n_2002;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_4817;
wire n_2371;
wire n_2935;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_4274;
wire n_2098;
wire n_2627;
wire n_3460;
wire n_3409;
wire n_2352;
wire n_4759;
wire n_3538;
wire n_1413;
wire n_4040;
wire n_2207;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_4849;
wire n_4867;
wire n_4474;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2574;
wire n_4728;
wire n_4316;
wire n_3697;
wire n_2361;
wire n_3393;
wire n_1603;
wire n_4247;
wire n_2638;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4887;
wire n_4617;
wire n_4062;
wire n_4524;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_4843;
wire n_2492;
wire n_1998;
wire n_4686;
wire n_4518;
wire n_3759;
wire n_4409;
wire n_4411;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_2034;
wire n_1637;
wire n_1687;
wire n_1419;
wire n_2711;
wire n_4336;
wire n_3933;
wire n_2270;
wire n_1653;
wire n_1506;
wire n_3206;
wire n_4777;
wire n_4792;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_2794;
wire n_2259;
wire n_1702;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_4068;
wire n_4290;
wire n_4253;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_4709;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_4398;
wire n_3155;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1659;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_1834;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_3914;
wire n_4304;
wire n_3911;
wire n_4625;
wire n_2558;
wire n_1371;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_4431;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_3736;
wire n_4656;
wire n_4805;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_4819;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_4885;
wire n_4729;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4900;
wire n_4679;
wire n_4115;
wire n_3174;
wire n_4701;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_2217;
wire n_1453;
wire n_1731;
wire n_3746;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_2745;
wire n_2722;
wire n_2201;
wire n_1737;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_4167;
wire n_2640;
wire n_1993;
wire n_4823;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_4875;
wire n_1777;
wire n_1514;
wire n_1957;
wire n_3967;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_4537;
wire n_3090;
wire n_2067;
wire n_2437;
wire n_2219;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_4730;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_3839;
wire n_1440;
wire n_4631;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_4659;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1774;
wire n_4713;
wire n_1725;
wire n_1491;
wire n_3972;
wire n_4579;
wire n_4616;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_2532;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4747;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1543;
wire n_2224;
wire n_1399;
wire n_1979;
wire n_1991;
wire n_1533;
wire n_3368;
wire n_2924;
wire n_4772;
wire n_3467;
wire n_2484;
wire n_4111;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_4587;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_4743;
wire n_2994;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_4538;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_3928;
wire n_4653;
wire n_4859;
wire n_2692;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_4654;
wire n_2264;
wire n_4677;
wire n_2754;
wire n_3534;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_4632;
wire n_4552;
wire n_2489;
wire n_4275;
wire n_3970;
wire n_3757;
wire n_3438;
wire n_4098;
wire n_2012;
wire n_3792;
wire n_4733;
wire n_4272;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_2245;
wire n_1782;
wire n_3561;
wire n_1418;
wire n_4789;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_2184;
wire n_4695;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_4878;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_3973;
wire n_2814;
wire n_1570;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_4442;
wire n_3968;
wire n_4698;
wire n_4634;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_4704;
wire n_1602;
wire n_2498;
wire n_1461;
wire n_2697;
wire n_4551;
wire n_3074;
wire n_3204;
wire n_4779;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_4072;
wire n_2430;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_4380;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1783;
wire n_4781;
wire n_2977;
wire n_3606;
wire n_4738;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1531;
wire n_4880;
wire n_4424;
wire n_4852;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1388;
wire n_4869;
wire n_1417;
wire n_4700;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_3055;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_4426;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_2817;
wire n_3239;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3172;
wire n_2598;
wire n_4436;
wire n_3878;
wire n_1762;
wire n_4450;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_4601;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_4746;
wire n_1791;
wire n_1890;
wire n_2850;
wire n_1747;
wire n_4220;
wire n_4251;
wire n_1683;
wire n_1944;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_4193;
wire n_4075;
wire n_3982;
wire n_2654;
wire n_3431;
wire n_4621;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_4737;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_4459;
wire n_3176;
wire n_2884;
wire n_2996;
wire n_4351;
wire n_4515;
wire n_2819;
wire n_3126;
wire n_4559;
wire n_4403;
wire n_1981;
wire n_2186;
wire n_1663;
wire n_4368;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_4509;
wire n_4740;
wire n_3609;
wire n_4136;
wire n_4858;
wire n_2315;
wire n_3228;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1952;
wire n_4223;
wire n_4077;
wire n_4642;
wire n_4393;
wire n_2221;
wire n_3576;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_4535;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_4853;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_2326;
wire n_2560;
wire n_3862;
wire n_1569;
wire n_4522;
wire n_2188;
wire n_4794;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_4724;
wire n_4644;
wire n_4456;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_4520;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_2898;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_1861;
wire n_1395;
wire n_3345;
wire n_4546;
wire n_3584;
wire n_1425;
wire n_4592;
wire n_3858;
wire n_4675;
wire n_1901;
wire n_3069;
wire n_4502;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_3691;
wire n_2889;
wire n_4851;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1727;
wire n_1554;
wire n_4382;
wire n_4435;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_4571;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_4764;
wire n_4833;
wire n_3439;
wire n_4889;
wire n_2014;
wire n_3056;
wire n_2345;
wire n_2986;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4723;
wire n_2382;
wire n_4719;
wire n_1707;
wire n_4828;
wire n_4178;
wire n_4655;
wire n_3062;
wire n_3161;
wire n_4581;
wire n_2317;
wire n_3289;
wire n_4558;
wire n_4827;
wire n_2799;
wire n_4454;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_4739;
wire n_2376;
wire n_2488;
wire n_4722;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_4768;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_2778;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_4782;
wire n_1716;
wire n_2788;
wire n_4838;
wire n_2872;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_4363;
wire n_4879;
wire n_4864;
wire n_2691;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_1550;
wire n_4465;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_4605;
wire n_3302;
wire n_4877;
wire n_3235;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_4808;
wire n_1648;
wire n_4015;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4482;
wire n_4865;
wire n_4153;
wire n_2041;
wire n_4564;
wire n_3627;
wire n_3840;
wire n_4300;
wire n_1478;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_3903;
wire n_4783;
wire n_4834;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_4530;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_2173;
wire n_3865;
wire n_3722;
wire n_3859;
wire n_4171;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_4526;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_4417;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_3428;
wire n_2961;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_4899;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_2030;
wire n_2453;
wire n_2883;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_3115;
wire n_4287;
wire n_4749;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_2234;
wire n_4825;
wire n_3251;
wire n_4440;
wire n_4549;
wire n_4804;
wire n_1910;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_4516;
wire n_2209;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4270;
wire n_4505;
wire n_2797;
wire n_1676;
wire n_3118;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_4574;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_4839;
wire n_3497;
wire n_4602;
wire n_1487;
wire n_4449;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_4750;
wire n_1495;
wire n_4445;
wire n_4566;
wire n_4231;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_4576;
wire n_3652;
wire n_4870;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_3114;
wire n_2594;
wire n_3125;
wire n_3234;
wire n_2394;
wire n_4461;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_4835;
wire n_4430;
wire n_2381;
wire n_4767;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_4407;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4676;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_4544;
wire n_4894;
wire n_2170;
wire n_2823;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_3267;
wire n_1595;
wire n_4897;
wire n_2161;
wire n_4429;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_4591;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_4646;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4446;
wire n_4185;
wire n_2642;
wire n_2500;
wire n_4797;
wire n_2366;
wire n_4563;
wire n_4725;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_3247;
wire n_3997;
wire n_2513;
wire n_2525;
wire n_1604;
wire n_3091;
wire n_4831;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4343;
wire n_4319;
wire n_1493;
wire n_4212;
wire n_4320;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_4881;
wire n_4314;
wire n_4596;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_4492;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_3694;
wire n_2586;
wire n_1448;
wire n_4364;
wire n_4288;
wire n_4245;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_4378;
wire n_4726;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_1879;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_4751;
wire n_1505;
wire n_4216;
wire n_4222;
wire n_1634;
wire n_3939;
wire n_4012;
wire n_2019;
wire n_4636;
wire n_2274;
wire n_2972;
wire n_1558;
wire n_3225;
wire n_4584;
wire n_4241;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_4711;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_4680;
wire n_2109;
wire n_2044;
wire n_2013;
wire n_2689;
wire n_1990;
wire n_2920;
wire n_3259;
wire n_4265;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_4560;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_4884;
wire n_3699;
wire n_1827;
wire n_4671;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_3693;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_4705;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;
wire n_4580;

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_612),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_665),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_866),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1328),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_297),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1275),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_816),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1072),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1162),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1310),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_551),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1125),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1064),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_426),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_449),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_710),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_294),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_966),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_783),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_561),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_494),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_34),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_443),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_619),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_43),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_884),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1330),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1115),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_701),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1323),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_442),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_496),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1304),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_391),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1231),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_958),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1317),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_476),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_584),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1237),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_440),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_682),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_733),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_92),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1083),
.Y(n_1403)
);

INVxp33_ASAP7_75t_R g1404 ( 
.A(n_350),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_906),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_911),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1200),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1040),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_771),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_150),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_650),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_918),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1338),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_433),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_931),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_365),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1249),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_364),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_844),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1224),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1287),
.Y(n_1421)
);

BUFx10_ASAP7_75t_L g1422 ( 
.A(n_1290),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_123),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_238),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_691),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_35),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_403),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1340),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_636),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_485),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1202),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_195),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_637),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_460),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1082),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_731),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_703),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_669),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_234),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_921),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_973),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1136),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1321),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1331),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_358),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_876),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_140),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1345),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_569),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_970),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1081),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_18),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_293),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_846),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1327),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_420),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1288),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1156),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_320),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1295),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_183),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_824),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_26),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_697),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_483),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_108),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_885),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_671),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1187),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_750),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1333),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_916),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_604),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_169),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1011),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_853),
.Y(n_1476)
);

BUFx10_ASAP7_75t_L g1477 ( 
.A(n_985),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_79),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_5),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1336),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_728),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_666),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_601),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_95),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_294),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_124),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1013),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1086),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_142),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_983),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1173),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_705),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1265),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1281),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_104),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_605),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_672),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1305),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_548),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_667),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1028),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_81),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1320),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_755),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_584),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_723),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_845),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_725),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_154),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_542),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_842),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1222),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_78),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_607),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1289),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_420),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1343),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_301),
.Y(n_1518)
);

CKINVDCx14_ASAP7_75t_R g1519 ( 
.A(n_305),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1302),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_235),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_258),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_715),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_960),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1141),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_686),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_334),
.Y(n_1527)
);

BUFx8_ASAP7_75t_SL g1528 ( 
.A(n_689),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1352),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_240),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_901),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1088),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_446),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1307),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_832),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_440),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_667),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_897),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1248),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1068),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1241),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1316),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_799),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_718),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_412),
.Y(n_1545)
);

BUFx10_ASAP7_75t_L g1546 ( 
.A(n_1036),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1245),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1020),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_336),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_476),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_849),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_746),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1032),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_708),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_653),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1143),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_16),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1201),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1092),
.Y(n_1559)
);

CKINVDCx16_ASAP7_75t_R g1560 ( 
.A(n_1152),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_325),
.Y(n_1561)
);

BUFx10_ASAP7_75t_L g1562 ( 
.A(n_269),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_706),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_345),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_712),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_570),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1292),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_674),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_92),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_260),
.Y(n_1570)
);

BUFx10_ASAP7_75t_L g1571 ( 
.A(n_1045),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_34),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_681),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_176),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_346),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1108),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_767),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_459),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_790),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1007),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_676),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_927),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_881),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_398),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1144),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_571),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_720),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_873),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_732),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1354),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_329),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_618),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_328),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_452),
.Y(n_1594)
);

BUFx5_ASAP7_75t_L g1595 ( 
.A(n_427),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_415),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1299),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_708),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_681),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_604),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_665),
.Y(n_1601)
);

CKINVDCx16_ASAP7_75t_R g1602 ( 
.A(n_625),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1100),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_811),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_283),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_347),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_682),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_51),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_331),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1116),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_834),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_300),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_670),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1319),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_673),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_722),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_744),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_84),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_364),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_507),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_719),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1257),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1300),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_734),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1058),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_315),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1091),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_124),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_574),
.Y(n_1630)
);

BUFx10_ASAP7_75t_L g1631 ( 
.A(n_647),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_965),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_64),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_695),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_900),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1221),
.Y(n_1636)
);

BUFx5_ASAP7_75t_L g1637 ( 
.A(n_638),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_113),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_208),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_726),
.Y(n_1640)
);

BUFx2_ASAP7_75t_SL g1641 ( 
.A(n_336),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_817),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1104),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_687),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_102),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_143),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_349),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_451),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_634),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_510),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_265),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_629),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1284),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_659),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1066),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1337),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_437),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_886),
.Y(n_1658)
);

CKINVDCx16_ASAP7_75t_R g1659 ( 
.A(n_303),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_422),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_28),
.Y(n_1661)
);

BUFx5_ASAP7_75t_L g1662 ( 
.A(n_167),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_407),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_510),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1301),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_678),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_617),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_205),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_27),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_134),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_150),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_541),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_869),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1314),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_457),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_567),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_321),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_152),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_629),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_625),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_497),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_977),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1075),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_778),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1230),
.Y(n_1685)
);

BUFx10_ASAP7_75t_L g1686 ( 
.A(n_1326),
.Y(n_1686)
);

BUFx10_ASAP7_75t_L g1687 ( 
.A(n_1348),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1087),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_265),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_214),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_378),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_699),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1329),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1324),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_12),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_62),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1286),
.Y(n_1697)
);

CKINVDCx14_ASAP7_75t_R g1698 ( 
.A(n_262),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_992),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_766),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_703),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_540),
.Y(n_1702)
);

BUFx10_ASAP7_75t_L g1703 ( 
.A(n_1318),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_716),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_445),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1151),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1121),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_201),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_548),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1132),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_942),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_692),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1357),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_930),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_630),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1054),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_154),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1306),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_88),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_69),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_529),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_441),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_979),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1255),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_635),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_991),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_630),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1026),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_764),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_377),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_137),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_702),
.Y(n_1732)
);

CKINVDCx20_ASAP7_75t_R g1733 ( 
.A(n_827),
.Y(n_1733)
);

CKINVDCx20_ASAP7_75t_R g1734 ( 
.A(n_724),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_978),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_694),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1065),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1128),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1234),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_558),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_923),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_542),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1315),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1178),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_874),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_309),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_882),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1235),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1350),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_913),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_166),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_239),
.Y(n_1752)
);

BUFx10_ASAP7_75t_L g1753 ( 
.A(n_1262),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_81),
.Y(n_1754)
);

BUFx10_ASAP7_75t_L g1755 ( 
.A(n_281),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1272),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_358),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_250),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_228),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_486),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_627),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1166),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_552),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_306),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_293),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_941),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1096),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1313),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_605),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_717),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_870),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_310),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_489),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_431),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_280),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_247),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1015),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_599),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_506),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_392),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_290),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_288),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_138),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1090),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_238),
.Y(n_1785)
);

BUFx10_ASAP7_75t_L g1786 ( 
.A(n_113),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_212),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_956),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_868),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_518),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1171),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1311),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1349),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_677),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_684),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_362),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1182),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_585),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_700),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_934),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_925),
.Y(n_1801)
);

BUFx10_ASAP7_75t_L g1802 ( 
.A(n_65),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1283),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_728),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_23),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_292),
.Y(n_1806)
);

CKINVDCx16_ASAP7_75t_R g1807 ( 
.A(n_21),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1043),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_745),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_729),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_713),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1027),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1308),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1341),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_512),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1000),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_356),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_266),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1029),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_441),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1062),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_658),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_319),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1332),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_444),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_79),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_789),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_182),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1296),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1334),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_329),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_560),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_371),
.Y(n_1833)
);

BUFx10_ASAP7_75t_L g1834 ( 
.A(n_88),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_591),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1118),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_946),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1344),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_411),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_351),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_902),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_354),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_98),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_707),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_920),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_802),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_46),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_686),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_203),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_67),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_19),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_675),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_679),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_928),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_18),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_458),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1347),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_322),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_939),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_685),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_735),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_413),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_401),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_402),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1037),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_666),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_5),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1033),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_141),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_696),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_696),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_984),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_796),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1285),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1322),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_756),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_475),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_688),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_567),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_591),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_356),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_668),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_535),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_610),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_352),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1303),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_680),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_349),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_831),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_3),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_288),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_12),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_711),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_89),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_819),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1312),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_190),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1291),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_178),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_194),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_341),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1207),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_963),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_286),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_230),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_467),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1212),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_676),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_513),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_883),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_289),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1335),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_601),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_700),
.Y(n_1914)
);

CKINVDCx20_ASAP7_75t_R g1915 ( 
.A(n_683),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_310),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_343),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_971),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1227),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_2),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_835),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1176),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_557),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_709),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_207),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_546),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1069),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1220),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_353),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_944),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_393),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_684),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_209),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_28),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_112),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_218),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_205),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_210),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_375),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_808),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_343),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_839),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_540),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_779),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_908),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1298),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_776),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_144),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_49),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_668),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_71),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1078),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_417),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1080),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1005),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_610),
.Y(n_1956)
);

BUFx8_ASAP7_75t_SL g1957 ( 
.A(n_638),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_653),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_457),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_436),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1353),
.Y(n_1961)
);

INVx2_ASAP7_75t_SL g1962 ( 
.A(n_27),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_843),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_714),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1294),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_721),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_472),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1358),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1325),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_704),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_312),
.Y(n_1971)
);

BUFx10_ASAP7_75t_L g1972 ( 
.A(n_720),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_277),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1071),
.Y(n_1974)
);

CKINVDCx16_ASAP7_75t_R g1975 ( 
.A(n_210),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_416),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1084),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1309),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1351),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1022),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_698),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_35),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1051),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_118),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_153),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_313),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_53),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_171),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_693),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_673),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1183),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_507),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_547),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_533),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_258),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1105),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_19),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_275),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_142),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_741),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_622),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1297),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_103),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_753),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_354),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_773),
.Y(n_2006)
);

BUFx10_ASAP7_75t_L g2007 ( 
.A(n_348),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_324),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1145),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_235),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_348),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_969),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_564),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_495),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_727),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_840),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1196),
.Y(n_2017)
);

CKINVDCx16_ASAP7_75t_R g2018 ( 
.A(n_730),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1010),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_177),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_372),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_211),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_426),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_286),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1293),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_690),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_571),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_654),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_21),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_863),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_312),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1228),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1595),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1595),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1595),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1528),
.Y(n_2036)
);

BUFx2_ASAP7_75t_L g2037 ( 
.A(n_1957),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_1362),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_2018),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1595),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1595),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1637),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1637),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1637),
.Y(n_2044)
);

CKINVDCx16_ASAP7_75t_R g2045 ( 
.A(n_1602),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1364),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1637),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1637),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1662),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1365),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1662),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1502),
.Y(n_2052)
);

CKINVDCx20_ASAP7_75t_R g2053 ( 
.A(n_1395),
.Y(n_2053)
);

BUFx10_ASAP7_75t_L g2054 ( 
.A(n_1964),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1662),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1662),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1662),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1401),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_1421),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1401),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1401),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1506),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1506),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1366),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1506),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1533),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1659),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1533),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1533),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1654),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1654),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_1435),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1654),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1725),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1361),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_1441),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1361),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_1367),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1722),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1725),
.Y(n_2080)
);

CKINVDCx16_ASAP7_75t_R g2081 ( 
.A(n_1779),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_1982),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1807),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_1446),
.Y(n_2084)
);

INVxp33_ASAP7_75t_L g2085 ( 
.A(n_1372),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1725),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1975),
.Y(n_2087)
);

INVxp33_ASAP7_75t_L g2088 ( 
.A(n_1381),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1754),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_1359),
.Y(n_2090)
);

INVxp33_ASAP7_75t_L g2091 ( 
.A(n_1382),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1754),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1368),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1754),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_1519),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1820),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1820),
.Y(n_2097)
);

CKINVDCx20_ASAP7_75t_R g2098 ( 
.A(n_1450),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1820),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1371),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1863),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1422),
.Y(n_2102)
);

INVxp33_ASAP7_75t_SL g2103 ( 
.A(n_1360),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1376),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_1442),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_1374),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1384),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1863),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1385),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1863),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_1386),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1883),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1883),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1424),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1883),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1388),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1920),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1374),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1920),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1920),
.Y(n_2120)
);

CKINVDCx16_ASAP7_75t_R g2121 ( 
.A(n_1560),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2005),
.Y(n_2122)
);

CKINVDCx20_ASAP7_75t_R g2123 ( 
.A(n_1467),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1394),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2005),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2005),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1485),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1598),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_1562),
.Y(n_2129)
);

INVxp33_ASAP7_75t_SL g2130 ( 
.A(n_1363),
.Y(n_2130)
);

CKINVDCx20_ASAP7_75t_R g2131 ( 
.A(n_1475),
.Y(n_2131)
);

INVxp67_ASAP7_75t_SL g2132 ( 
.A(n_1582),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1613),
.Y(n_2133)
);

BUFx2_ASAP7_75t_L g2134 ( 
.A(n_1698),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1622),
.Y(n_2135)
);

BUFx3_ASAP7_75t_L g2136 ( 
.A(n_1422),
.Y(n_2136)
);

BUFx2_ASAP7_75t_SL g2137 ( 
.A(n_1498),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1403),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_SL g2139 ( 
.A(n_1562),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1631),
.Y(n_2140)
);

CKINVDCx20_ASAP7_75t_R g2141 ( 
.A(n_1512),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1407),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1406),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1409),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1625),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1826),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1840),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1415),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2008),
.Y(n_2149)
);

CKINVDCx20_ASAP7_75t_R g2150 ( 
.A(n_1532),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1400),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1420),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1411),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1418),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1430),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_1541),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1440),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1463),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1464),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1473),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1443),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1478),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1444),
.Y(n_2163)
);

CKINVDCx16_ASAP7_75t_R g2164 ( 
.A(n_1623),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1482),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1484),
.Y(n_2166)
);

INVxp33_ASAP7_75t_SL g2167 ( 
.A(n_1369),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1454),
.Y(n_2168)
);

CKINVDCx20_ASAP7_75t_R g2169 ( 
.A(n_1559),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1455),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1458),
.Y(n_2171)
);

CKINVDCx20_ASAP7_75t_R g2172 ( 
.A(n_1580),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1486),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1500),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1549),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_1457),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_1462),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1570),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1575),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1581),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1592),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1601),
.Y(n_2182)
);

CKINVDCx16_ASAP7_75t_R g2183 ( 
.A(n_1750),
.Y(n_2183)
);

CKINVDCx20_ASAP7_75t_R g2184 ( 
.A(n_1585),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1607),
.Y(n_2185)
);

CKINVDCx16_ASAP7_75t_R g2186 ( 
.A(n_1631),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1469),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1470),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1608),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1621),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_1655),
.Y(n_2191)
);

CKINVDCx20_ASAP7_75t_R g2192 ( 
.A(n_1684),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1627),
.Y(n_2193)
);

INVxp67_ASAP7_75t_SL g2194 ( 
.A(n_1624),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1471),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1630),
.Y(n_2196)
);

CKINVDCx20_ASAP7_75t_R g2197 ( 
.A(n_1733),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1634),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1638),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1639),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_1762),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1644),
.Y(n_2202)
);

CKINVDCx20_ASAP7_75t_R g2203 ( 
.A(n_1903),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1476),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1646),
.Y(n_2205)
);

INVxp67_ASAP7_75t_SL g2206 ( 
.A(n_1642),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1648),
.Y(n_2207)
);

CKINVDCx20_ASAP7_75t_R g2208 ( 
.A(n_1912),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1650),
.Y(n_2209)
);

INVxp67_ASAP7_75t_SL g2210 ( 
.A(n_1767),
.Y(n_2210)
);

INVxp33_ASAP7_75t_SL g2211 ( 
.A(n_1375),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_1755),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1480),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1652),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1663),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1667),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_2029),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1670),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1671),
.Y(n_2219)
);

INVxp33_ASAP7_75t_L g2220 ( 
.A(n_1690),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1696),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1704),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1712),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1717),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1487),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_1452),
.Y(n_2226)
);

INVxp33_ASAP7_75t_SL g2227 ( 
.A(n_1378),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1490),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1719),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1491),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1736),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1740),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1757),
.Y(n_2233)
);

CKINVDCx16_ASAP7_75t_R g2234 ( 
.A(n_1755),
.Y(n_2234)
);

CKINVDCx16_ASAP7_75t_R g2235 ( 
.A(n_1786),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2045),
.A2(n_1557),
.B1(n_1647),
.B2(n_1392),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2095),
.B(n_1501),
.Y(n_2237)
);

AND2x6_ASAP7_75t_L g2238 ( 
.A(n_2034),
.B(n_1406),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2058),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2143),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2060),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2061),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2143),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2062),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2046),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2054),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2134),
.B(n_1665),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_2143),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2063),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2050),
.B(n_1714),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2065),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_2075),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2066),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2068),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2039),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_2069),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2070),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_2064),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2071),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2073),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2121),
.A2(n_1947),
.B1(n_1600),
.B2(n_1555),
.Y(n_2261)
);

INVx2_ASAP7_75t_SL g2262 ( 
.A(n_2054),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2078),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2164),
.B(n_1457),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2074),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2217),
.B(n_1683),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2080),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2105),
.A2(n_1456),
.B1(n_1499),
.B2(n_1437),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2086),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2093),
.B(n_2017),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2132),
.B(n_1838),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_2089),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2092),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2094),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2096),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2077),
.B(n_1921),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2097),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2183),
.B(n_1477),
.Y(n_2278)
);

BUFx3_ASAP7_75t_L g2279 ( 
.A(n_2127),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2099),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2102),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_2101),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2108),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2100),
.B(n_1408),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_2103),
.B(n_2130),
.Y(n_2285)
);

INVx5_ASAP7_75t_L g2286 ( 
.A(n_2140),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2136),
.B(n_1534),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_2110),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2112),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2194),
.B(n_1477),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2067),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2113),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2115),
.Y(n_2293)
);

BUFx6f_ASAP7_75t_L g2294 ( 
.A(n_2117),
.Y(n_2294)
);

BUFx2_ASAP7_75t_L g2295 ( 
.A(n_2176),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2119),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2120),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2122),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2079),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2083),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2125),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2126),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2035),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2040),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_2104),
.Y(n_2305)
);

HB1xp67_ASAP7_75t_L g2306 ( 
.A(n_2087),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2033),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2042),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2041),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2043),
.Y(n_2310)
);

AND2x2_ASAP7_75t_SL g2311 ( 
.A(n_2081),
.B(n_2037),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2044),
.Y(n_2312)
);

AND2x2_ASAP7_75t_SL g2313 ( 
.A(n_2186),
.B(n_1373),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2107),
.B(n_1520),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2047),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2206),
.B(n_1548),
.Y(n_2316)
);

BUFx6f_ASAP7_75t_L g2317 ( 
.A(n_2155),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2048),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2049),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_2109),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2181),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2051),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2111),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2055),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_2210),
.B(n_1738),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2182),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2056),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2057),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2116),
.B(n_1551),
.Y(n_2329)
);

XOR2xp5_ASAP7_75t_L g2330 ( 
.A(n_2038),
.B(n_2053),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2226),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2151),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2153),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2124),
.B(n_1729),
.Y(n_2334)
);

AND2x6_ASAP7_75t_L g2335 ( 
.A(n_2154),
.B(n_1406),
.Y(n_2335)
);

HB1xp67_ASAP7_75t_L g2336 ( 
.A(n_2106),
.Y(n_2336)
);

NOR2x1_ASAP7_75t_L g2337 ( 
.A(n_2128),
.B(n_1370),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2133),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_2052),
.B(n_1391),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2158),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2159),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2160),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2162),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2165),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2166),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2138),
.B(n_1965),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_2082),
.B(n_1393),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2118),
.Y(n_2348)
);

NAND2xp33_ASAP7_75t_L g2349 ( 
.A(n_2142),
.B(n_1379),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2173),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2174),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2135),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2175),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2178),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2179),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2180),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2090),
.B(n_1546),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2114),
.B(n_1546),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2144),
.B(n_1919),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2129),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2185),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_2145),
.Y(n_2362)
);

AOI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2234),
.A2(n_1380),
.B1(n_1389),
.B2(n_1387),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2148),
.B(n_1377),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_2152),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2189),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2212),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2157),
.Y(n_2368)
);

AND2x2_ASAP7_75t_SL g2369 ( 
.A(n_2235),
.B(n_1383),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2190),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_2193),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2196),
.Y(n_2372)
);

INVx6_ASAP7_75t_L g2373 ( 
.A(n_2139),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2161),
.B(n_1944),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2198),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_2163),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2168),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2167),
.A2(n_1396),
.B1(n_1397),
.B2(n_1390),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2199),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2200),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2202),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2170),
.B(n_1398),
.Y(n_2382)
);

CKINVDCx20_ASAP7_75t_R g2383 ( 
.A(n_2059),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2171),
.B(n_1571),
.Y(n_2384)
);

CKINVDCx8_ASAP7_75t_R g2385 ( 
.A(n_2137),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_2177),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2187),
.B(n_1405),
.Y(n_2387)
);

OAI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2211),
.A2(n_1926),
.B1(n_1402),
.B2(n_1410),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2205),
.Y(n_2389)
);

AND3x2_ASAP7_75t_L g2390 ( 
.A(n_2207),
.B(n_1495),
.C(n_1468),
.Y(n_2390)
);

OAI22x1_ASAP7_75t_SL g2391 ( 
.A1(n_2036),
.A2(n_1679),
.B1(n_1734),
.B2(n_1668),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2209),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2188),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2227),
.B(n_1412),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2195),
.B(n_1571),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2214),
.Y(n_2396)
);

AND2x6_ASAP7_75t_L g2397 ( 
.A(n_2233),
.B(n_1577),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2204),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2215),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2213),
.B(n_2225),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_SL g2401 ( 
.A(n_2139),
.B(n_1686),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2216),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2228),
.B(n_1686),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2218),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_2230),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2072),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2243),
.Y(n_2407)
);

NAND3xp33_ASAP7_75t_L g2408 ( 
.A(n_2394),
.B(n_2147),
.C(n_2146),
.Y(n_2408)
);

INVx4_ASAP7_75t_L g2409 ( 
.A(n_2245),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2240),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2307),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2359),
.B(n_1687),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2308),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2248),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2254),
.Y(n_2415)
);

INVx8_ASAP7_75t_L g2416 ( 
.A(n_2258),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2284),
.B(n_2085),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2254),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2333),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2340),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2282),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2237),
.Y(n_2422)
);

CKINVDCx16_ASAP7_75t_R g2423 ( 
.A(n_2331),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2374),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2383),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2344),
.Y(n_2426)
);

INVxp33_ASAP7_75t_L g2427 ( 
.A(n_2255),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2345),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2314),
.B(n_2088),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2282),
.Y(n_2430)
);

BUFx4f_ASAP7_75t_L g2431 ( 
.A(n_2373),
.Y(n_2431)
);

INVx1_ASAP7_75t_SL g2432 ( 
.A(n_2252),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_SL g2433 ( 
.A(n_2311),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2303),
.A2(n_1565),
.B1(n_1593),
.B2(n_1496),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2288),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2332),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2350),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2288),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2263),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2351),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2385),
.Y(n_2441)
);

BUFx4f_ASAP7_75t_L g2442 ( 
.A(n_2332),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2339),
.A2(n_2084),
.B1(n_2098),
.B2(n_2076),
.Y(n_2443)
);

INVxp67_ASAP7_75t_SL g2444 ( 
.A(n_2304),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2329),
.B(n_1493),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2334),
.B(n_1494),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2294),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2294),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2309),
.A2(n_1681),
.B1(n_1720),
.B2(n_1633),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2347),
.B(n_1687),
.Y(n_2450)
);

AOI22xp33_ASAP7_75t_L g2451 ( 
.A1(n_2312),
.A2(n_1763),
.B1(n_1849),
.B2(n_1742),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2354),
.Y(n_2452)
);

INVx2_ASAP7_75t_SL g2453 ( 
.A(n_2357),
.Y(n_2453)
);

INVx3_ASAP7_75t_L g2454 ( 
.A(n_2317),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_2317),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2346),
.B(n_2364),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2253),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2370),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2382),
.B(n_2091),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2257),
.Y(n_2460)
);

INVxp67_ASAP7_75t_L g2461 ( 
.A(n_2336),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2372),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2341),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2260),
.Y(n_2464)
);

INVx2_ASAP7_75t_SL g2465 ( 
.A(n_2358),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2387),
.B(n_2220),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2375),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2269),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2274),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2321),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2286),
.B(n_1703),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_2276),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2275),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2283),
.Y(n_2474)
);

AND2x4_ASAP7_75t_L g2475 ( 
.A(n_2247),
.B(n_2149),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2292),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2286),
.B(n_1703),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2296),
.Y(n_2478)
);

NOR2xp67_ASAP7_75t_L g2479 ( 
.A(n_2305),
.B(n_2320),
.Y(n_2479)
);

INVx5_ASAP7_75t_L g2480 ( 
.A(n_2341),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2268),
.B(n_2221),
.C(n_2219),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2301),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_2321),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2313),
.B(n_1753),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2326),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2326),
.Y(n_2486)
);

NAND3xp33_ASAP7_75t_L g2487 ( 
.A(n_2271),
.B(n_2223),
.C(n_2222),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2239),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2371),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2369),
.B(n_1753),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2241),
.Y(n_2491)
);

INVx5_ASAP7_75t_L g2492 ( 
.A(n_2371),
.Y(n_2492)
);

INVx3_ASAP7_75t_L g2493 ( 
.A(n_2279),
.Y(n_2493)
);

INVx2_ASAP7_75t_SL g2494 ( 
.A(n_2266),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2250),
.B(n_1503),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2379),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2380),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2242),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2244),
.Y(n_2499)
);

INVx4_ASAP7_75t_L g2500 ( 
.A(n_2368),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2270),
.B(n_1504),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2384),
.B(n_1507),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2249),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2389),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_L g2505 ( 
.A(n_2238),
.B(n_1577),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2251),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2395),
.B(n_1515),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2315),
.B(n_1517),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2318),
.B(n_2319),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2265),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2396),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2324),
.B(n_1525),
.Y(n_2512)
);

OAI21xp33_ASAP7_75t_SL g2513 ( 
.A1(n_2290),
.A2(n_1606),
.B(n_1561),
.Y(n_2513)
);

CKINVDCx12_ASAP7_75t_R g2514 ( 
.A(n_2236),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2285),
.B(n_1529),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2267),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2273),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_2377),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2401),
.B(n_1538),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2400),
.B(n_1539),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2316),
.A2(n_1933),
.B1(n_1935),
.B2(n_1870),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2310),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2322),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2277),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2256),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2327),
.Y(n_2526)
);

BUFx2_ASAP7_75t_L g2527 ( 
.A(n_2291),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2299),
.B(n_1554),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2280),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2328),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2342),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2343),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2353),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2281),
.B(n_2224),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2289),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2355),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2356),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2361),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2366),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2378),
.B(n_1540),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2293),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2381),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2297),
.Y(n_2543)
);

INVx2_ASAP7_75t_SL g2544 ( 
.A(n_2287),
.Y(n_2544)
);

INVx8_ASAP7_75t_L g2545 ( 
.A(n_2386),
.Y(n_2545)
);

BUFx4f_ASAP7_75t_L g2546 ( 
.A(n_2335),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2295),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2392),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2399),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2298),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2302),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2393),
.B(n_1542),
.Y(n_2552)
);

INVx4_ASAP7_75t_L g2553 ( 
.A(n_2405),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2259),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2272),
.Y(n_2555)
);

INVx3_ASAP7_75t_L g2556 ( 
.A(n_2338),
.Y(n_2556)
);

CKINVDCx20_ASAP7_75t_R g2557 ( 
.A(n_2406),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2325),
.A2(n_1990),
.B1(n_1950),
.B2(n_1609),
.Y(n_2558)
);

INVx4_ASAP7_75t_L g2559 ( 
.A(n_2323),
.Y(n_2559)
);

NAND2xp33_ASAP7_75t_L g2560 ( 
.A(n_2238),
.B(n_1577),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2402),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2238),
.B(n_1543),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2404),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2352),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2362),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2337),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2390),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2335),
.Y(n_2568)
);

NAND2xp33_ASAP7_75t_SL g2569 ( 
.A(n_2348),
.B(n_1746),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_2300),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_2388),
.A2(n_1752),
.B1(n_1962),
.B2(n_1615),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2335),
.B(n_1547),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2397),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2397),
.B(n_1553),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2397),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2403),
.B(n_2123),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2360),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2367),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2246),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2349),
.B(n_1556),
.Y(n_2580)
);

INVx5_ASAP7_75t_L g2581 ( 
.A(n_2262),
.Y(n_2581)
);

NOR2x1p5_ASAP7_75t_L g2582 ( 
.A(n_2264),
.B(n_1399),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2365),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2376),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2398),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2363),
.B(n_2131),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2306),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2278),
.Y(n_2588)
);

INVx4_ASAP7_75t_L g2589 ( 
.A(n_2330),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2261),
.B(n_2141),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2391),
.Y(n_2591)
);

INVx1_ASAP7_75t_SL g2592 ( 
.A(n_2331),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2237),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2243),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2333),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2333),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2411),
.Y(n_2597)
);

BUFx6f_ASAP7_75t_SL g2598 ( 
.A(n_2441),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_SL g2599 ( 
.A(n_2494),
.B(n_2150),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_2453),
.B(n_2156),
.Y(n_2600)
);

OR2x6_ASAP7_75t_L g2601 ( 
.A(n_2416),
.B(n_1641),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2465),
.B(n_2169),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2456),
.B(n_1413),
.Y(n_2603)
);

OR2x6_ASAP7_75t_L g2604 ( 
.A(n_2416),
.B(n_1764),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2419),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2420),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2459),
.B(n_1417),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2466),
.B(n_1419),
.Y(n_2608)
);

INVx2_ASAP7_75t_SL g2609 ( 
.A(n_2592),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2417),
.B(n_1428),
.Y(n_2610)
);

INVxp67_ASAP7_75t_L g2611 ( 
.A(n_2429),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_SL g2612 ( 
.A(n_2422),
.B(n_2593),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2413),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2588),
.B(n_2172),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2424),
.B(n_2184),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2520),
.B(n_2191),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2561),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_L g2618 ( 
.A(n_2461),
.B(n_2192),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2445),
.B(n_1431),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2581),
.B(n_2436),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2426),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2428),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2457),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2427),
.B(n_2446),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2444),
.B(n_1448),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2571),
.A2(n_1460),
.B1(n_1472),
.B2(n_1451),
.Y(n_2626)
);

AND2x4_ASAP7_75t_SL g2627 ( 
.A(n_2557),
.B(n_2197),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2460),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2436),
.Y(n_2629)
);

INVxp67_ASAP7_75t_L g2630 ( 
.A(n_2528),
.Y(n_2630)
);

NOR2x1p5_ASAP7_75t_L g2631 ( 
.A(n_2579),
.B(n_1414),
.Y(n_2631)
);

AND2x6_ASAP7_75t_SL g2632 ( 
.A(n_2590),
.B(n_1770),
.Y(n_2632)
);

O2A1O1Ixp33_ASAP7_75t_L g2633 ( 
.A1(n_2513),
.A2(n_2540),
.B(n_2509),
.C(n_2440),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2437),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2452),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2495),
.B(n_1488),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2458),
.Y(n_2637)
);

AOI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2569),
.A2(n_1660),
.B1(n_1702),
.B2(n_1620),
.C(n_1596),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2464),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2501),
.B(n_1511),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2462),
.A2(n_1531),
.B1(n_1535),
.B2(n_1524),
.Y(n_2641)
);

NAND3xp33_ASAP7_75t_L g2642 ( 
.A(n_2408),
.B(n_1423),
.C(n_1416),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2468),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2467),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2480),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_2527),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2496),
.B(n_1552),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_SL g2648 ( 
.A(n_2409),
.B(n_2201),
.Y(n_2648)
);

NOR2xp67_ASAP7_75t_SL g2649 ( 
.A(n_2575),
.B(n_1694),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2469),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2515),
.B(n_2203),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2497),
.B(n_1656),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2439),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2596),
.A2(n_2208),
.B1(n_1567),
.B2(n_1576),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2581),
.B(n_1558),
.Y(n_2655)
);

AND2x6_ASAP7_75t_L g2656 ( 
.A(n_2573),
.B(n_1697),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2504),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2511),
.B(n_1699),
.Y(n_2658)
);

INVxp67_ASAP7_75t_L g2659 ( 
.A(n_2534),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2595),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2531),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2463),
.B(n_1579),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2580),
.A2(n_1718),
.B1(n_1735),
.B2(n_1716),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2523),
.B(n_1737),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2473),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2526),
.B(n_1743),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2532),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2530),
.A2(n_1745),
.B1(n_1748),
.B2(n_1747),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2474),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2566),
.B(n_1766),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2476),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2463),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2583),
.B(n_2229),
.Y(n_2673)
);

INVx8_ASAP7_75t_L g2674 ( 
.A(n_2545),
.Y(n_2674)
);

AO221x1_ASAP7_75t_L g2675 ( 
.A1(n_2556),
.A2(n_1756),
.B1(n_1836),
.B2(n_1821),
.C(n_1694),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2533),
.Y(n_2676)
);

OR2x6_ASAP7_75t_L g2677 ( 
.A(n_2545),
.B(n_2584),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2570),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2508),
.B(n_1777),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2484),
.B(n_1404),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2489),
.B(n_1583),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2478),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2490),
.B(n_1708),
.Y(n_2683)
);

NOR2xp67_ASAP7_75t_L g2684 ( 
.A(n_2500),
.B(n_2231),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2412),
.B(n_1760),
.Y(n_2685)
);

AO221x1_ASAP7_75t_L g2686 ( 
.A1(n_2567),
.A2(n_1821),
.B1(n_1836),
.B2(n_1756),
.C(n_1694),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2512),
.B(n_1792),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2536),
.B(n_1800),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2537),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2539),
.B(n_1803),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2450),
.B(n_1880),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2552),
.B(n_1913),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2542),
.B(n_1812),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2487),
.A2(n_1813),
.B1(n_1816),
.B2(n_1814),
.Y(n_2694)
);

INVxp67_ASAP7_75t_L g2695 ( 
.A(n_2577),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2548),
.B(n_1827),
.Y(n_2696)
);

INVxp67_ASAP7_75t_L g2697 ( 
.A(n_2578),
.Y(n_2697)
);

AO221x1_ASAP7_75t_L g2698 ( 
.A1(n_2525),
.A2(n_1836),
.B1(n_1837),
.B2(n_1821),
.C(n_1756),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2549),
.B(n_1830),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2563),
.Y(n_2700)
);

NOR3xp33_ASAP7_75t_SL g2701 ( 
.A(n_2423),
.B(n_1426),
.C(n_1425),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2587),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2488),
.B(n_1841),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2576),
.A2(n_1590),
.B1(n_1597),
.B2(n_1588),
.Y(n_2704)
);

INVxp67_ASAP7_75t_L g2705 ( 
.A(n_2432),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_2475),
.Y(n_2706)
);

INVxp67_ASAP7_75t_L g2707 ( 
.A(n_2547),
.Y(n_2707)
);

INVxp67_ASAP7_75t_L g2708 ( 
.A(n_2586),
.Y(n_2708)
);

INVx2_ASAP7_75t_SL g2709 ( 
.A(n_2485),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2491),
.B(n_1845),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2498),
.B(n_1854),
.Y(n_2711)
);

AOI22xp5_ASAP7_75t_L g2712 ( 
.A1(n_2582),
.A2(n_2502),
.B1(n_2507),
.B2(n_2544),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2499),
.B(n_2503),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2482),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2493),
.B(n_1914),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2481),
.A2(n_1857),
.B1(n_1902),
.B2(n_1859),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2559),
.B(n_1923),
.Y(n_2717)
);

AOI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2506),
.A2(n_1604),
.B1(n_1610),
.B2(n_1603),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2489),
.B(n_1611),
.Y(n_2719)
);

OAI221xp5_ASAP7_75t_L g2720 ( 
.A1(n_2521),
.A2(n_1776),
.B1(n_1785),
.B2(n_1774),
.C(n_1772),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2510),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2442),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2516),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2517),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2524),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2529),
.B(n_1918),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2535),
.B(n_1928),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2585),
.B(n_2479),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2541),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_R g2730 ( 
.A(n_2431),
.B(n_1614),
.Y(n_2730)
);

OAI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2472),
.A2(n_2558),
.B1(n_2562),
.B2(n_2572),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2543),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2550),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2551),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2425),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2522),
.B(n_1617),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2522),
.B(n_1626),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2407),
.B(n_1963),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2594),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2564),
.B(n_1974),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_2538),
.B(n_1628),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2414),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2538),
.B(n_1632),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2415),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2565),
.B(n_1978),
.Y(n_2745)
);

AOI22xp33_ASAP7_75t_L g2746 ( 
.A1(n_2568),
.A2(n_1983),
.B1(n_2012),
.B2(n_2002),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2554),
.B(n_2025),
.Y(n_2747)
);

INVx2_ASAP7_75t_SL g2748 ( 
.A(n_2454),
.Y(n_2748)
);

AOI22xp33_ASAP7_75t_L g2749 ( 
.A1(n_2519),
.A2(n_2030),
.B1(n_2032),
.B2(n_1837),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2418),
.Y(n_2750)
);

BUFx5_ASAP7_75t_L g2751 ( 
.A(n_2480),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2492),
.B(n_1635),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2492),
.B(n_1636),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2555),
.B(n_1643),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2421),
.B(n_1653),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2430),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2435),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2438),
.B(n_1658),
.Y(n_2758)
);

INVx8_ASAP7_75t_L g2759 ( 
.A(n_2433),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2518),
.B(n_1673),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2447),
.B(n_2448),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2455),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2574),
.B(n_1674),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2410),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2553),
.A2(n_1685),
.B1(n_1688),
.B2(n_1682),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2546),
.B(n_1693),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2470),
.B(n_2028),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2483),
.B(n_1427),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2434),
.A2(n_1837),
.B1(n_1798),
.B2(n_1810),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2486),
.B(n_1429),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2449),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_L g2772 ( 
.A(n_2451),
.B(n_1700),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2471),
.B(n_1706),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_L g2774 ( 
.A1(n_2505),
.A2(n_1811),
.B1(n_1817),
.B2(n_1787),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2443),
.B(n_1707),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2560),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2477),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2591),
.A2(n_1832),
.B1(n_1833),
.B2(n_1831),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2589),
.B(n_1710),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2514),
.B(n_1711),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2456),
.B(n_1713),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_SL g2782 ( 
.A(n_2409),
.B(n_1773),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2494),
.B(n_1723),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2411),
.Y(n_2784)
);

INVx8_ASAP7_75t_L g2785 ( 
.A(n_2416),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2456),
.B(n_1724),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2494),
.B(n_1726),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2419),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2459),
.B(n_1432),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2494),
.B(n_1728),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2456),
.A2(n_1741),
.B1(n_1744),
.B2(n_1739),
.Y(n_2791)
);

NAND2xp33_ASAP7_75t_L g2792 ( 
.A(n_2456),
.B(n_1749),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2459),
.B(n_1433),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2456),
.B(n_1768),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2456),
.B(n_1771),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2419),
.Y(n_2796)
);

AND3x1_ASAP7_75t_L g2797 ( 
.A(n_2590),
.B(n_1839),
.C(n_1835),
.Y(n_2797)
);

INVx5_ASAP7_75t_L g2798 ( 
.A(n_2436),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2419),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2494),
.B(n_1784),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2494),
.B(n_1788),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2419),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2456),
.B(n_1789),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2456),
.B(n_1791),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2423),
.B(n_2232),
.C(n_1436),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_L g2806 ( 
.A(n_2459),
.B(n_1434),
.Y(n_2806)
);

NOR2x1p5_ASAP7_75t_L g2807 ( 
.A(n_2441),
.B(n_1438),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2459),
.B(n_1439),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2592),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2456),
.B(n_1793),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2459),
.B(n_1445),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2419),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2459),
.B(n_1447),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2411),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2459),
.B(n_1449),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2411),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2411),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2419),
.Y(n_2818)
);

AOI22xp33_ASAP7_75t_L g2819 ( 
.A1(n_2456),
.A2(n_1850),
.B1(n_1851),
.B2(n_1848),
.Y(n_2819)
);

NOR3xp33_ASAP7_75t_L g2820 ( 
.A(n_2423),
.B(n_1459),
.C(n_1453),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2419),
.Y(n_2821)
);

NAND3xp33_ASAP7_75t_L g2822 ( 
.A(n_2459),
.B(n_1465),
.C(n_1461),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_2459),
.B(n_1466),
.Y(n_2823)
);

NOR2xp67_ASAP7_75t_SL g2824 ( 
.A(n_2575),
.B(n_1855),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2419),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2456),
.B(n_1797),
.Y(n_2826)
);

OAI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2456),
.A2(n_1860),
.B1(n_1869),
.B2(n_1844),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2456),
.B(n_1801),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2411),
.Y(n_2829)
);

NAND2xp33_ASAP7_75t_L g2830 ( 
.A(n_2456),
.B(n_1808),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2456),
.B(n_1809),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2411),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_2494),
.B(n_1819),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2456),
.B(n_1824),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2456),
.B(n_1829),
.Y(n_2835)
);

INVxp67_ASAP7_75t_L g2836 ( 
.A(n_2592),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2419),
.Y(n_2837)
);

NAND2xp33_ASAP7_75t_SL g2838 ( 
.A(n_2582),
.B(n_1877),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2597),
.Y(n_2839)
);

AND2x4_ASAP7_75t_L g2840 ( 
.A(n_2609),
.B(n_2809),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2605),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_SL g2842 ( 
.A(n_2653),
.Y(n_2842)
);

OAI22xp5_ASAP7_75t_SL g2843 ( 
.A1(n_2708),
.A2(n_1915),
.B1(n_1916),
.B2(n_1911),
.Y(n_2843)
);

INVx2_ASAP7_75t_SL g2844 ( 
.A(n_2673),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2629),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2613),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_2611),
.B(n_1846),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2789),
.B(n_2793),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2806),
.B(n_1865),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2808),
.A2(n_1970),
.B1(n_1993),
.B2(n_1966),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2781),
.B(n_1868),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2784),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2814),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2606),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_SL g2855 ( 
.A(n_2836),
.B(n_2011),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2705),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2786),
.B(n_1872),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2715),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2811),
.B(n_1873),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2813),
.B(n_2020),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2815),
.B(n_1474),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2823),
.B(n_2794),
.Y(n_2862)
);

INVx2_ASAP7_75t_SL g2863 ( 
.A(n_2702),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2621),
.Y(n_2864)
);

NAND2xp33_ASAP7_75t_L g2865 ( 
.A(n_2751),
.B(n_1874),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2622),
.Y(n_2866)
);

BUFx3_ASAP7_75t_L g2867 ( 
.A(n_2674),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2634),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2627),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2816),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2817),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2829),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2635),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2795),
.B(n_1875),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2637),
.Y(n_2875)
);

HB1xp67_ASAP7_75t_L g2876 ( 
.A(n_2646),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2803),
.B(n_1876),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2672),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2804),
.B(n_1886),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2630),
.B(n_1479),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2798),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2810),
.A2(n_1895),
.B1(n_1896),
.B2(n_1889),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2826),
.B(n_1898),
.Y(n_2883)
);

BUFx4f_ASAP7_75t_L g2884 ( 
.A(n_2674),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2828),
.B(n_1907),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2722),
.B(n_1864),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2831),
.B(n_1910),
.Y(n_2887)
);

NOR3xp33_ASAP7_75t_SL g2888 ( 
.A(n_2827),
.B(n_1483),
.C(n_1481),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2834),
.B(n_1922),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2835),
.B(n_1927),
.Y(n_2890)
);

INVx4_ASAP7_75t_L g2891 ( 
.A(n_2785),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2832),
.Y(n_2892)
);

A2O1A1Ixp33_ASAP7_75t_L g2893 ( 
.A1(n_2692),
.A2(n_1881),
.B(n_1897),
.C(n_1878),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2617),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_R g2895 ( 
.A(n_2648),
.B(n_1930),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2603),
.B(n_1940),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2706),
.B(n_2677),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2785),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2623),
.Y(n_2899)
);

A2O1A1Ixp33_ASAP7_75t_L g2900 ( 
.A1(n_2683),
.A2(n_1905),
.B(n_1909),
.C(n_1899),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2644),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2767),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2657),
.Y(n_2903)
);

INVx1_ASAP7_75t_SL g2904 ( 
.A(n_2735),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2628),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2660),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2610),
.B(n_1942),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2798),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2788),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2607),
.B(n_1945),
.Y(n_2910)
);

A2O1A1Ixp33_ASAP7_75t_L g2911 ( 
.A1(n_2633),
.A2(n_1939),
.B(n_1948),
.C(n_1934),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2624),
.B(n_1946),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2796),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2799),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2608),
.B(n_1952),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2802),
.Y(n_2916)
);

AND3x1_ASAP7_75t_SL g2917 ( 
.A(n_2638),
.B(n_1956),
.C(n_1953),
.Y(n_2917)
);

NAND2x1p5_ASAP7_75t_L g2918 ( 
.A(n_2798),
.B(n_1960),
.Y(n_2918)
);

CKINVDCx5p33_ASAP7_75t_R g2919 ( 
.A(n_2598),
.Y(n_2919)
);

CKINVDCx5p33_ASAP7_75t_R g2920 ( 
.A(n_2677),
.Y(n_2920)
);

OR2x6_ASAP7_75t_L g2921 ( 
.A(n_2759),
.B(n_1981),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2619),
.B(n_1954),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2616),
.A2(n_1961),
.B1(n_1968),
.B2(n_1955),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2812),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2818),
.Y(n_2925)
);

NAND2xp33_ASAP7_75t_L g2926 ( 
.A(n_2751),
.B(n_1969),
.Y(n_2926)
);

INVxp67_ASAP7_75t_L g2927 ( 
.A(n_2717),
.Y(n_2927)
);

OAI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2636),
.A2(n_1979),
.B(n_1977),
.Y(n_2928)
);

AOI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2792),
.A2(n_2830),
.B1(n_2731),
.B2(n_2771),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2651),
.A2(n_1991),
.B1(n_1996),
.B2(n_1980),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2640),
.B(n_2000),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2821),
.A2(n_1987),
.B1(n_1989),
.B2(n_1986),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2707),
.B(n_1998),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2825),
.B(n_2837),
.Y(n_2934)
);

BUFx12f_ASAP7_75t_L g2935 ( 
.A(n_2601),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2639),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2661),
.Y(n_2937)
);

INVxp67_ASAP7_75t_L g2938 ( 
.A(n_2691),
.Y(n_2938)
);

OR2x2_ASAP7_75t_SL g2939 ( 
.A(n_2780),
.B(n_2010),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2667),
.Y(n_2940)
);

NOR3xp33_ASAP7_75t_SL g2941 ( 
.A(n_2838),
.B(n_1492),
.C(n_1489),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2684),
.B(n_2004),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2643),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2759),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2659),
.B(n_1786),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2782),
.B(n_2006),
.Y(n_2946)
);

AOI21x1_ASAP7_75t_L g2947 ( 
.A1(n_2679),
.A2(n_2015),
.B(n_2014),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2678),
.B(n_1497),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2676),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2689),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2695),
.B(n_1505),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2730),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2700),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2687),
.B(n_2009),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2728),
.B(n_2016),
.Y(n_2955)
);

INVx3_ASAP7_75t_L g2956 ( 
.A(n_2764),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2713),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2625),
.B(n_2019),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2650),
.Y(n_2959)
);

CKINVDCx20_ASAP7_75t_R g2960 ( 
.A(n_2615),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2712),
.B(n_1508),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2665),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2669),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2671),
.Y(n_2964)
);

BUFx2_ASAP7_75t_L g2965 ( 
.A(n_2601),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_SL g2966 ( 
.A1(n_2680),
.A2(n_1834),
.B1(n_1972),
.B2(n_1802),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2748),
.B(n_1509),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2744),
.Y(n_2968)
);

HB1xp67_ASAP7_75t_L g2969 ( 
.A(n_2697),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2791),
.B(n_1510),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2682),
.B(n_1513),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2604),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2714),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2721),
.B(n_1514),
.Y(n_2974)
);

AO22x1_ASAP7_75t_L g2975 ( 
.A1(n_2685),
.A2(n_1518),
.B1(n_1521),
.B2(n_1516),
.Y(n_2975)
);

AOI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2822),
.A2(n_1523),
.B1(n_1526),
.B2(n_1522),
.Y(n_2976)
);

NAND3xp33_ASAP7_75t_L g2977 ( 
.A(n_2618),
.B(n_1530),
.C(n_1527),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_2701),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2724),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2729),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2632),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2807),
.B(n_1802),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2797),
.B(n_1834),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2723),
.B(n_1536),
.Y(n_2984)
);

CKINVDCx16_ASAP7_75t_R g2985 ( 
.A(n_2604),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2663),
.A2(n_2626),
.B1(n_2716),
.B2(n_2819),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2725),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2762),
.B(n_1537),
.Y(n_2988)
);

A2O1A1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2670),
.A2(n_1545),
.B(n_1550),
.C(n_1544),
.Y(n_2989)
);

OAI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2704),
.A2(n_1599),
.B1(n_1645),
.B2(n_1574),
.Y(n_2990)
);

INVx4_ASAP7_75t_L g2991 ( 
.A(n_2645),
.Y(n_2991)
);

INVx2_ASAP7_75t_SL g2992 ( 
.A(n_2750),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2733),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2734),
.B(n_2732),
.Y(n_2994)
);

INVx1_ASAP7_75t_SL g2995 ( 
.A(n_2599),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2739),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2742),
.Y(n_2997)
);

INVxp67_ASAP7_75t_L g2998 ( 
.A(n_2768),
.Y(n_2998)
);

BUFx2_ASAP7_75t_L g2999 ( 
.A(n_2656),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2756),
.Y(n_3000)
);

AND2x2_ASAP7_75t_SL g3001 ( 
.A(n_2820),
.B(n_1972),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2757),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2647),
.B(n_1563),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2709),
.Y(n_3004)
);

OAI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2763),
.A2(n_2003),
.B(n_2001),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_SL g3006 ( 
.A1(n_2777),
.A2(n_1566),
.B1(n_1568),
.B2(n_1564),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2652),
.B(n_1569),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2779),
.B(n_1572),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2658),
.B(n_1573),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2751),
.B(n_1578),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2703),
.B(n_1584),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2710),
.B(n_1586),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2614),
.A2(n_1589),
.B1(n_1591),
.B2(n_1587),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2612),
.B(n_2007),
.Y(n_3014)
);

INVx5_ASAP7_75t_L g3015 ( 
.A(n_2656),
.Y(n_3015)
);

INVx2_ASAP7_75t_SL g3016 ( 
.A(n_2631),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2761),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2656),
.A2(n_1605),
.B1(n_1612),
.B2(n_1594),
.Y(n_3018)
);

BUFx2_ASAP7_75t_L g3019 ( 
.A(n_2755),
.Y(n_3019)
);

BUFx2_ASAP7_75t_L g3020 ( 
.A(n_2758),
.Y(n_3020)
);

BUFx8_ASAP7_75t_L g3021 ( 
.A(n_2751),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2664),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2711),
.B(n_1616),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2776),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2726),
.B(n_1618),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2727),
.B(n_1619),
.Y(n_3026)
);

INVx2_ASAP7_75t_SL g3027 ( 
.A(n_2747),
.Y(n_3027)
);

INVx5_ASAP7_75t_L g3028 ( 
.A(n_2805),
.Y(n_3028)
);

INVx4_ASAP7_75t_L g3029 ( 
.A(n_2620),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2754),
.A2(n_1640),
.B(n_1629),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2738),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2600),
.B(n_1649),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2740),
.B(n_1651),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2666),
.Y(n_3034)
);

AO22x1_ASAP7_75t_L g3035 ( 
.A1(n_2773),
.A2(n_1661),
.B1(n_1664),
.B2(n_1657),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2688),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2642),
.A2(n_2654),
.B(n_2745),
.C(n_2770),
.Y(n_3037)
);

NAND2x1p5_ASAP7_75t_L g3038 ( 
.A(n_2602),
.B(n_736),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2765),
.B(n_1666),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2718),
.B(n_1669),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2775),
.B(n_1994),
.Y(n_3041)
);

INVxp67_ASAP7_75t_L g3042 ( 
.A(n_2783),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2690),
.Y(n_3043)
);

INVx4_ASAP7_75t_L g3044 ( 
.A(n_2824),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2693),
.B(n_1672),
.Y(n_3045)
);

AND2x6_ASAP7_75t_SL g3046 ( 
.A(n_2696),
.B(n_2007),
.Y(n_3046)
);

BUFx3_ASAP7_75t_L g3047 ( 
.A(n_2699),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2833),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2686),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2694),
.A2(n_1676),
.B1(n_1677),
.B2(n_1675),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2641),
.B(n_1678),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2787),
.A2(n_1689),
.B(n_1680),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2746),
.B(n_1691),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2801),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2790),
.Y(n_3055)
);

INVx2_ASAP7_75t_SL g3056 ( 
.A(n_2800),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2720),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2749),
.A2(n_1695),
.B1(n_1701),
.B2(n_1692),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2736),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2760),
.B(n_1705),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2737),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2668),
.B(n_2766),
.Y(n_3062)
);

INVxp67_ASAP7_75t_SL g3063 ( 
.A(n_2741),
.Y(n_3063)
);

NAND2x1p5_ASAP7_75t_L g3064 ( 
.A(n_2662),
.B(n_737),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2675),
.A2(n_1715),
.B1(n_1721),
.B2(n_1709),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2769),
.B(n_1727),
.Y(n_3066)
);

AND2x4_ASAP7_75t_L g3067 ( 
.A(n_2681),
.B(n_1730),
.Y(n_3067)
);

AO22x1_ASAP7_75t_L g3068 ( 
.A1(n_2778),
.A2(n_1732),
.B1(n_1751),
.B2(n_1731),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2655),
.B(n_2719),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2698),
.B(n_1758),
.Y(n_3070)
);

NOR2x2_ASAP7_75t_L g3071 ( 
.A(n_2772),
.B(n_1759),
.Y(n_3071)
);

INVx2_ASAP7_75t_SL g3072 ( 
.A(n_2743),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_SL g3073 ( 
.A1(n_2774),
.A2(n_1765),
.B1(n_1769),
.B2(n_1761),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_2752),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2753),
.B(n_1775),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2649),
.B(n_1778),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2611),
.B(n_1780),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2609),
.B(n_1781),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2605),
.Y(n_3079)
);

NAND2x1p5_ASAP7_75t_L g3080 ( 
.A(n_2798),
.B(n_738),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2605),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2605),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2597),
.Y(n_3083)
);

INVx4_ASAP7_75t_L g3084 ( 
.A(n_2674),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_2609),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2611),
.B(n_1782),
.Y(n_3086)
);

OR2x6_ASAP7_75t_L g3087 ( 
.A(n_2674),
.B(n_0),
.Y(n_3087)
);

INVx4_ASAP7_75t_L g3088 ( 
.A(n_2674),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2611),
.B(n_1783),
.Y(n_3089)
);

BUFx3_ASAP7_75t_L g3090 ( 
.A(n_2702),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_2653),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_R g3092 ( 
.A(n_2653),
.B(n_1790),
.Y(n_3092)
);

HB1xp67_ASAP7_75t_L g3093 ( 
.A(n_2609),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2611),
.B(n_1794),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2611),
.B(n_1795),
.Y(n_3095)
);

NAND3xp33_ASAP7_75t_L g3096 ( 
.A(n_2789),
.B(n_1799),
.C(n_1796),
.Y(n_3096)
);

INVx3_ASAP7_75t_L g3097 ( 
.A(n_2629),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2611),
.B(n_1804),
.Y(n_3098)
);

INVx5_ASAP7_75t_L g3099 ( 
.A(n_2674),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2611),
.B(n_1805),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2605),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2597),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2611),
.B(n_1806),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2611),
.B(n_1815),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_2611),
.B(n_1818),
.Y(n_3105)
);

AO22x1_ASAP7_75t_L g3106 ( 
.A1(n_2683),
.A2(n_1823),
.B1(n_1825),
.B2(n_1822),
.Y(n_3106)
);

O2A1O1Ixp5_ASAP7_75t_L g3107 ( 
.A1(n_2848),
.A2(n_740),
.B(n_742),
.C(n_739),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2862),
.B(n_1828),
.Y(n_3108)
);

AOI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_2860),
.A2(n_1843),
.B1(n_1847),
.B2(n_1842),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2861),
.B(n_1852),
.Y(n_3110)
);

AOI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2849),
.A2(n_747),
.B(n_743),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2986),
.A2(n_1856),
.B1(n_1858),
.B2(n_1853),
.Y(n_3112)
);

INVxp67_ASAP7_75t_L g3113 ( 
.A(n_2856),
.Y(n_3113)
);

INVx3_ASAP7_75t_SL g3114 ( 
.A(n_2842),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2839),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2844),
.B(n_1861),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2841),
.Y(n_3117)
);

AOI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_3008),
.A2(n_1866),
.B1(n_1867),
.B2(n_1862),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2859),
.A2(n_749),
.B(n_748),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_3036),
.A2(n_752),
.B(n_751),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2846),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2881),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2852),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2854),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2864),
.Y(n_3125)
);

NOR2xp67_ASAP7_75t_L g3126 ( 
.A(n_3099),
.B(n_754),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2881),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2866),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2927),
.B(n_1871),
.Y(n_3129)
);

OAI22x1_ASAP7_75t_L g3130 ( 
.A1(n_2938),
.A2(n_1882),
.B1(n_1884),
.B2(n_1879),
.Y(n_3130)
);

O2A1O1Ixp5_ASAP7_75t_L g3131 ( 
.A1(n_2911),
.A2(n_758),
.B(n_759),
.C(n_757),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_2998),
.B(n_1885),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2858),
.B(n_1887),
.Y(n_3133)
);

O2A1O1Ixp33_ASAP7_75t_L g3134 ( 
.A1(n_2900),
.A2(n_2893),
.B(n_2902),
.C(n_2989),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2868),
.Y(n_3135)
);

INVxp67_ASAP7_75t_SL g3136 ( 
.A(n_3093),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2873),
.Y(n_3137)
);

AND2x4_ASAP7_75t_L g3138 ( 
.A(n_3090),
.B(n_760),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_SL g3139 ( 
.A(n_3091),
.B(n_1988),
.Y(n_3139)
);

BUFx8_ASAP7_75t_SL g3140 ( 
.A(n_2944),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_3031),
.A2(n_762),
.B(n_761),
.Y(n_3141)
);

A2O1A1Ixp33_ASAP7_75t_L g3142 ( 
.A1(n_2929),
.A2(n_1890),
.B(n_1891),
.C(n_1888),
.Y(n_3142)
);

INVxp67_ASAP7_75t_L g3143 ( 
.A(n_2840),
.Y(n_3143)
);

O2A1O1Ixp5_ASAP7_75t_L g3144 ( 
.A1(n_2851),
.A2(n_765),
.B(n_768),
.C(n_763),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2957),
.B(n_1892),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2877),
.A2(n_770),
.B(n_769),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_3042),
.A2(n_1894),
.B1(n_1900),
.B2(n_1893),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2883),
.A2(n_774),
.B(n_772),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_3022),
.B(n_1901),
.Y(n_3149)
);

O2A1O1Ixp33_ASAP7_75t_SL g3150 ( 
.A1(n_3037),
.A2(n_777),
.B(n_780),
.C(n_775),
.Y(n_3150)
);

OR2x2_ASAP7_75t_L g3151 ( 
.A(n_2904),
.B(n_1904),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3034),
.B(n_1906),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2885),
.A2(n_782),
.B(n_781),
.Y(n_3153)
);

O2A1O1Ixp33_ASAP7_75t_L g3154 ( 
.A1(n_3077),
.A2(n_1917),
.B(n_1924),
.C(n_1908),
.Y(n_3154)
);

NAND3xp33_ASAP7_75t_L g3155 ( 
.A(n_2850),
.B(n_1929),
.C(n_1925),
.Y(n_3155)
);

NOR2xp33_ASAP7_75t_L g3156 ( 
.A(n_3089),
.B(n_1931),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2887),
.A2(n_785),
.B(n_784),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2853),
.Y(n_3158)
);

AOI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_3055),
.A2(n_1936),
.B1(n_1937),
.B2(n_1932),
.Y(n_3159)
);

BUFx6f_ASAP7_75t_L g3160 ( 
.A(n_2944),
.Y(n_3160)
);

BUFx3_ASAP7_75t_L g3161 ( 
.A(n_2867),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_3043),
.B(n_1938),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3017),
.B(n_1941),
.Y(n_3163)
);

INVx4_ASAP7_75t_L g3164 ( 
.A(n_3099),
.Y(n_3164)
);

A2O1A1Ixp33_ASAP7_75t_SL g3165 ( 
.A1(n_3060),
.A2(n_787),
.B(n_788),
.C(n_786),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2875),
.Y(n_3166)
);

BUFx6f_ASAP7_75t_L g3167 ( 
.A(n_2908),
.Y(n_3167)
);

AOI33xp33_ASAP7_75t_L g3168 ( 
.A1(n_2966),
.A2(n_1958),
.A3(n_1949),
.B1(n_1959),
.B2(n_1951),
.B3(n_1943),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_3094),
.B(n_1967),
.Y(n_3169)
);

A2O1A1Ixp33_ASAP7_75t_L g3170 ( 
.A1(n_3062),
.A2(n_1973),
.B(n_1976),
.C(n_1971),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2901),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_R g3172 ( 
.A(n_2898),
.B(n_1984),
.Y(n_3172)
);

OAI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_3049),
.A2(n_1992),
.B(n_1985),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_2889),
.A2(n_792),
.B(n_791),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2870),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3047),
.B(n_1995),
.Y(n_3176)
);

AND2x4_ASAP7_75t_L g3177 ( 
.A(n_2891),
.B(n_793),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2934),
.A2(n_795),
.B(n_794),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2903),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_3069),
.A2(n_1999),
.B(n_2013),
.C(n_1997),
.Y(n_3180)
);

A2O1A1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_3048),
.A2(n_2022),
.B(n_2023),
.C(n_2021),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3027),
.B(n_2024),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2871),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_2876),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2906),
.B(n_2909),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_3063),
.A2(n_798),
.B(n_797),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_3024),
.A2(n_2027),
.B1(n_2031),
.B2(n_2026),
.Y(n_3187)
);

NOR2x1_ASAP7_75t_R g3188 ( 
.A(n_3084),
.B(n_0),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2872),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2913),
.B(n_2914),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2857),
.A2(n_801),
.B(n_800),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2916),
.B(n_1),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2924),
.Y(n_3193)
);

HB1xp67_ASAP7_75t_L g3194 ( 
.A(n_3085),
.Y(n_3194)
);

OAI22xp5_ASAP7_75t_L g3195 ( 
.A1(n_3054),
.A2(n_804),
.B1(n_805),
.B2(n_803),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2925),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3079),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3081),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2892),
.Y(n_3199)
);

O2A1O1Ixp5_ASAP7_75t_SL g3200 ( 
.A1(n_2961),
.A2(n_2915),
.B(n_2912),
.C(n_2879),
.Y(n_3200)
);

AOI21x1_ASAP7_75t_L g3201 ( 
.A1(n_2874),
.A2(n_807),
.B(n_806),
.Y(n_3201)
);

A2O1A1Ixp33_ASAP7_75t_L g3202 ( 
.A1(n_3075),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_3202)
);

BUFx3_ASAP7_75t_L g3203 ( 
.A(n_2884),
.Y(n_3203)
);

INVxp67_ASAP7_75t_L g3204 ( 
.A(n_2969),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3082),
.B(n_4),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3056),
.A2(n_810),
.B1(n_812),
.B2(n_809),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3101),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2907),
.B(n_6),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_R g3209 ( 
.A(n_2869),
.B(n_813),
.Y(n_3209)
);

BUFx6f_ASAP7_75t_L g3210 ( 
.A(n_2863),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2890),
.A2(n_815),
.B(n_814),
.Y(n_3211)
);

O2A1O1Ixp33_ASAP7_75t_SL g3212 ( 
.A1(n_3070),
.A2(n_820),
.B(n_821),
.C(n_818),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2896),
.A2(n_823),
.B(n_822),
.Y(n_3213)
);

AOI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_2995),
.A2(n_826),
.B1(n_828),
.B2(n_825),
.Y(n_3214)
);

O2A1O1Ixp33_ASAP7_75t_SL g3215 ( 
.A1(n_2970),
.A2(n_830),
.B(n_833),
.C(n_829),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_2910),
.A2(n_837),
.B1(n_838),
.B2(n_836),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3019),
.B(n_6),
.Y(n_3217)
);

NOR2xp67_ASAP7_75t_SL g3218 ( 
.A(n_3015),
.B(n_7),
.Y(n_3218)
);

NAND2x1p5_ASAP7_75t_L g3219 ( 
.A(n_3088),
.B(n_841),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2994),
.A2(n_848),
.B(n_847),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2958),
.A2(n_851),
.B(n_850),
.Y(n_3221)
);

BUFx2_ASAP7_75t_SL g3222 ( 
.A(n_2897),
.Y(n_3222)
);

OR2x6_ASAP7_75t_L g3223 ( 
.A(n_2935),
.B(n_7),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2894),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_3020),
.A2(n_854),
.B(n_852),
.Y(n_3225)
);

O2A1O1Ixp5_ASAP7_75t_L g3226 ( 
.A1(n_3005),
.A2(n_3010),
.B(n_2928),
.C(n_3044),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2845),
.Y(n_3227)
);

O2A1O1Ixp33_ASAP7_75t_L g3228 ( 
.A1(n_3086),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_3228)
);

INVx3_ASAP7_75t_L g3229 ( 
.A(n_3097),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2886),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_2933),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2937),
.Y(n_3232)
);

NAND2x1_ASAP7_75t_L g3233 ( 
.A(n_2899),
.B(n_855),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_2940),
.A2(n_857),
.B1(n_858),
.B2(n_856),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3057),
.B(n_8),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2949),
.Y(n_3236)
);

BUFx12f_ASAP7_75t_L g3237 ( 
.A(n_2919),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_2960),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_2855),
.B(n_859),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2950),
.B(n_9),
.Y(n_3240)
);

BUFx3_ASAP7_75t_L g3241 ( 
.A(n_3021),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2953),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2991),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_SL g3244 ( 
.A(n_2952),
.B(n_860),
.Y(n_3244)
);

INVx5_ASAP7_75t_L g3245 ( 
.A(n_3087),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2922),
.B(n_2931),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_SL g3247 ( 
.A(n_3096),
.B(n_861),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2954),
.B(n_10),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_3000),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_2865),
.A2(n_864),
.B(n_862),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_2926),
.A2(n_867),
.B(n_865),
.Y(n_3251)
);

INVxp67_ASAP7_75t_L g3252 ( 
.A(n_2945),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3095),
.B(n_11),
.Y(n_3253)
);

AOI221xp5_ASAP7_75t_L g3254 ( 
.A1(n_2843),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.C(n_15),
.Y(n_3254)
);

O2A1O1Ixp33_ASAP7_75t_L g3255 ( 
.A1(n_3098),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_3255)
);

BUFx6f_ASAP7_75t_L g3256 ( 
.A(n_3016),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3100),
.B(n_16),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3103),
.B(n_17),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3059),
.A2(n_872),
.B(n_871),
.Y(n_3259)
);

AO21x2_ASAP7_75t_L g3260 ( 
.A1(n_2955),
.A2(n_3007),
.B(n_3003),
.Y(n_3260)
);

AOI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3061),
.A2(n_877),
.B(n_875),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2996),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_3072),
.A2(n_2977),
.B1(n_2882),
.B2(n_3039),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_SL g3264 ( 
.A(n_3104),
.B(n_878),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2987),
.A2(n_880),
.B(n_879),
.Y(n_3265)
);

A2O1A1Ixp33_ASAP7_75t_SL g3266 ( 
.A1(n_3065),
.A2(n_888),
.B(n_889),
.C(n_887),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2979),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2980),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_SL g3269 ( 
.A1(n_2981),
.A2(n_22),
.B1(n_17),
.B2(n_20),
.Y(n_3269)
);

OAI22xp5_ASAP7_75t_L g3270 ( 
.A1(n_3041),
.A2(n_891),
.B1(n_892),
.B2(n_890),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2997),
.Y(n_3271)
);

NAND3xp33_ASAP7_75t_SL g3272 ( 
.A(n_2895),
.B(n_20),
.C(n_22),
.Y(n_3272)
);

O2A1O1Ixp33_ASAP7_75t_L g3273 ( 
.A1(n_2990),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3273)
);

NOR3xp33_ASAP7_75t_SL g3274 ( 
.A(n_2978),
.B(n_24),
.C(n_25),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2905),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_2993),
.A2(n_894),
.B(n_893),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2936),
.Y(n_3277)
);

INVx5_ASAP7_75t_L g3278 ( 
.A(n_3087),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3009),
.B(n_26),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_2943),
.A2(n_896),
.B(n_895),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2959),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_2880),
.B(n_29),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2962),
.A2(n_899),
.B(n_898),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2963),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_SL g3285 ( 
.A(n_3015),
.B(n_903),
.Y(n_3285)
);

AOI21x1_ASAP7_75t_L g3286 ( 
.A1(n_2964),
.A2(n_905),
.B(n_904),
.Y(n_3286)
);

NOR3xp33_ASAP7_75t_SL g3287 ( 
.A(n_2985),
.B(n_29),
.C(n_30),
.Y(n_3287)
);

CKINVDCx11_ASAP7_75t_R g3288 ( 
.A(n_3046),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2973),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_3105),
.A2(n_2946),
.B(n_2847),
.C(n_3040),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_3083),
.A2(n_909),
.B(n_907),
.Y(n_3291)
);

OAI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3004),
.A2(n_3102),
.B1(n_3045),
.B2(n_3033),
.Y(n_3292)
);

BUFx12f_ASAP7_75t_L g3293 ( 
.A(n_2920),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3011),
.B(n_30),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2971),
.A2(n_912),
.B(n_910),
.Y(n_3295)
);

AND2x4_ASAP7_75t_SL g3296 ( 
.A(n_3029),
.B(n_914),
.Y(n_3296)
);

AND2x4_ASAP7_75t_L g3297 ( 
.A(n_2878),
.B(n_2956),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3028),
.B(n_915),
.Y(n_3298)
);

AOI21x1_ASAP7_75t_L g3299 ( 
.A1(n_2947),
.A2(n_919),
.B(n_917),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3012),
.B(n_31),
.Y(n_3300)
);

BUFx2_ASAP7_75t_L g3301 ( 
.A(n_2972),
.Y(n_3301)
);

AOI21x1_ASAP7_75t_L g3302 ( 
.A1(n_2942),
.A2(n_924),
.B(n_922),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_2951),
.B(n_31),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3002),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2968),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_2992),
.A2(n_3025),
.B1(n_3026),
.B2(n_3023),
.Y(n_3306)
);

INVx4_ASAP7_75t_L g3307 ( 
.A(n_3028),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3246),
.A2(n_2984),
.B(n_2974),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3306),
.A2(n_3038),
.B(n_3074),
.Y(n_3309)
);

OAI22x1_ASAP7_75t_L g3310 ( 
.A1(n_3282),
.A2(n_2983),
.B1(n_3032),
.B2(n_2965),
.Y(n_3310)
);

AOI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_3156),
.A2(n_2948),
.B1(n_2982),
.B2(n_3001),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_3161),
.B(n_2999),
.Y(n_3312)
);

OR2x6_ASAP7_75t_L g3313 ( 
.A(n_3160),
.B(n_3080),
.Y(n_3313)
);

AO31x2_ASAP7_75t_L g3314 ( 
.A1(n_3170),
.A2(n_3030),
.A3(n_3076),
.B(n_3052),
.Y(n_3314)
);

A2O1A1Ixp33_ASAP7_75t_L g3315 ( 
.A1(n_3169),
.A2(n_2888),
.B(n_2941),
.C(n_3006),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3117),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3110),
.A2(n_2930),
.B1(n_2923),
.B2(n_3078),
.Y(n_3317)
);

OAI21x1_ASAP7_75t_L g3318 ( 
.A1(n_3201),
.A2(n_3064),
.B(n_2918),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3226),
.A2(n_3066),
.B(n_3051),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3185),
.A2(n_3190),
.B1(n_3263),
.B2(n_3108),
.Y(n_3320)
);

OAI21x1_ASAP7_75t_L g3321 ( 
.A1(n_3302),
.A2(n_2932),
.B(n_3053),
.Y(n_3321)
);

NAND3x1_ASAP7_75t_L g3322 ( 
.A(n_3254),
.B(n_3013),
.C(n_2976),
.Y(n_3322)
);

A2O1A1Ixp33_ASAP7_75t_L g3323 ( 
.A1(n_3173),
.A2(n_3067),
.B(n_3014),
.C(n_3018),
.Y(n_3323)
);

O2A1O1Ixp5_ASAP7_75t_L g3324 ( 
.A1(n_3208),
.A2(n_3035),
.B(n_3106),
.C(n_2975),
.Y(n_3324)
);

AO31x2_ASAP7_75t_L g3325 ( 
.A1(n_3142),
.A2(n_3058),
.A3(n_2917),
.B(n_3071),
.Y(n_3325)
);

INVx5_ASAP7_75t_L g3326 ( 
.A(n_3140),
.Y(n_3326)
);

NAND2x1p5_ASAP7_75t_L g3327 ( 
.A(n_3210),
.B(n_2967),
.Y(n_3327)
);

OR2x6_ASAP7_75t_L g3328 ( 
.A(n_3160),
.B(n_2921),
.Y(n_3328)
);

OAI21x1_ASAP7_75t_L g3329 ( 
.A1(n_3200),
.A2(n_3286),
.B(n_3299),
.Y(n_3329)
);

INVx3_ASAP7_75t_SL g3330 ( 
.A(n_3114),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3290),
.A2(n_2988),
.B(n_2921),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3124),
.Y(n_3332)
);

OAI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_3248),
.A2(n_3073),
.B(n_3050),
.Y(n_3333)
);

NAND2x1p5_ASAP7_75t_L g3334 ( 
.A(n_3210),
.B(n_3092),
.Y(n_3334)
);

OAI21x1_ASAP7_75t_L g3335 ( 
.A1(n_3233),
.A2(n_3131),
.B(n_3107),
.Y(n_3335)
);

NAND2x1p5_ASAP7_75t_L g3336 ( 
.A(n_3164),
.B(n_2939),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3125),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3145),
.B(n_3068),
.Y(n_3338)
);

AOI21x1_ASAP7_75t_L g3339 ( 
.A1(n_3247),
.A2(n_929),
.B(n_926),
.Y(n_3339)
);

CKINVDCx5p33_ASAP7_75t_R g3340 ( 
.A(n_3237),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_SL g3341 ( 
.A1(n_3250),
.A2(n_933),
.B(n_932),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_3139),
.B(n_32),
.Y(n_3342)
);

OA21x2_ASAP7_75t_L g3343 ( 
.A1(n_3144),
.A2(n_936),
.B(n_935),
.Y(n_3343)
);

O2A1O1Ixp5_ASAP7_75t_SL g3344 ( 
.A1(n_3264),
.A2(n_3298),
.B(n_3239),
.C(n_3216),
.Y(n_3344)
);

CKINVDCx5p33_ASAP7_75t_R g3345 ( 
.A(n_3293),
.Y(n_3345)
);

OAI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3134),
.A2(n_938),
.B(n_937),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3129),
.B(n_32),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3128),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3163),
.B(n_33),
.Y(n_3349)
);

OAI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_3279),
.A2(n_943),
.B(n_940),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3260),
.A2(n_947),
.B(n_945),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3149),
.B(n_33),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3152),
.B(n_36),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3135),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3162),
.B(n_36),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3292),
.A2(n_949),
.B(n_948),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3137),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_L g3358 ( 
.A1(n_3251),
.A2(n_951),
.B(n_950),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_3203),
.B(n_952),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3303),
.B(n_37),
.Y(n_3360)
);

AND2x6_ASAP7_75t_L g3361 ( 
.A(n_3177),
.B(n_953),
.Y(n_3361)
);

AO21x2_ASAP7_75t_L g3362 ( 
.A1(n_3165),
.A2(n_955),
.B(n_954),
.Y(n_3362)
);

INVxp67_ASAP7_75t_SL g3363 ( 
.A(n_3204),
.Y(n_3363)
);

A2O1A1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3253),
.A2(n_3258),
.B(n_3257),
.C(n_3154),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3166),
.B(n_37),
.Y(n_3365)
);

OAI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3294),
.A2(n_959),
.B(n_957),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3133),
.B(n_38),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3252),
.B(n_38),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3111),
.A2(n_962),
.B(n_961),
.Y(n_3369)
);

NOR2xp67_ASAP7_75t_L g3370 ( 
.A(n_3243),
.B(n_964),
.Y(n_3370)
);

OAI21x1_ASAP7_75t_L g3371 ( 
.A1(n_3186),
.A2(n_968),
.B(n_967),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3171),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_3372)
);

OAI21x1_ASAP7_75t_L g3373 ( 
.A1(n_3141),
.A2(n_974),
.B(n_972),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3179),
.B(n_39),
.Y(n_3374)
);

OAI21x1_ASAP7_75t_L g3375 ( 
.A1(n_3120),
.A2(n_976),
.B(n_975),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_3184),
.B(n_40),
.Y(n_3376)
);

AOI21x1_ASAP7_75t_SL g3377 ( 
.A1(n_3235),
.A2(n_41),
.B(n_42),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3193),
.B(n_3196),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3197),
.B(n_42),
.Y(n_3379)
);

OAI21x1_ASAP7_75t_L g3380 ( 
.A1(n_3119),
.A2(n_981),
.B(n_980),
.Y(n_3380)
);

A2O1A1Ixp33_ASAP7_75t_L g3381 ( 
.A1(n_3300),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_3381)
);

OAI21x1_ASAP7_75t_L g3382 ( 
.A1(n_3146),
.A2(n_986),
.B(n_982),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3198),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3207),
.B(n_3232),
.Y(n_3384)
);

NOR3xp33_ASAP7_75t_SL g3385 ( 
.A(n_3272),
.B(n_3269),
.C(n_3181),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3236),
.Y(n_3386)
);

AOI21x1_ASAP7_75t_L g3387 ( 
.A1(n_3148),
.A2(n_988),
.B(n_987),
.Y(n_3387)
);

AO31x2_ASAP7_75t_L g3388 ( 
.A1(n_3202),
.A2(n_990),
.A3(n_993),
.B(n_989),
.Y(n_3388)
);

OAI21x1_ASAP7_75t_L g3389 ( 
.A1(n_3153),
.A2(n_995),
.B(n_994),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3242),
.B(n_44),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3227),
.Y(n_3391)
);

INVx2_ASAP7_75t_SL g3392 ( 
.A(n_3122),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_3209),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_3157),
.A2(n_997),
.B(n_996),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3262),
.B(n_45),
.Y(n_3395)
);

AOI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_3231),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_3396)
);

AO31x2_ASAP7_75t_L g3397 ( 
.A1(n_3270),
.A2(n_999),
.A3(n_1001),
.B(n_998),
.Y(n_3397)
);

OAI21x1_ASAP7_75t_SL g3398 ( 
.A1(n_3191),
.A2(n_1003),
.B(n_1002),
.Y(n_3398)
);

A2O1A1Ixp33_ASAP7_75t_L g3399 ( 
.A1(n_3273),
.A2(n_3180),
.B(n_3155),
.C(n_3225),
.Y(n_3399)
);

NAND2x1p5_ASAP7_75t_L g3400 ( 
.A(n_3227),
.B(n_1008),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3267),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3174),
.A2(n_1006),
.B(n_1004),
.Y(n_3402)
);

A2O1A1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_3118),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_3403)
);

NAND3xp33_ASAP7_75t_L g3404 ( 
.A(n_3109),
.B(n_50),
.C(n_51),
.Y(n_3404)
);

OAI21x1_ASAP7_75t_L g3405 ( 
.A1(n_3259),
.A2(n_1012),
.B(n_1009),
.Y(n_3405)
);

AOI21x1_ASAP7_75t_L g3406 ( 
.A1(n_3213),
.A2(n_1016),
.B(n_1014),
.Y(n_3406)
);

NOR3xp33_ASAP7_75t_L g3407 ( 
.A(n_3168),
.B(n_50),
.C(n_52),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3268),
.B(n_52),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3271),
.B(n_53),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3249),
.B(n_54),
.Y(n_3410)
);

OAI21x1_ASAP7_75t_L g3411 ( 
.A1(n_3261),
.A2(n_1018),
.B(n_1017),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3221),
.A2(n_3150),
.B(n_3295),
.Y(n_3412)
);

NAND2x1p5_ASAP7_75t_L g3413 ( 
.A(n_3122),
.B(n_1021),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3113),
.B(n_54),
.Y(n_3414)
);

NOR4xp25_ASAP7_75t_L g3415 ( 
.A(n_3228),
.B(n_57),
.C(n_55),
.D(n_56),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3281),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3176),
.B(n_3284),
.Y(n_3417)
);

INVx3_ASAP7_75t_L g3418 ( 
.A(n_3167),
.Y(n_3418)
);

OAI21x1_ASAP7_75t_L g3419 ( 
.A1(n_3265),
.A2(n_1023),
.B(n_1019),
.Y(n_3419)
);

O2A1O1Ixp5_ASAP7_75t_SL g3420 ( 
.A1(n_3195),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3289),
.B(n_58),
.Y(n_3421)
);

AO31x2_ASAP7_75t_L g3422 ( 
.A1(n_3234),
.A2(n_1025),
.A3(n_1030),
.B(n_1024),
.Y(n_3422)
);

CKINVDCx20_ASAP7_75t_R g3423 ( 
.A(n_3238),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3115),
.Y(n_3424)
);

INVx2_ASAP7_75t_SL g3425 ( 
.A(n_3127),
.Y(n_3425)
);

AO31x2_ASAP7_75t_L g3426 ( 
.A1(n_3178),
.A2(n_1034),
.A3(n_1035),
.B(n_1031),
.Y(n_3426)
);

AOI221x1_ASAP7_75t_L g3427 ( 
.A1(n_3130),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_62),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_3211),
.A2(n_1039),
.B(n_1038),
.Y(n_3428)
);

OAI21x1_ASAP7_75t_L g3429 ( 
.A1(n_3276),
.A2(n_1042),
.B(n_1041),
.Y(n_3429)
);

CKINVDCx5p33_ASAP7_75t_R g3430 ( 
.A(n_3241),
.Y(n_3430)
);

AOI211x1_ASAP7_75t_L g3431 ( 
.A1(n_3192),
.A2(n_64),
.B(n_61),
.C(n_63),
.Y(n_3431)
);

BUFx4f_ASAP7_75t_L g3432 ( 
.A(n_3127),
.Y(n_3432)
);

INVxp67_ASAP7_75t_SL g3433 ( 
.A(n_3136),
.Y(n_3433)
);

BUFx2_ASAP7_75t_L g3434 ( 
.A(n_3301),
.Y(n_3434)
);

OAI21x1_ASAP7_75t_L g3435 ( 
.A1(n_3280),
.A2(n_1046),
.B(n_1044),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3205),
.B(n_63),
.Y(n_3436)
);

A2O1A1Ixp33_ASAP7_75t_L g3437 ( 
.A1(n_3240),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_3437)
);

O2A1O1Ixp5_ASAP7_75t_L g3438 ( 
.A1(n_3266),
.A2(n_69),
.B(n_66),
.C(n_68),
.Y(n_3438)
);

OAI21x1_ASAP7_75t_L g3439 ( 
.A1(n_3283),
.A2(n_1048),
.B(n_1047),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_3220),
.A2(n_1050),
.B(n_1049),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3121),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_SL g3442 ( 
.A(n_3307),
.B(n_1053),
.Y(n_3442)
);

OAI21x1_ASAP7_75t_L g3443 ( 
.A1(n_3291),
.A2(n_1055),
.B(n_1052),
.Y(n_3443)
);

OAI21x1_ASAP7_75t_L g3444 ( 
.A1(n_3123),
.A2(n_1057),
.B(n_1056),
.Y(n_3444)
);

O2A1O1Ixp5_ASAP7_75t_SL g3445 ( 
.A1(n_3285),
.A2(n_71),
.B(n_68),
.C(n_70),
.Y(n_3445)
);

BUFx2_ASAP7_75t_L g3446 ( 
.A(n_3194),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3158),
.Y(n_3447)
);

CKINVDCx20_ASAP7_75t_R g3448 ( 
.A(n_3172),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_3305),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_3449)
);

BUFx3_ASAP7_75t_L g3450 ( 
.A(n_3167),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3304),
.B(n_72),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3217),
.B(n_3182),
.Y(n_3452)
);

INVx3_ASAP7_75t_L g3453 ( 
.A(n_3256),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3215),
.A2(n_1060),
.B(n_1059),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3175),
.B(n_73),
.Y(n_3455)
);

OAI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3183),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_3456)
);

OR2x6_ASAP7_75t_L g3457 ( 
.A(n_3222),
.B(n_1061),
.Y(n_3457)
);

AO21x2_ASAP7_75t_L g3458 ( 
.A1(n_3212),
.A2(n_1067),
.B(n_1063),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_3151),
.B(n_74),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3189),
.Y(n_3460)
);

OAI21x1_ASAP7_75t_L g3461 ( 
.A1(n_3199),
.A2(n_1073),
.B(n_1070),
.Y(n_3461)
);

OAI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_3224),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3275),
.B(n_77),
.Y(n_3463)
);

AOI21xp33_ASAP7_75t_L g3464 ( 
.A1(n_3112),
.A2(n_78),
.B(n_80),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3277),
.A2(n_1076),
.B(n_1074),
.Y(n_3465)
);

AOI21x1_ASAP7_75t_SL g3466 ( 
.A1(n_3138),
.A2(n_80),
.B(n_82),
.Y(n_3466)
);

OAI21x1_ASAP7_75t_L g3467 ( 
.A1(n_3219),
.A2(n_1079),
.B(n_1077),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3229),
.B(n_82),
.Y(n_3468)
);

OAI21x1_ASAP7_75t_L g3469 ( 
.A1(n_3206),
.A2(n_1089),
.B(n_1085),
.Y(n_3469)
);

OAI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3132),
.A2(n_1094),
.B(n_1093),
.Y(n_3470)
);

OAI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3116),
.A2(n_1097),
.B(n_1095),
.Y(n_3471)
);

OA21x2_ASAP7_75t_L g3472 ( 
.A1(n_3214),
.A2(n_1099),
.B(n_1098),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3143),
.B(n_83),
.Y(n_3473)
);

AND2x4_ASAP7_75t_L g3474 ( 
.A(n_3256),
.B(n_1101),
.Y(n_3474)
);

A2O1A1Ixp33_ASAP7_75t_L g3475 ( 
.A1(n_3255),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_3475)
);

AO31x2_ASAP7_75t_L g3476 ( 
.A1(n_3187),
.A2(n_1103),
.A3(n_1106),
.B(n_1102),
.Y(n_3476)
);

HB1xp67_ASAP7_75t_L g3477 ( 
.A(n_3230),
.Y(n_3477)
);

AOI21x1_ASAP7_75t_L g3478 ( 
.A1(n_3218),
.A2(n_1109),
.B(n_1107),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3244),
.A2(n_1111),
.B(n_1110),
.Y(n_3479)
);

AOI21x1_ASAP7_75t_L g3480 ( 
.A1(n_3126),
.A2(n_3297),
.B(n_3223),
.Y(n_3480)
);

AO31x2_ASAP7_75t_L g3481 ( 
.A1(n_3274),
.A2(n_3287),
.A3(n_3159),
.B(n_3296),
.Y(n_3481)
);

NOR2x1_ASAP7_75t_SL g3482 ( 
.A(n_3245),
.B(n_1112),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3147),
.B(n_85),
.Y(n_3483)
);

AO31x2_ASAP7_75t_L g3484 ( 
.A1(n_3245),
.A2(n_1114),
.A3(n_1117),
.B(n_1113),
.Y(n_3484)
);

INVx8_ASAP7_75t_L g3485 ( 
.A(n_3230),
.Y(n_3485)
);

INVxp67_ASAP7_75t_L g3486 ( 
.A(n_3188),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3278),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3278),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3223),
.Y(n_3489)
);

OAI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3288),
.A2(n_1120),
.B(n_1119),
.Y(n_3490)
);

NOR2xp33_ASAP7_75t_L g3491 ( 
.A(n_3156),
.B(n_86),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_3210),
.B(n_86),
.Y(n_3492)
);

AO22x2_ASAP7_75t_L g3493 ( 
.A1(n_3272),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_3493)
);

AO22x2_ASAP7_75t_L g3494 ( 
.A1(n_3272),
.A2(n_91),
.B1(n_87),
.B2(n_90),
.Y(n_3494)
);

OAI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_3226),
.A2(n_1123),
.B(n_1122),
.Y(n_3495)
);

OAI21x1_ASAP7_75t_L g3496 ( 
.A1(n_3201),
.A2(n_1126),
.B(n_1124),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3246),
.A2(n_1129),
.B(n_1127),
.Y(n_3497)
);

OAI21x1_ASAP7_75t_L g3498 ( 
.A1(n_3201),
.A2(n_1131),
.B(n_1130),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3129),
.B(n_91),
.Y(n_3499)
);

AOI21x1_ASAP7_75t_L g3500 ( 
.A1(n_3247),
.A2(n_1134),
.B(n_1133),
.Y(n_3500)
);

OAI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3226),
.A2(n_1137),
.B(n_1135),
.Y(n_3501)
);

OAI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3226),
.A2(n_1139),
.B(n_1138),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3108),
.B(n_93),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3347),
.B(n_93),
.Y(n_3504)
);

OAI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3491),
.A2(n_94),
.B(n_95),
.Y(n_3505)
);

INVxp67_ASAP7_75t_L g3506 ( 
.A(n_3446),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3464),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3322),
.A2(n_96),
.B(n_97),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3452),
.B(n_98),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_3453),
.B(n_1140),
.Y(n_3510)
);

OAI21x1_ASAP7_75t_L g3511 ( 
.A1(n_3329),
.A2(n_1146),
.B(n_1142),
.Y(n_3511)
);

BUFx3_ASAP7_75t_L g3512 ( 
.A(n_3432),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3434),
.Y(n_3513)
);

OAI21x1_ASAP7_75t_L g3514 ( 
.A1(n_3335),
.A2(n_1148),
.B(n_1147),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3378),
.Y(n_3515)
);

HB1xp67_ASAP7_75t_L g3516 ( 
.A(n_3363),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3311),
.B(n_99),
.Y(n_3517)
);

OAI21x1_ASAP7_75t_L g3518 ( 
.A1(n_3412),
.A2(n_1150),
.B(n_1149),
.Y(n_3518)
);

AND2x2_ASAP7_75t_SL g3519 ( 
.A(n_3415),
.B(n_99),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3384),
.Y(n_3520)
);

INVxp67_ASAP7_75t_SL g3521 ( 
.A(n_3433),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3450),
.Y(n_3522)
);

OAI21x1_ASAP7_75t_L g3523 ( 
.A1(n_3496),
.A2(n_1154),
.B(n_1153),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3332),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_SL g3525 ( 
.A1(n_3367),
.A2(n_3333),
.B1(n_3404),
.B2(n_3490),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3348),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3354),
.Y(n_3527)
);

OAI21x1_ASAP7_75t_L g3528 ( 
.A1(n_3498),
.A2(n_1157),
.B(n_1155),
.Y(n_3528)
);

OAI21x1_ASAP7_75t_L g3529 ( 
.A1(n_3371),
.A2(n_1159),
.B(n_1158),
.Y(n_3529)
);

AND2x4_ASAP7_75t_L g3530 ( 
.A(n_3418),
.B(n_1160),
.Y(n_3530)
);

AOI221xp5_ASAP7_75t_L g3531 ( 
.A1(n_3323),
.A2(n_3407),
.B1(n_3310),
.B2(n_3475),
.C(n_3483),
.Y(n_3531)
);

HB1xp67_ASAP7_75t_L g3532 ( 
.A(n_3392),
.Y(n_3532)
);

OAI21x1_ASAP7_75t_L g3533 ( 
.A1(n_3405),
.A2(n_1163),
.B(n_1161),
.Y(n_3533)
);

OAI21x1_ASAP7_75t_L g3534 ( 
.A1(n_3411),
.A2(n_1165),
.B(n_1164),
.Y(n_3534)
);

OA21x2_ASAP7_75t_L g3535 ( 
.A1(n_3495),
.A2(n_1168),
.B(n_1167),
.Y(n_3535)
);

AOI22xp33_ASAP7_75t_L g3536 ( 
.A1(n_3320),
.A2(n_3346),
.B1(n_3338),
.B2(n_3342),
.Y(n_3536)
);

OA21x2_ASAP7_75t_L g3537 ( 
.A1(n_3501),
.A2(n_1170),
.B(n_1169),
.Y(n_3537)
);

AND2x4_ASAP7_75t_SL g3538 ( 
.A(n_3312),
.B(n_1172),
.Y(n_3538)
);

CKINVDCx5p33_ASAP7_75t_R g3539 ( 
.A(n_3330),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3308),
.A2(n_1346),
.B(n_1342),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3503),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_3541)
);

NAND3xp33_ASAP7_75t_L g3542 ( 
.A(n_3385),
.B(n_100),
.C(n_101),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_SL g3543 ( 
.A1(n_3309),
.A2(n_103),
.B(n_104),
.Y(n_3543)
);

HB1xp67_ASAP7_75t_L g3544 ( 
.A(n_3425),
.Y(n_3544)
);

OAI221xp5_ASAP7_75t_L g3545 ( 
.A1(n_3317),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.C(n_108),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3417),
.A2(n_3364),
.B1(n_3399),
.B2(n_3315),
.Y(n_3546)
);

OAI21x1_ASAP7_75t_L g3547 ( 
.A1(n_3373),
.A2(n_1175),
.B(n_1174),
.Y(n_3547)
);

AO21x2_ASAP7_75t_L g3548 ( 
.A1(n_3502),
.A2(n_1179),
.B(n_1177),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3357),
.Y(n_3549)
);

OAI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3344),
.A2(n_3319),
.B(n_3324),
.Y(n_3550)
);

O2A1O1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_3403),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_3551)
);

OAI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3331),
.A2(n_3352),
.B(n_3349),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3360),
.A2(n_3353),
.B1(n_3355),
.B2(n_3350),
.Y(n_3553)
);

OAI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3375),
.A2(n_1181),
.B(n_1180),
.Y(n_3554)
);

O2A1O1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_3381),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_3555)
);

OAI22xp5_ASAP7_75t_L g3556 ( 
.A1(n_3436),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3556)
);

AO21x2_ASAP7_75t_L g3557 ( 
.A1(n_3351),
.A2(n_1185),
.B(n_1184),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3423),
.B(n_1186),
.Y(n_3558)
);

BUFx3_ASAP7_75t_L g3559 ( 
.A(n_3485),
.Y(n_3559)
);

OAI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3366),
.A2(n_112),
.B(n_114),
.Y(n_3560)
);

AO32x2_ASAP7_75t_L g3561 ( 
.A1(n_3372),
.A2(n_116),
.A3(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_3561)
);

BUFx2_ASAP7_75t_R g3562 ( 
.A(n_3340),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3383),
.Y(n_3563)
);

AOI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3499),
.A2(n_3494),
.B1(n_3493),
.B2(n_3470),
.Y(n_3564)
);

OAI21x1_ASAP7_75t_L g3565 ( 
.A1(n_3380),
.A2(n_1189),
.B(n_1188),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_L g3566 ( 
.A1(n_3471),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3316),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_3489),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3568)
);

AOI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3492),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_3424),
.B(n_121),
.Y(n_3570)
);

OAI22xp33_ASAP7_75t_L g3571 ( 
.A1(n_3396),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3451),
.B(n_122),
.Y(n_3572)
);

BUFx3_ASAP7_75t_L g3573 ( 
.A(n_3485),
.Y(n_3573)
);

INVx1_ASAP7_75t_SL g3574 ( 
.A(n_3391),
.Y(n_3574)
);

BUFx6f_ASAP7_75t_SL g3575 ( 
.A(n_3328),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3337),
.Y(n_3576)
);

OAI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3321),
.A2(n_125),
.B(n_126),
.Y(n_3577)
);

AND2x4_ASAP7_75t_L g3578 ( 
.A(n_3477),
.B(n_1190),
.Y(n_3578)
);

A2O1A1Ixp33_ASAP7_75t_L g3579 ( 
.A1(n_3356),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_3579)
);

BUFx6f_ASAP7_75t_L g3580 ( 
.A(n_3326),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_3326),
.Y(n_3581)
);

BUFx2_ASAP7_75t_R g3582 ( 
.A(n_3345),
.Y(n_3582)
);

INVx3_ASAP7_75t_L g3583 ( 
.A(n_3334),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3368),
.B(n_3473),
.Y(n_3584)
);

OAI21x1_ASAP7_75t_L g3585 ( 
.A1(n_3382),
.A2(n_1192),
.B(n_1191),
.Y(n_3585)
);

OAI21x1_ASAP7_75t_L g3586 ( 
.A1(n_3389),
.A2(n_1194),
.B(n_1193),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_3361),
.A2(n_3456),
.B1(n_3462),
.B2(n_3459),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3386),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_3393),
.B(n_1195),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3401),
.Y(n_3590)
);

OAI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3394),
.A2(n_1198),
.B(n_1197),
.Y(n_3591)
);

NOR2x1_ASAP7_75t_SL g3592 ( 
.A(n_3313),
.B(n_1199),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3361),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_3593)
);

HB1xp67_ASAP7_75t_L g3594 ( 
.A(n_3327),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_3487),
.B(n_1203),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3410),
.B(n_1204),
.Y(n_3596)
);

OR2x2_ASAP7_75t_L g3597 ( 
.A(n_3441),
.B(n_129),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3447),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3460),
.Y(n_3599)
);

AO31x2_ASAP7_75t_L g3600 ( 
.A1(n_3454),
.A2(n_1206),
.A3(n_1208),
.B(n_1205),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3358),
.A2(n_1356),
.B(n_1355),
.Y(n_3601)
);

NAND2xp33_ASAP7_75t_L g3602 ( 
.A(n_3361),
.B(n_131),
.Y(n_3602)
);

OAI21x1_ASAP7_75t_L g3603 ( 
.A1(n_3419),
.A2(n_1210),
.B(n_1209),
.Y(n_3603)
);

OR2x6_ASAP7_75t_L g3604 ( 
.A(n_3457),
.B(n_1211),
.Y(n_3604)
);

AO21x1_ASAP7_75t_L g3605 ( 
.A1(n_3369),
.A2(n_130),
.B(n_131),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3455),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3429),
.A2(n_1214),
.B(n_1213),
.Y(n_3607)
);

OR2x6_ASAP7_75t_SL g3608 ( 
.A(n_3430),
.B(n_130),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3435),
.A2(n_1216),
.B(n_1215),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3439),
.A2(n_1218),
.B(n_1217),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3463),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3325),
.B(n_132),
.Y(n_3612)
);

OA21x2_ASAP7_75t_L g3613 ( 
.A1(n_3438),
.A2(n_1223),
.B(n_1219),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3365),
.Y(n_3614)
);

OA21x2_ASAP7_75t_L g3615 ( 
.A1(n_3444),
.A2(n_1226),
.B(n_1225),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3374),
.Y(n_3616)
);

CKINVDCx5p33_ASAP7_75t_R g3617 ( 
.A(n_3448),
.Y(n_3617)
);

AOI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3486),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3443),
.A2(n_1232),
.B(n_1229),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3421),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3461),
.A2(n_1236),
.B(n_1233),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3481),
.B(n_135),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3481),
.B(n_136),
.Y(n_3623)
);

AND2x4_ASAP7_75t_L g3624 ( 
.A(n_3488),
.B(n_1238),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3325),
.B(n_137),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3465),
.A2(n_1240),
.B(n_1239),
.Y(n_3626)
);

OAI21x1_ASAP7_75t_L g3627 ( 
.A1(n_3387),
.A2(n_1243),
.B(n_1242),
.Y(n_3627)
);

BUFx6f_ASAP7_75t_L g3628 ( 
.A(n_3328),
.Y(n_3628)
);

CKINVDCx5p33_ASAP7_75t_R g3629 ( 
.A(n_3376),
.Y(n_3629)
);

CKINVDCx5p33_ASAP7_75t_R g3630 ( 
.A(n_3414),
.Y(n_3630)
);

OA21x2_ASAP7_75t_L g3631 ( 
.A1(n_3469),
.A2(n_1246),
.B(n_1244),
.Y(n_3631)
);

INVxp67_ASAP7_75t_SL g3632 ( 
.A(n_3379),
.Y(n_3632)
);

HB1xp67_ASAP7_75t_L g3633 ( 
.A(n_3313),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3416),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3634)
);

BUFx3_ASAP7_75t_L g3635 ( 
.A(n_3359),
.Y(n_3635)
);

O2A1O1Ixp33_ASAP7_75t_SL g3636 ( 
.A1(n_3437),
.A2(n_143),
.B(n_139),
.C(n_141),
.Y(n_3636)
);

BUFx3_ASAP7_75t_L g3637 ( 
.A(n_3474),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3390),
.Y(n_3638)
);

AND2x4_ASAP7_75t_L g3639 ( 
.A(n_3480),
.B(n_1247),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3395),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3406),
.A2(n_1251),
.B(n_1250),
.Y(n_3641)
);

BUFx4_ASAP7_75t_SL g3642 ( 
.A(n_3457),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3408),
.B(n_144),
.Y(n_3643)
);

CKINVDCx16_ASAP7_75t_R g3644 ( 
.A(n_3442),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3409),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3468),
.Y(n_3646)
);

AO31x2_ASAP7_75t_L g3647 ( 
.A1(n_3427),
.A2(n_1253),
.A3(n_1254),
.B(n_1252),
.Y(n_3647)
);

AO21x2_ASAP7_75t_L g3648 ( 
.A1(n_3362),
.A2(n_3318),
.B(n_3458),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_3336),
.Y(n_3649)
);

INVx3_ASAP7_75t_L g3650 ( 
.A(n_3400),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3500),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3339),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3632),
.B(n_3431),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3516),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_SL g3655 ( 
.A1(n_3560),
.A2(n_3479),
.B(n_3472),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3645),
.B(n_3449),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3584),
.B(n_3484),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3614),
.B(n_3482),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3616),
.B(n_3445),
.Y(n_3659)
);

OA21x2_ASAP7_75t_L g3660 ( 
.A1(n_3550),
.A2(n_3402),
.B(n_3440),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3622),
.B(n_3484),
.Y(n_3661)
);

OA21x2_ASAP7_75t_L g3662 ( 
.A1(n_3577),
.A2(n_3497),
.B(n_3478),
.Y(n_3662)
);

INVxp67_ASAP7_75t_SL g3663 ( 
.A(n_3521),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3635),
.B(n_3370),
.Y(n_3664)
);

OAI22xp5_ASAP7_75t_L g3665 ( 
.A1(n_3525),
.A2(n_3413),
.B1(n_3428),
.B2(n_3343),
.Y(n_3665)
);

AND2x4_ASAP7_75t_L g3666 ( 
.A(n_3583),
.B(n_3467),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3526),
.Y(n_3667)
);

INVx1_ASAP7_75t_SL g3668 ( 
.A(n_3513),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3567),
.Y(n_3669)
);

AOI211xp5_ASAP7_75t_L g3670 ( 
.A1(n_3505),
.A2(n_3341),
.B(n_3466),
.C(n_3377),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_3512),
.Y(n_3671)
);

BUFx3_ASAP7_75t_L g3672 ( 
.A(n_3559),
.Y(n_3672)
);

AND2x2_ASAP7_75t_SL g3673 ( 
.A(n_3602),
.B(n_3420),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3637),
.B(n_3388),
.Y(n_3674)
);

O2A1O1Ixp5_ASAP7_75t_L g3675 ( 
.A1(n_3605),
.A2(n_3397),
.B(n_3388),
.C(n_3422),
.Y(n_3675)
);

AOI21xp5_ASAP7_75t_SL g3676 ( 
.A1(n_3604),
.A2(n_3398),
.B(n_3314),
.Y(n_3676)
);

O2A1O1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3517),
.A2(n_3397),
.B(n_3422),
.C(n_3476),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3506),
.B(n_3314),
.Y(n_3678)
);

OA21x2_ASAP7_75t_L g3679 ( 
.A1(n_3552),
.A2(n_3476),
.B(n_3426),
.Y(n_3679)
);

A2O1A1Ixp33_ASAP7_75t_L g3680 ( 
.A1(n_3531),
.A2(n_3426),
.B(n_147),
.C(n_145),
.Y(n_3680)
);

A2O1A1Ixp33_ASAP7_75t_L g3681 ( 
.A1(n_3551),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3564),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.Y(n_3682)
);

AOI21x1_ASAP7_75t_SL g3683 ( 
.A1(n_3612),
.A2(n_3625),
.B(n_3623),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3576),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3572),
.B(n_1256),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3504),
.B(n_1258),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3638),
.B(n_3640),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3644),
.A2(n_151),
.B1(n_148),
.B2(n_149),
.Y(n_3688)
);

AOI21x1_ASAP7_75t_SL g3689 ( 
.A1(n_3639),
.A2(n_151),
.B(n_152),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3646),
.B(n_1259),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3508),
.B(n_1260),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3588),
.Y(n_3692)
);

AND2x4_ASAP7_75t_L g3693 ( 
.A(n_3522),
.B(n_1261),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3590),
.Y(n_3694)
);

INVxp67_ASAP7_75t_L g3695 ( 
.A(n_3532),
.Y(n_3695)
);

AOI21x1_ASAP7_75t_SL g3696 ( 
.A1(n_3509),
.A2(n_153),
.B(n_155),
.Y(n_3696)
);

OR2x2_ASAP7_75t_L g3697 ( 
.A(n_3515),
.B(n_155),
.Y(n_3697)
);

AOI21x1_ASAP7_75t_SL g3698 ( 
.A1(n_3643),
.A2(n_156),
.B(n_157),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3520),
.B(n_156),
.Y(n_3699)
);

O2A1O1Ixp33_ASAP7_75t_L g3700 ( 
.A1(n_3545),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3598),
.Y(n_3701)
);

OR2x2_ASAP7_75t_L g3702 ( 
.A(n_3524),
.B(n_158),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3527),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3549),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3606),
.B(n_1263),
.Y(n_3705)
);

INVx1_ASAP7_75t_SL g3706 ( 
.A(n_3574),
.Y(n_3706)
);

AOI21x1_ASAP7_75t_SL g3707 ( 
.A1(n_3595),
.A2(n_159),
.B(n_160),
.Y(n_3707)
);

BUFx4f_ASAP7_75t_SL g3708 ( 
.A(n_3580),
.Y(n_3708)
);

AOI21xp5_ASAP7_75t_SL g3709 ( 
.A1(n_3604),
.A2(n_1277),
.B(n_1267),
.Y(n_3709)
);

HB1xp67_ASAP7_75t_L g3710 ( 
.A(n_3563),
.Y(n_3710)
);

OA21x2_ASAP7_75t_L g3711 ( 
.A1(n_3514),
.A2(n_160),
.B(n_161),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3546),
.A2(n_1266),
.B(n_1264),
.Y(n_3712)
);

NOR2xp67_ASAP7_75t_L g3713 ( 
.A(n_3594),
.B(n_3611),
.Y(n_3713)
);

AOI21x1_ASAP7_75t_SL g3714 ( 
.A1(n_3624),
.A2(n_161),
.B(n_162),
.Y(n_3714)
);

INVx2_ASAP7_75t_SL g3715 ( 
.A(n_3573),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3536),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3599),
.Y(n_3717)
);

O2A1O1Ixp33_ASAP7_75t_L g3718 ( 
.A1(n_3579),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3570),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3553),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_3720)
);

OAI22xp5_ASAP7_75t_L g3721 ( 
.A1(n_3587),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_3721)
);

OAI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3630),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3558),
.B(n_1268),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3597),
.B(n_172),
.Y(n_3724)
);

OAI22xp5_ASAP7_75t_L g3725 ( 
.A1(n_3629),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_3725)
);

OAI22x1_ASAP7_75t_L g3726 ( 
.A1(n_3542),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3543),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3519),
.B(n_1269),
.Y(n_3728)
);

AOI21x1_ASAP7_75t_SL g3729 ( 
.A1(n_3633),
.A2(n_3578),
.B(n_3510),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3651),
.Y(n_3730)
);

AOI21xp5_ASAP7_75t_SL g3731 ( 
.A1(n_3555),
.A2(n_1282),
.B(n_1271),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3566),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3596),
.B(n_1270),
.Y(n_3733)
);

CKINVDCx5p33_ASAP7_75t_R g3734 ( 
.A(n_3617),
.Y(n_3734)
);

AOI221x1_ASAP7_75t_SL g3735 ( 
.A1(n_3556),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.C(n_181),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3593),
.B(n_1273),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_3544),
.Y(n_3737)
);

OAI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_3569),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3652),
.Y(n_3739)
);

AOI21x1_ASAP7_75t_SL g3740 ( 
.A1(n_3530),
.A2(n_182),
.B(n_183),
.Y(n_3740)
);

AOI211xp5_ASAP7_75t_L g3741 ( 
.A1(n_3571),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_3741)
);

HB1xp67_ASAP7_75t_L g3742 ( 
.A(n_3628),
.Y(n_3742)
);

CKINVDCx16_ASAP7_75t_R g3743 ( 
.A(n_3580),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3538),
.B(n_1274),
.Y(n_3744)
);

NOR2xp67_ASAP7_75t_L g3745 ( 
.A(n_3539),
.B(n_1339),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3647),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3581),
.Y(n_3747)
);

AND2x4_ASAP7_75t_L g3748 ( 
.A(n_3668),
.B(n_3628),
.Y(n_3748)
);

AO21x2_ASAP7_75t_L g3749 ( 
.A1(n_3746),
.A2(n_3648),
.B(n_3511),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3657),
.B(n_3649),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3717),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3669),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3654),
.B(n_3541),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3661),
.B(n_3649),
.Y(n_3754)
);

BUFx3_ASAP7_75t_L g3755 ( 
.A(n_3671),
.Y(n_3755)
);

OA21x2_ASAP7_75t_L g3756 ( 
.A1(n_3659),
.A2(n_3641),
.B(n_3627),
.Y(n_3756)
);

INVx3_ASAP7_75t_L g3757 ( 
.A(n_3672),
.Y(n_3757)
);

AO21x2_ASAP7_75t_L g3758 ( 
.A1(n_3676),
.A2(n_3540),
.B(n_3548),
.Y(n_3758)
);

BUFx3_ASAP7_75t_L g3759 ( 
.A(n_3747),
.Y(n_3759)
);

INVx3_ASAP7_75t_L g3760 ( 
.A(n_3708),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3684),
.Y(n_3761)
);

INVxp33_ASAP7_75t_L g3762 ( 
.A(n_3742),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3743),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3680),
.A2(n_3518),
.B(n_3601),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3704),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3719),
.Y(n_3766)
);

AND2x4_ASAP7_75t_L g3767 ( 
.A(n_3674),
.B(n_3650),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3703),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3710),
.Y(n_3769)
);

AO21x2_ASAP7_75t_L g3770 ( 
.A1(n_3677),
.A2(n_3626),
.B(n_3621),
.Y(n_3770)
);

INVx2_ASAP7_75t_SL g3771 ( 
.A(n_3715),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3663),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3692),
.B(n_3647),
.Y(n_3773)
);

NOR3xp33_ASAP7_75t_L g3774 ( 
.A(n_3700),
.B(n_3636),
.C(n_3618),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3694),
.Y(n_3775)
);

BUFx3_ASAP7_75t_L g3776 ( 
.A(n_3734),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3706),
.B(n_3589),
.Y(n_3777)
);

BUFx12f_ASAP7_75t_L g3778 ( 
.A(n_3724),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3701),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3678),
.B(n_3608),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3730),
.Y(n_3781)
);

AO21x2_ASAP7_75t_L g3782 ( 
.A1(n_3655),
.A2(n_3529),
.B(n_3565),
.Y(n_3782)
);

INVxp67_ASAP7_75t_L g3783 ( 
.A(n_3737),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3664),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3739),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3667),
.Y(n_3786)
);

INVx8_ASAP7_75t_L g3787 ( 
.A(n_3693),
.Y(n_3787)
);

AO21x2_ASAP7_75t_L g3788 ( 
.A1(n_3665),
.A2(n_3586),
.B(n_3585),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3713),
.B(n_3685),
.Y(n_3789)
);

OA21x2_ASAP7_75t_L g3790 ( 
.A1(n_3675),
.A2(n_3591),
.B(n_3534),
.Y(n_3790)
);

OA21x2_ASAP7_75t_L g3791 ( 
.A1(n_3653),
.A2(n_3533),
.B(n_3607),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3681),
.A2(n_3507),
.B(n_3620),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3687),
.Y(n_3793)
);

HB1xp67_ASAP7_75t_L g3794 ( 
.A(n_3695),
.Y(n_3794)
);

BUFx8_ASAP7_75t_SL g3795 ( 
.A(n_3723),
.Y(n_3795)
);

OA21x2_ASAP7_75t_L g3796 ( 
.A1(n_3658),
.A2(n_3619),
.B(n_3554),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3679),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3744),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3679),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3699),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3702),
.B(n_3600),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3727),
.Y(n_3802)
);

BUFx2_ASAP7_75t_L g3803 ( 
.A(n_3666),
.Y(n_3803)
);

AO21x2_ASAP7_75t_L g3804 ( 
.A1(n_3731),
.A2(n_3603),
.B(n_3547),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3686),
.B(n_3728),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3697),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3711),
.Y(n_3807)
);

HB1xp67_ASAP7_75t_L g3808 ( 
.A(n_3656),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3711),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3690),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3673),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3691),
.B(n_3592),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3726),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3705),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3660),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3733),
.B(n_3535),
.Y(n_3816)
);

AND2x4_ASAP7_75t_L g3817 ( 
.A(n_3745),
.B(n_3581),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3662),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3660),
.Y(n_3819)
);

AND2x4_ASAP7_75t_L g3820 ( 
.A(n_3736),
.B(n_3600),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3732),
.A2(n_3634),
.B1(n_3568),
.B2(n_3575),
.Y(n_3821)
);

OR2x6_ASAP7_75t_L g3822 ( 
.A(n_3709),
.B(n_3642),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3662),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3720),
.Y(n_3824)
);

BUFx6f_ASAP7_75t_L g3825 ( 
.A(n_3729),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3718),
.Y(n_3826)
);

BUFx2_ASAP7_75t_L g3827 ( 
.A(n_3682),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3670),
.B(n_3537),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3716),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3721),
.B(n_3561),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3735),
.Y(n_3831)
);

AOI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_3741),
.A2(n_3738),
.B1(n_3725),
.B2(n_3688),
.Y(n_3832)
);

AO21x2_ASAP7_75t_L g3833 ( 
.A1(n_3712),
.A2(n_3610),
.B(n_3609),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3803),
.B(n_3557),
.Y(n_3834)
);

BUFx3_ASAP7_75t_L g3835 ( 
.A(n_3755),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3750),
.B(n_3562),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3754),
.B(n_3582),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3752),
.Y(n_3838)
);

INVx2_ASAP7_75t_SL g3839 ( 
.A(n_3757),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3751),
.B(n_3613),
.Y(n_3840)
);

BUFx3_ASAP7_75t_L g3841 ( 
.A(n_3759),
.Y(n_3841)
);

OR2x2_ASAP7_75t_L g3842 ( 
.A(n_3765),
.B(n_3631),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3761),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3775),
.Y(n_3844)
);

OAI222xp33_ASAP7_75t_L g3845 ( 
.A1(n_3831),
.A2(n_3722),
.B1(n_3683),
.B2(n_3689),
.C1(n_3561),
.C2(n_3740),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3766),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3769),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3780),
.B(n_3615),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3768),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3793),
.B(n_3523),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3794),
.B(n_3528),
.Y(n_3851)
);

HB1xp67_ASAP7_75t_L g3852 ( 
.A(n_3772),
.Y(n_3852)
);

BUFx2_ASAP7_75t_L g3853 ( 
.A(n_3783),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3762),
.B(n_184),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3781),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3789),
.B(n_185),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3811),
.B(n_186),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3779),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3786),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3785),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3773),
.Y(n_3861)
);

OR2x2_ASAP7_75t_L g3862 ( 
.A(n_3808),
.B(n_187),
.Y(n_3862)
);

BUFx3_ASAP7_75t_L g3863 ( 
.A(n_3760),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3800),
.B(n_187),
.Y(n_3864)
);

BUFx2_ASAP7_75t_L g3865 ( 
.A(n_3802),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3763),
.B(n_188),
.Y(n_3866)
);

OR2x2_ASAP7_75t_L g3867 ( 
.A(n_3801),
.B(n_188),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3807),
.Y(n_3868)
);

HB1xp67_ASAP7_75t_L g3869 ( 
.A(n_3806),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3809),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3805),
.B(n_189),
.Y(n_3871)
);

INVx2_ASAP7_75t_SL g3872 ( 
.A(n_3748),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3797),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3784),
.B(n_189),
.Y(n_3874)
);

AO21x2_ASAP7_75t_L g3875 ( 
.A1(n_3823),
.A2(n_3696),
.B(n_3698),
.Y(n_3875)
);

HB1xp67_ASAP7_75t_L g3876 ( 
.A(n_3813),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3799),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3818),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3815),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3812),
.B(n_190),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3828),
.B(n_191),
.Y(n_3881)
);

INVx1_ASAP7_75t_SL g3882 ( 
.A(n_3771),
.Y(n_3882)
);

HB1xp67_ASAP7_75t_L g3883 ( 
.A(n_3810),
.Y(n_3883)
);

HB1xp67_ASAP7_75t_L g3884 ( 
.A(n_3791),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3819),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3749),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3798),
.B(n_191),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3753),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_L g3889 ( 
.A(n_3777),
.B(n_192),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_3776),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3798),
.B(n_192),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3756),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3767),
.B(n_193),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3778),
.B(n_193),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3796),
.Y(n_3895)
);

BUFx2_ASAP7_75t_L g3896 ( 
.A(n_3814),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3770),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3820),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3816),
.B(n_194),
.Y(n_3899)
);

BUFx3_ASAP7_75t_L g3900 ( 
.A(n_3795),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3788),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3790),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3826),
.B(n_3824),
.Y(n_3903)
);

HB1xp67_ASAP7_75t_L g3904 ( 
.A(n_3825),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3817),
.B(n_195),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3825),
.B(n_196),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3758),
.Y(n_3907)
);

AOI222xp33_ASAP7_75t_L g3908 ( 
.A1(n_3792),
.A2(n_3714),
.B1(n_3707),
.B2(n_222),
.C1(n_204),
.C2(n_230),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3830),
.B(n_3782),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3822),
.B(n_196),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3804),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3829),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3764),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3827),
.B(n_197),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3787),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3833),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3832),
.B(n_197),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3774),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3821),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3752),
.Y(n_3920)
);

BUFx2_ASAP7_75t_L g3921 ( 
.A(n_3803),
.Y(n_3921)
);

AO21x2_ASAP7_75t_L g3922 ( 
.A1(n_3823),
.A2(n_198),
.B(n_199),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3752),
.Y(n_3923)
);

INVxp67_ASAP7_75t_SL g3924 ( 
.A(n_3808),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3751),
.B(n_198),
.Y(n_3925)
);

AND2x4_ASAP7_75t_L g3926 ( 
.A(n_3803),
.B(n_1276),
.Y(n_3926)
);

INVx2_ASAP7_75t_SL g3927 ( 
.A(n_3755),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3752),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3808),
.B(n_199),
.Y(n_3929)
);

INVx3_ASAP7_75t_L g3930 ( 
.A(n_3755),
.Y(n_3930)
);

INVx3_ASAP7_75t_L g3931 ( 
.A(n_3755),
.Y(n_3931)
);

AOI221xp5_ASAP7_75t_L g3932 ( 
.A1(n_3918),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_3932)
);

AOI221xp5_ASAP7_75t_L g3933 ( 
.A1(n_3889),
.A2(n_204),
.B1(n_200),
.B2(n_202),
.C(n_206),
.Y(n_3933)
);

AOI22xp33_ASAP7_75t_L g3934 ( 
.A1(n_3908),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_3934)
);

INVx4_ASAP7_75t_L g3935 ( 
.A(n_3890),
.Y(n_3935)
);

NAND3xp33_ASAP7_75t_L g3936 ( 
.A(n_3913),
.B(n_3907),
.C(n_3888),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3838),
.Y(n_3937)
);

AOI221xp5_ASAP7_75t_L g3938 ( 
.A1(n_3917),
.A2(n_3845),
.B1(n_3876),
.B2(n_3881),
.C(n_3919),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3865),
.Y(n_3939)
);

NAND4xp25_ASAP7_75t_L g3940 ( 
.A(n_3903),
.B(n_212),
.C(n_209),
.D(n_211),
.Y(n_3940)
);

AOI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3848),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3843),
.Y(n_3942)
);

OAI22xp5_ASAP7_75t_SL g3943 ( 
.A1(n_3900),
.A2(n_216),
.B1(n_213),
.B2(n_215),
.Y(n_3943)
);

OAI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3867),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3865),
.Y(n_3945)
);

AOI33xp33_ASAP7_75t_L g3946 ( 
.A1(n_3909),
.A2(n_220),
.A3(n_222),
.B1(n_217),
.B2(n_219),
.B3(n_221),
.Y(n_3946)
);

NOR2xp33_ASAP7_75t_L g3947 ( 
.A(n_3930),
.B(n_219),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3923),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3928),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3920),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3879),
.Y(n_3951)
);

NOR3xp33_ASAP7_75t_L g3952 ( 
.A(n_3929),
.B(n_220),
.C(n_221),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3844),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_SL g3954 ( 
.A(n_3931),
.B(n_223),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3859),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3873),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3877),
.Y(n_3957)
);

NAND3xp33_ASAP7_75t_L g3958 ( 
.A(n_3916),
.B(n_223),
.C(n_224),
.Y(n_3958)
);

OR2x6_ASAP7_75t_L g3959 ( 
.A(n_3927),
.B(n_224),
.Y(n_3959)
);

OAI211xp5_ASAP7_75t_SL g3960 ( 
.A1(n_3864),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3846),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3924),
.B(n_225),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3921),
.B(n_226),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3910),
.A2(n_229),
.B1(n_227),
.B2(n_228),
.Y(n_3964)
);

AND2x4_ASAP7_75t_L g3965 ( 
.A(n_3898),
.B(n_229),
.Y(n_3965)
);

OAI22xp5_ASAP7_75t_L g3966 ( 
.A1(n_3914),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3847),
.Y(n_3967)
);

AO21x2_ASAP7_75t_L g3968 ( 
.A1(n_3886),
.A2(n_231),
.B(n_232),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3852),
.B(n_233),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3901),
.A2(n_1279),
.B(n_1278),
.Y(n_3970)
);

HB1xp67_ASAP7_75t_L g3971 ( 
.A(n_3861),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3869),
.B(n_234),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3883),
.B(n_236),
.Y(n_3973)
);

INVx2_ASAP7_75t_SL g3974 ( 
.A(n_3841),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3885),
.Y(n_3975)
);

AOI221xp5_ASAP7_75t_SL g3976 ( 
.A1(n_3912),
.A2(n_3906),
.B1(n_3899),
.B2(n_3856),
.C(n_3880),
.Y(n_3976)
);

BUFx2_ASAP7_75t_SL g3977 ( 
.A(n_3835),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3896),
.B(n_236),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3853),
.B(n_237),
.Y(n_3979)
);

AOI221xp5_ASAP7_75t_L g3980 ( 
.A1(n_3854),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.C(n_241),
.Y(n_3980)
);

OAI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3882),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3834),
.A2(n_3875),
.B(n_3911),
.Y(n_3982)
);

HB1xp67_ASAP7_75t_L g3983 ( 
.A(n_3868),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3870),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3855),
.Y(n_3985)
);

OAI221xp5_ASAP7_75t_L g3986 ( 
.A1(n_3857),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3860),
.B(n_244),
.Y(n_3987)
);

OAI31xp33_ASAP7_75t_L g3988 ( 
.A1(n_3894),
.A2(n_247),
.A3(n_245),
.B(n_246),
.Y(n_3988)
);

NAND2xp33_ASAP7_75t_R g3989 ( 
.A(n_3862),
.B(n_246),
.Y(n_3989)
);

OAI22xp5_ASAP7_75t_L g3990 ( 
.A1(n_3904),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_3990)
);

AOI22xp5_ASAP7_75t_L g3991 ( 
.A1(n_3839),
.A2(n_251),
.B1(n_248),
.B2(n_249),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3849),
.Y(n_3992)
);

BUFx2_ASAP7_75t_L g3993 ( 
.A(n_3872),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3858),
.Y(n_3994)
);

NAND3xp33_ASAP7_75t_L g3995 ( 
.A(n_3851),
.B(n_251),
.C(n_252),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3878),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3895),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3863),
.Y(n_3998)
);

OAI221xp5_ASAP7_75t_L g3999 ( 
.A1(n_3925),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.C(n_255),
.Y(n_3999)
);

AND2x4_ASAP7_75t_L g4000 ( 
.A(n_3850),
.B(n_253),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3892),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3836),
.B(n_3837),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3915),
.B(n_254),
.Y(n_4003)
);

INVx1_ASAP7_75t_SL g4004 ( 
.A(n_3887),
.Y(n_4004)
);

NAND2x1p5_ASAP7_75t_L g4005 ( 
.A(n_3926),
.B(n_1280),
.Y(n_4005)
);

HB1xp67_ASAP7_75t_L g4006 ( 
.A(n_3884),
.Y(n_4006)
);

AOI33xp33_ASAP7_75t_L g4007 ( 
.A1(n_3871),
.A2(n_257),
.A3(n_260),
.B1(n_255),
.B2(n_256),
.B3(n_259),
.Y(n_4007)
);

OAI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3842),
.A2(n_259),
.B1(n_256),
.B2(n_257),
.Y(n_4008)
);

OR2x2_ASAP7_75t_L g4009 ( 
.A(n_3897),
.B(n_261),
.Y(n_4009)
);

OAI211xp5_ASAP7_75t_SL g4010 ( 
.A1(n_3902),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3840),
.Y(n_4011)
);

OR2x2_ASAP7_75t_L g4012 ( 
.A(n_3866),
.B(n_263),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3891),
.B(n_264),
.Y(n_4013)
);

OA21x2_ASAP7_75t_L g4014 ( 
.A1(n_3874),
.A2(n_264),
.B(n_266),
.Y(n_4014)
);

INVxp33_ASAP7_75t_L g4015 ( 
.A(n_3893),
.Y(n_4015)
);

INVx4_ASAP7_75t_SL g4016 ( 
.A(n_3905),
.Y(n_4016)
);

OAI33xp33_ASAP7_75t_L g4017 ( 
.A1(n_3922),
.A2(n_269),
.A3(n_271),
.B1(n_267),
.B2(n_268),
.B3(n_270),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3838),
.Y(n_4018)
);

OAI221xp5_ASAP7_75t_L g4019 ( 
.A1(n_3918),
.A2(n_270),
.B1(n_267),
.B2(n_268),
.C(n_271),
.Y(n_4019)
);

NOR3xp33_ASAP7_75t_SL g4020 ( 
.A(n_3918),
.B(n_272),
.C(n_273),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3838),
.Y(n_4021)
);

BUFx6f_ASAP7_75t_L g4022 ( 
.A(n_3841),
.Y(n_4022)
);

OAI31xp33_ASAP7_75t_L g4023 ( 
.A1(n_3918),
.A2(n_274),
.A3(n_272),
.B(n_273),
.Y(n_4023)
);

INVxp33_ASAP7_75t_L g4024 ( 
.A(n_3900),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_3890),
.Y(n_4025)
);

AOI221xp5_ASAP7_75t_L g4026 ( 
.A1(n_3918),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_4026)
);

OAI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3918),
.A2(n_279),
.B1(n_276),
.B2(n_278),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3888),
.B(n_278),
.Y(n_4028)
);

INVxp67_ASAP7_75t_L g4029 ( 
.A(n_3846),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3865),
.Y(n_4030)
);

AOI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3908),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3924),
.B(n_282),
.Y(n_4032)
);

OAI211xp5_ASAP7_75t_L g4033 ( 
.A1(n_3908),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_4033)
);

AND2x4_ASAP7_75t_L g4034 ( 
.A(n_3921),
.B(n_284),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3865),
.Y(n_4035)
);

OAI211xp5_ASAP7_75t_L g4036 ( 
.A1(n_3908),
.A2(n_289),
.B(n_285),
.C(n_287),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3921),
.B(n_285),
.Y(n_4037)
);

NOR2x1_ASAP7_75t_SL g4038 ( 
.A(n_3909),
.B(n_287),
.Y(n_4038)
);

INVxp67_ASAP7_75t_SL g4039 ( 
.A(n_3884),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_R g4040 ( 
.A(n_3890),
.B(n_290),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3838),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3838),
.Y(n_4042)
);

NAND2x1_ASAP7_75t_L g4043 ( 
.A(n_3865),
.B(n_291),
.Y(n_4043)
);

AOI22xp33_ASAP7_75t_L g4044 ( 
.A1(n_3908),
.A2(n_295),
.B1(n_291),
.B2(n_292),
.Y(n_4044)
);

HB1xp67_ASAP7_75t_L g4045 ( 
.A(n_3846),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3838),
.Y(n_4046)
);

OAI221xp5_ASAP7_75t_L g4047 ( 
.A1(n_3918),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_4047)
);

AND2x4_ASAP7_75t_L g4048 ( 
.A(n_3921),
.B(n_296),
.Y(n_4048)
);

AOI221xp5_ASAP7_75t_L g4049 ( 
.A1(n_3918),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.C(n_301),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_3890),
.Y(n_4050)
);

AOI221xp5_ASAP7_75t_L g4051 ( 
.A1(n_3918),
.A2(n_303),
.B1(n_299),
.B2(n_302),
.C(n_304),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3908),
.A2(n_305),
.B1(n_302),
.B2(n_304),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3888),
.B(n_306),
.Y(n_4053)
);

INVx1_ASAP7_75t_SL g4054 ( 
.A(n_3882),
.Y(n_4054)
);

OA21x2_ASAP7_75t_L g4055 ( 
.A1(n_3879),
.A2(n_307),
.B(n_308),
.Y(n_4055)
);

AOI222xp33_ASAP7_75t_L g4056 ( 
.A1(n_3918),
.A2(n_309),
.B1(n_313),
.B2(n_307),
.C1(n_308),
.C2(n_311),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3838),
.Y(n_4057)
);

A2O1A1Ixp33_ASAP7_75t_SL g4058 ( 
.A1(n_3918),
.A2(n_315),
.B(n_311),
.C(n_314),
.Y(n_4058)
);

AO21x2_ASAP7_75t_L g4059 ( 
.A1(n_3886),
.A2(n_314),
.B(n_316),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3838),
.Y(n_4060)
);

OAI211xp5_ASAP7_75t_SL g4061 ( 
.A1(n_3918),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3865),
.Y(n_4062)
);

AND2x6_ASAP7_75t_SL g4063 ( 
.A(n_3889),
.B(n_317),
.Y(n_4063)
);

OAI211xp5_ASAP7_75t_SL g4064 ( 
.A1(n_3918),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_4064)
);

INVx1_ASAP7_75t_SL g4065 ( 
.A(n_3882),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3838),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_3921),
.B(n_321),
.Y(n_4067)
);

OA21x2_ASAP7_75t_L g4068 ( 
.A1(n_3982),
.A2(n_4039),
.B(n_4001),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_3997),
.Y(n_4069)
);

INVx3_ASAP7_75t_L g4070 ( 
.A(n_4022),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_3993),
.B(n_322),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_3961),
.B(n_4045),
.Y(n_4072)
);

BUFx12f_ASAP7_75t_L g4073 ( 
.A(n_4025),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3938),
.B(n_323),
.Y(n_4074)
);

AND2x4_ASAP7_75t_L g4075 ( 
.A(n_4029),
.B(n_323),
.Y(n_4075)
);

INVxp67_ASAP7_75t_SL g4076 ( 
.A(n_4006),
.Y(n_4076)
);

INVx2_ASAP7_75t_SL g4077 ( 
.A(n_4022),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_SL g4078 ( 
.A1(n_4038),
.A2(n_324),
.B(n_325),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3996),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3951),
.Y(n_4080)
);

OA21x2_ASAP7_75t_L g4081 ( 
.A1(n_3936),
.A2(n_326),
.B(n_327),
.Y(n_4081)
);

OR2x6_ASAP7_75t_L g4082 ( 
.A(n_3977),
.B(n_326),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3939),
.Y(n_4083)
);

BUFx2_ASAP7_75t_L g4084 ( 
.A(n_3998),
.Y(n_4084)
);

OR2x2_ASAP7_75t_L g4085 ( 
.A(n_4011),
.B(n_327),
.Y(n_4085)
);

INVx3_ASAP7_75t_L g4086 ( 
.A(n_3935),
.Y(n_4086)
);

INVx4_ASAP7_75t_SL g4087 ( 
.A(n_3959),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3975),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3945),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_4030),
.Y(n_4090)
);

INVx3_ASAP7_75t_L g4091 ( 
.A(n_4035),
.Y(n_4091)
);

BUFx2_ASAP7_75t_L g4092 ( 
.A(n_4062),
.Y(n_4092)
);

AOI21xp33_ASAP7_75t_L g4093 ( 
.A1(n_4033),
.A2(n_328),
.B(n_330),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3971),
.Y(n_4094)
);

INVx1_ASAP7_75t_SL g4095 ( 
.A(n_4040),
.Y(n_4095)
);

NOR2x1p5_ASAP7_75t_L g4096 ( 
.A(n_3940),
.B(n_330),
.Y(n_4096)
);

AOI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_4036),
.A2(n_331),
.B(n_332),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3967),
.B(n_332),
.Y(n_4098)
);

OR2x6_ASAP7_75t_L g4099 ( 
.A(n_3974),
.B(n_333),
.Y(n_4099)
);

INVx2_ASAP7_75t_SL g4100 ( 
.A(n_4054),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3956),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3957),
.Y(n_4102)
);

INVx2_ASAP7_75t_L g4103 ( 
.A(n_3984),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3955),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_SL g4105 ( 
.A(n_3976),
.B(n_333),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_4065),
.B(n_334),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3983),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3985),
.B(n_335),
.Y(n_4108)
);

INVx1_ASAP7_75t_SL g4109 ( 
.A(n_4050),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4004),
.B(n_335),
.Y(n_4110)
);

AOI21x1_ASAP7_75t_L g4111 ( 
.A1(n_4043),
.A2(n_337),
.B(n_338),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_3994),
.B(n_3953),
.Y(n_4112)
);

AO21x1_ASAP7_75t_L g4113 ( 
.A1(n_3989),
.A2(n_337),
.B(n_338),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3937),
.Y(n_4114)
);

HB1xp67_ASAP7_75t_L g4115 ( 
.A(n_3992),
.Y(n_4115)
);

INVx4_ASAP7_75t_SL g4116 ( 
.A(n_3959),
.Y(n_4116)
);

OA21x2_ASAP7_75t_L g4117 ( 
.A1(n_3942),
.A2(n_339),
.B(n_340),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3948),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3949),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_4034),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4018),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4021),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3950),
.B(n_339),
.Y(n_4123)
);

BUFx8_ASAP7_75t_L g4124 ( 
.A(n_4003),
.Y(n_4124)
);

NAND3xp33_ASAP7_75t_SL g4125 ( 
.A(n_3952),
.B(n_340),
.C(n_341),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4041),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4042),
.Y(n_4127)
);

OA21x2_ASAP7_75t_L g4128 ( 
.A1(n_4046),
.A2(n_342),
.B(n_344),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_4057),
.Y(n_4129)
);

AND2x4_ASAP7_75t_SL g4130 ( 
.A(n_4048),
.B(n_342),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4060),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_4066),
.Y(n_4132)
);

NAND3xp33_ASAP7_75t_L g4133 ( 
.A(n_3933),
.B(n_344),
.C(n_345),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4009),
.Y(n_4134)
);

OA21x2_ASAP7_75t_L g4135 ( 
.A1(n_3962),
.A2(n_346),
.B(n_347),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3987),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3965),
.Y(n_4137)
);

HB1xp67_ASAP7_75t_L g4138 ( 
.A(n_3972),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4015),
.B(n_350),
.Y(n_4139)
);

INVx2_ASAP7_75t_SL g4140 ( 
.A(n_4016),
.Y(n_4140)
);

OAI21x1_ASAP7_75t_L g4141 ( 
.A1(n_3969),
.A2(n_351),
.B(n_352),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_4032),
.Y(n_4142)
);

OA21x2_ASAP7_75t_L g4143 ( 
.A1(n_3973),
.A2(n_353),
.B(n_355),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4000),
.Y(n_4144)
);

OAI21x1_ASAP7_75t_L g4145 ( 
.A1(n_3978),
.A2(n_4055),
.B(n_4053),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4028),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4014),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3979),
.B(n_355),
.Y(n_4148)
);

INVx5_ASAP7_75t_L g4149 ( 
.A(n_4063),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3963),
.Y(n_4150)
);

INVxp67_ASAP7_75t_L g4151 ( 
.A(n_3947),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4037),
.Y(n_4152)
);

INVx2_ASAP7_75t_SL g4153 ( 
.A(n_4016),
.Y(n_4153)
);

INVxp67_ASAP7_75t_SL g4154 ( 
.A(n_4067),
.Y(n_4154)
);

INVx1_ASAP7_75t_SL g4155 ( 
.A(n_4002),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_3968),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4059),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4012),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3995),
.Y(n_4159)
);

OA21x2_ASAP7_75t_L g4160 ( 
.A1(n_3958),
.A2(n_357),
.B(n_359),
.Y(n_4160)
);

OAI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_3934),
.A2(n_357),
.B(n_359),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_4013),
.Y(n_4162)
);

INVx3_ASAP7_75t_L g4163 ( 
.A(n_4005),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3954),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3946),
.B(n_360),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_4024),
.B(n_360),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4008),
.Y(n_4167)
);

AO21x2_ASAP7_75t_L g4168 ( 
.A1(n_4058),
.A2(n_361),
.B(n_362),
.Y(n_4168)
);

BUFx2_ASAP7_75t_L g4169 ( 
.A(n_4020),
.Y(n_4169)
);

OA21x2_ASAP7_75t_L g4170 ( 
.A1(n_3970),
.A2(n_361),
.B(n_363),
.Y(n_4170)
);

OAI21x1_ASAP7_75t_L g4171 ( 
.A1(n_3941),
.A2(n_363),
.B(n_365),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3944),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3966),
.Y(n_4173)
);

HB1xp67_ASAP7_75t_L g4174 ( 
.A(n_3999),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4007),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_3986),
.Y(n_4176)
);

INVx2_ASAP7_75t_SL g4177 ( 
.A(n_3990),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_3991),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_4019),
.Y(n_4179)
);

INVx2_ASAP7_75t_SL g4180 ( 
.A(n_3981),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4047),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3960),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4010),
.Y(n_4183)
);

INVx4_ASAP7_75t_SL g4184 ( 
.A(n_3943),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4027),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4017),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_3988),
.B(n_366),
.Y(n_4187)
);

INVx2_ASAP7_75t_L g4188 ( 
.A(n_4023),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4061),
.Y(n_4189)
);

OR2x2_ASAP7_75t_L g4190 ( 
.A(n_3964),
.B(n_4031),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4064),
.Y(n_4191)
);

INVxp67_ASAP7_75t_SL g4192 ( 
.A(n_3980),
.Y(n_4192)
);

BUFx3_ASAP7_75t_L g4193 ( 
.A(n_4056),
.Y(n_4193)
);

INVx4_ASAP7_75t_SL g4194 ( 
.A(n_3932),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4052),
.B(n_366),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_4044),
.B(n_367),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4026),
.B(n_4049),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_SL g4198 ( 
.A(n_4051),
.B(n_367),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4001),
.Y(n_4199)
);

NAND3xp33_ASAP7_75t_L g4200 ( 
.A(n_3938),
.B(n_368),
.C(n_369),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4001),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4001),
.Y(n_4202)
);

INVx2_ASAP7_75t_SL g4203 ( 
.A(n_4022),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4001),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4001),
.Y(n_4205)
);

BUFx2_ASAP7_75t_L g4206 ( 
.A(n_3961),
.Y(n_4206)
);

OAI21x1_ASAP7_75t_L g4207 ( 
.A1(n_3982),
.A2(n_368),
.B(n_369),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4001),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3961),
.B(n_370),
.Y(n_4209)
);

INVx4_ASAP7_75t_SL g4210 ( 
.A(n_3959),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_3997),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_3993),
.B(n_370),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4001),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4001),
.Y(n_4214)
);

AOI21x1_ASAP7_75t_L g4215 ( 
.A1(n_4043),
.A2(n_371),
.B(n_372),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4001),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3997),
.Y(n_4217)
);

INVx4_ASAP7_75t_SL g4218 ( 
.A(n_3959),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4001),
.Y(n_4219)
);

BUFx2_ASAP7_75t_L g4220 ( 
.A(n_3961),
.Y(n_4220)
);

INVx5_ASAP7_75t_L g4221 ( 
.A(n_3959),
.Y(n_4221)
);

AOI21x1_ASAP7_75t_L g4222 ( 
.A1(n_4043),
.A2(n_373),
.B(n_374),
.Y(n_4222)
);

OA21x2_ASAP7_75t_L g4223 ( 
.A1(n_3982),
.A2(n_373),
.B(n_374),
.Y(n_4223)
);

OAI21x1_ASAP7_75t_L g4224 ( 
.A1(n_3982),
.A2(n_375),
.B(n_376),
.Y(n_4224)
);

BUFx2_ASAP7_75t_L g4225 ( 
.A(n_3961),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4145),
.B(n_376),
.Y(n_4226)
);

NAND2x1p5_ASAP7_75t_L g4227 ( 
.A(n_4206),
.B(n_377),
.Y(n_4227)
);

AND2x2_ASAP7_75t_L g4228 ( 
.A(n_4072),
.B(n_378),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4084),
.B(n_379),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4159),
.B(n_4146),
.Y(n_4230)
);

AND2x2_ASAP7_75t_L g4231 ( 
.A(n_4140),
.B(n_379),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_L g4232 ( 
.A1(n_4193),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_4232)
);

INVx2_ASAP7_75t_SL g4233 ( 
.A(n_4153),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4136),
.B(n_380),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4220),
.B(n_381),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4225),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4080),
.Y(n_4237)
);

INVx4_ASAP7_75t_L g4238 ( 
.A(n_4073),
.Y(n_4238)
);

NAND3xp33_ASAP7_75t_L g4239 ( 
.A(n_4149),
.B(n_382),
.C(n_383),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4088),
.Y(n_4240)
);

HB1xp67_ASAP7_75t_L g4241 ( 
.A(n_4223),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4118),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4091),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4121),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4158),
.B(n_383),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4138),
.B(n_384),
.Y(n_4246)
);

AOI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_4074),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4122),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4154),
.B(n_385),
.Y(n_4249)
);

BUFx2_ASAP7_75t_L g4250 ( 
.A(n_4076),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4147),
.B(n_386),
.Y(n_4251)
);

AND2x2_ASAP7_75t_L g4252 ( 
.A(n_4155),
.B(n_387),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4134),
.B(n_387),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4131),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4199),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_4142),
.B(n_388),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4094),
.B(n_4157),
.Y(n_4257)
);

NOR2xp67_ASAP7_75t_L g4258 ( 
.A(n_4221),
.B(n_388),
.Y(n_4258)
);

NAND2x1p5_ASAP7_75t_L g4259 ( 
.A(n_4100),
.B(n_389),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4164),
.B(n_389),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4092),
.B(n_390),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4150),
.B(n_390),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4201),
.Y(n_4263)
);

AND2x4_ASAP7_75t_L g4264 ( 
.A(n_4077),
.B(n_391),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4202),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4152),
.B(n_392),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4204),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4162),
.B(n_393),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_4083),
.B(n_394),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4089),
.B(n_394),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4156),
.B(n_395),
.Y(n_4271)
);

AND2x4_ASAP7_75t_SL g4272 ( 
.A(n_4082),
.B(n_395),
.Y(n_4272)
);

CKINVDCx20_ASAP7_75t_R g4273 ( 
.A(n_4124),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4090),
.B(n_396),
.Y(n_4274)
);

AND2x4_ASAP7_75t_L g4275 ( 
.A(n_4203),
.B(n_396),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4205),
.Y(n_4276)
);

OR2x2_ASAP7_75t_L g4277 ( 
.A(n_4107),
.B(n_397),
.Y(n_4277)
);

AOI22xp5_ASAP7_75t_L g4278 ( 
.A1(n_4194),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4208),
.Y(n_4279)
);

NOR3xp33_ASAP7_75t_L g4280 ( 
.A(n_4200),
.B(n_399),
.C(n_400),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4101),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_SL g4282 ( 
.A(n_4149),
.B(n_400),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4085),
.B(n_401),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4070),
.B(n_4086),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4102),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4213),
.Y(n_4286)
);

INVx3_ASAP7_75t_L g4287 ( 
.A(n_4120),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4104),
.Y(n_4288)
);

INVx2_ASAP7_75t_SL g4289 ( 
.A(n_4221),
.Y(n_4289)
);

INVxp67_ASAP7_75t_L g4290 ( 
.A(n_4135),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4144),
.B(n_402),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4112),
.B(n_403),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4137),
.B(n_404),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4214),
.Y(n_4294)
);

INVx2_ASAP7_75t_SL g4295 ( 
.A(n_4120),
.Y(n_4295)
);

HB1xp67_ASAP7_75t_L g4296 ( 
.A(n_4115),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4079),
.B(n_404),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4151),
.B(n_405),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4143),
.B(n_405),
.Y(n_4299)
);

AND2x4_ASAP7_75t_SL g4300 ( 
.A(n_4099),
.B(n_406),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_SL g4301 ( 
.A(n_4113),
.B(n_406),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_4114),
.B(n_407),
.Y(n_4302)
);

AND2x4_ASAP7_75t_L g4303 ( 
.A(n_4087),
.B(n_408),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4174),
.B(n_408),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4119),
.B(n_409),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4216),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4126),
.Y(n_4307)
);

INVxp67_ASAP7_75t_L g4308 ( 
.A(n_4169),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4127),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4105),
.B(n_409),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4123),
.B(n_410),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4129),
.B(n_410),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4219),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4132),
.B(n_411),
.Y(n_4314)
);

OR2x2_ASAP7_75t_L g4315 ( 
.A(n_4103),
.B(n_412),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_4108),
.B(n_413),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4069),
.B(n_414),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4211),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4217),
.B(n_414),
.Y(n_4319)
);

INVxp67_ASAP7_75t_L g4320 ( 
.A(n_4176),
.Y(n_4320)
);

OR2x2_ASAP7_75t_L g4321 ( 
.A(n_4167),
.B(n_415),
.Y(n_4321)
);

AND2x4_ASAP7_75t_L g4322 ( 
.A(n_4116),
.B(n_416),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4210),
.B(n_417),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4218),
.B(n_418),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4139),
.B(n_418),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4117),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4192),
.B(n_419),
.Y(n_4327)
);

NOR2x1_ASAP7_75t_L g4328 ( 
.A(n_4078),
.B(n_419),
.Y(n_4328)
);

INVx3_ASAP7_75t_L g4329 ( 
.A(n_4075),
.Y(n_4329)
);

INVx1_ASAP7_75t_SL g4330 ( 
.A(n_4095),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4128),
.Y(n_4331)
);

AND2x4_ASAP7_75t_L g4332 ( 
.A(n_4163),
.B(n_421),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4098),
.B(n_421),
.Y(n_4333)
);

OR2x2_ASAP7_75t_L g4334 ( 
.A(n_4209),
.B(n_422),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4172),
.B(n_423),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4071),
.B(n_423),
.Y(n_4336)
);

NOR2xp33_ASAP7_75t_L g4337 ( 
.A(n_4179),
.B(n_424),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4081),
.Y(n_4338)
);

INVx3_ASAP7_75t_L g4339 ( 
.A(n_4109),
.Y(n_4339)
);

AND2x2_ASAP7_75t_L g4340 ( 
.A(n_4212),
.B(n_424),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4173),
.B(n_425),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4207),
.Y(n_4342)
);

AND2x2_ASAP7_75t_L g4343 ( 
.A(n_4068),
.B(n_425),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4178),
.B(n_427),
.Y(n_4344)
);

INVx4_ASAP7_75t_L g4345 ( 
.A(n_4130),
.Y(n_4345)
);

AND2x4_ASAP7_75t_SL g4346 ( 
.A(n_4106),
.B(n_428),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4224),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4141),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4110),
.Y(n_4349)
);

OR2x2_ASAP7_75t_L g4350 ( 
.A(n_4185),
.B(n_428),
.Y(n_4350)
);

AOI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4198),
.A2(n_4197),
.B1(n_4188),
.B2(n_4133),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4177),
.B(n_429),
.Y(n_4352)
);

NOR2x1p5_ASAP7_75t_L g4353 ( 
.A(n_4125),
.B(n_429),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4166),
.B(n_430),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4180),
.B(n_430),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4111),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4181),
.B(n_4184),
.Y(n_4357)
);

NAND3xp33_ASAP7_75t_L g4358 ( 
.A(n_4189),
.B(n_431),
.C(n_432),
.Y(n_4358)
);

INVx1_ASAP7_75t_SL g4359 ( 
.A(n_4148),
.Y(n_4359)
);

NAND2x1_ASAP7_75t_L g4360 ( 
.A(n_4160),
.B(n_432),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4186),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4182),
.B(n_4175),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4183),
.B(n_433),
.Y(n_4363)
);

INVxp67_ASAP7_75t_L g4364 ( 
.A(n_4191),
.Y(n_4364)
);

INVx1_ASAP7_75t_SL g4365 ( 
.A(n_4187),
.Y(n_4365)
);

NAND5xp2_ASAP7_75t_L g4366 ( 
.A(n_4097),
.B(n_436),
.C(n_434),
.D(n_435),
.E(n_437),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4170),
.B(n_434),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4096),
.B(n_435),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4215),
.B(n_438),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4222),
.B(n_438),
.Y(n_4370)
);

AOI21xp33_ASAP7_75t_SL g4371 ( 
.A1(n_4093),
.A2(n_439),
.B(n_442),
.Y(n_4371)
);

NAND2xp33_ASAP7_75t_L g4372 ( 
.A(n_4165),
.B(n_439),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4168),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4190),
.Y(n_4374)
);

AND2x4_ASAP7_75t_L g4375 ( 
.A(n_4171),
.B(n_443),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4196),
.B(n_444),
.Y(n_4376)
);

NAND4xp25_ASAP7_75t_SL g4377 ( 
.A(n_4195),
.B(n_447),
.C(n_445),
.D(n_446),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_4161),
.B(n_447),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4145),
.B(n_448),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4072),
.B(n_448),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4145),
.B(n_449),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4145),
.B(n_450),
.Y(n_4382)
);

OR2x2_ASAP7_75t_L g4383 ( 
.A(n_4147),
.B(n_450),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4080),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4145),
.B(n_451),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4084),
.Y(n_4386)
);

OAI22xp5_ASAP7_75t_SL g4387 ( 
.A1(n_4149),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4145),
.B(n_453),
.Y(n_4388)
);

OAI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_4200),
.A2(n_454),
.B(n_455),
.Y(n_4389)
);

OAI31xp33_ASAP7_75t_SL g4390 ( 
.A1(n_4200),
.A2(n_458),
.A3(n_455),
.B(n_456),
.Y(n_4390)
);

OR2x2_ASAP7_75t_L g4391 ( 
.A(n_4147),
.B(n_456),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4080),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4072),
.B(n_459),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4080),
.Y(n_4394)
);

OR2x2_ASAP7_75t_L g4395 ( 
.A(n_4147),
.B(n_460),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4072),
.B(n_461),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4072),
.B(n_461),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4080),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4072),
.B(n_462),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4072),
.B(n_462),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4072),
.B(n_463),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4072),
.B(n_463),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4072),
.B(n_464),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4080),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4080),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4145),
.B(n_464),
.Y(n_4406)
);

OR2x2_ASAP7_75t_L g4407 ( 
.A(n_4147),
.B(n_465),
.Y(n_4407)
);

AOI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4074),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_4408)
);

INVxp67_ASAP7_75t_SL g4409 ( 
.A(n_4206),
.Y(n_4409)
);

OR2x2_ASAP7_75t_L g4410 ( 
.A(n_4147),
.B(n_466),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4080),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_4072),
.B(n_468),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4084),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4080),
.Y(n_4414)
);

INVx2_ASAP7_75t_SL g4415 ( 
.A(n_4140),
.Y(n_4415)
);

AND2x4_ASAP7_75t_L g4416 ( 
.A(n_4140),
.B(n_468),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4080),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4080),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_4072),
.B(n_469),
.Y(n_4419)
);

HB1xp67_ASAP7_75t_L g4420 ( 
.A(n_4206),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4080),
.Y(n_4421)
);

NAND3xp33_ASAP7_75t_L g4422 ( 
.A(n_4149),
.B(n_469),
.C(n_470),
.Y(n_4422)
);

OR2x2_ASAP7_75t_L g4423 ( 
.A(n_4147),
.B(n_470),
.Y(n_4423)
);

OAI33xp33_ASAP7_75t_L g4424 ( 
.A1(n_4074),
.A2(n_473),
.A3(n_475),
.B1(n_471),
.B2(n_472),
.B3(n_474),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4145),
.B(n_471),
.Y(n_4425)
);

BUFx3_ASAP7_75t_L g4426 ( 
.A(n_4073),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4080),
.Y(n_4427)
);

NOR2xp33_ASAP7_75t_SL g4428 ( 
.A(n_4149),
.B(n_473),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4080),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4072),
.B(n_474),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4145),
.B(n_477),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4080),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4080),
.Y(n_4433)
);

OAI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_4200),
.A2(n_477),
.B(n_478),
.Y(n_4434)
);

OR2x2_ASAP7_75t_L g4435 ( 
.A(n_4147),
.B(n_478),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4072),
.B(n_479),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4080),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4084),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4080),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4237),
.Y(n_4440)
);

NAND2x1p5_ASAP7_75t_L g4441 ( 
.A(n_4250),
.B(n_479),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4240),
.Y(n_4442)
);

NOR2xp33_ASAP7_75t_SL g4443 ( 
.A(n_4238),
.B(n_480),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4242),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4244),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4248),
.Y(n_4446)
);

INVxp67_ASAP7_75t_L g4447 ( 
.A(n_4428),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4289),
.B(n_480),
.Y(n_4448)
);

HB1xp67_ASAP7_75t_L g4449 ( 
.A(n_4250),
.Y(n_4449)
);

AOI31xp33_ASAP7_75t_L g4450 ( 
.A1(n_4328),
.A2(n_4301),
.A3(n_4434),
.B(n_4389),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4361),
.B(n_481),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4254),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4255),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4263),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4233),
.B(n_481),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4265),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4267),
.Y(n_4457)
);

OR2x2_ASAP7_75t_L g4458 ( 
.A(n_4374),
.B(n_482),
.Y(n_4458)
);

BUFx2_ASAP7_75t_L g4459 ( 
.A(n_4409),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4308),
.B(n_482),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4415),
.B(n_483),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4276),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4386),
.B(n_484),
.Y(n_4463)
);

NAND2x1p5_ASAP7_75t_L g4464 ( 
.A(n_4360),
.B(n_484),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4279),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4365),
.B(n_485),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4286),
.Y(n_4467)
);

NOR2x1_ASAP7_75t_L g4468 ( 
.A(n_4258),
.B(n_486),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4320),
.B(n_487),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4294),
.Y(n_4470)
);

NOR2x1_ASAP7_75t_L g4471 ( 
.A(n_4343),
.B(n_487),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4290),
.B(n_488),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4413),
.B(n_488),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4287),
.Y(n_4474)
);

AND2x4_ASAP7_75t_L g4475 ( 
.A(n_4284),
.B(n_4295),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4438),
.B(n_489),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4306),
.Y(n_4477)
);

INVx3_ASAP7_75t_SL g4478 ( 
.A(n_4273),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4313),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4330),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4384),
.Y(n_4481)
);

HB1xp67_ASAP7_75t_L g4482 ( 
.A(n_4420),
.Y(n_4482)
);

NAND2xp33_ASAP7_75t_SL g4483 ( 
.A(n_4387),
.B(n_490),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4392),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4394),
.Y(n_4485)
);

AND2x4_ASAP7_75t_SL g4486 ( 
.A(n_4345),
.B(n_490),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4243),
.B(n_491),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_4426),
.B(n_4364),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4236),
.B(n_491),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4398),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4359),
.B(n_492),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4342),
.B(n_492),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4349),
.B(n_493),
.Y(n_4493)
);

OAI21xp33_ASAP7_75t_L g4494 ( 
.A1(n_4390),
.A2(n_493),
.B(n_494),
.Y(n_4494)
);

INVxp67_ASAP7_75t_L g4495 ( 
.A(n_4357),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4347),
.B(n_495),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4404),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4405),
.Y(n_4498)
);

INVxp67_ASAP7_75t_L g4499 ( 
.A(n_4241),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4411),
.Y(n_4500)
);

NAND4xp25_ASAP7_75t_L g4501 ( 
.A(n_4366),
.B(n_498),
.C(n_496),
.D(n_497),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4230),
.B(n_498),
.Y(n_4502)
);

OR2x6_ASAP7_75t_L g4503 ( 
.A(n_4303),
.B(n_499),
.Y(n_4503)
);

AND2x4_ASAP7_75t_L g4504 ( 
.A(n_4339),
.B(n_499),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4414),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4417),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4418),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4338),
.B(n_500),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4329),
.B(n_500),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4348),
.B(n_501),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4421),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4281),
.Y(n_4512)
);

OR2x2_ASAP7_75t_L g4513 ( 
.A(n_4326),
.B(n_501),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4373),
.B(n_502),
.Y(n_4514)
);

OR2x2_ASAP7_75t_L g4515 ( 
.A(n_4331),
.B(n_502),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4427),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4226),
.B(n_503),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4228),
.B(n_503),
.Y(n_4518)
);

OR2x2_ASAP7_75t_L g4519 ( 
.A(n_4285),
.B(n_504),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4379),
.B(n_504),
.Y(n_4520)
);

O2A1O1Ixp5_ASAP7_75t_L g4521 ( 
.A1(n_4282),
.A2(n_508),
.B(n_505),
.C(n_506),
.Y(n_4521)
);

OR2x2_ASAP7_75t_L g4522 ( 
.A(n_4288),
.B(n_505),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4429),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4307),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4381),
.B(n_508),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4382),
.B(n_509),
.Y(n_4526)
);

NAND2x1p5_ASAP7_75t_L g4527 ( 
.A(n_4235),
.B(n_509),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4432),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4385),
.B(n_511),
.Y(n_4529)
);

INVxp67_ASAP7_75t_SL g4530 ( 
.A(n_4227),
.Y(n_4530)
);

AND2x4_ASAP7_75t_SL g4531 ( 
.A(n_4322),
.B(n_511),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4380),
.B(n_512),
.Y(n_4532)
);

INVx2_ASAP7_75t_SL g4533 ( 
.A(n_4416),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_4257),
.B(n_513),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4393),
.B(n_514),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4309),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_4323),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4388),
.B(n_514),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4433),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4396),
.B(n_515),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4315),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4437),
.Y(n_4542)
);

NAND3x1_ASAP7_75t_L g4543 ( 
.A(n_4351),
.B(n_515),
.C(n_516),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4406),
.B(n_516),
.Y(n_4544)
);

OR2x2_ASAP7_75t_L g4545 ( 
.A(n_4318),
.B(n_517),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4425),
.B(n_517),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4397),
.B(n_518),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4399),
.B(n_519),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4439),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4431),
.B(n_519),
.Y(n_4550)
);

AND2x2_ASAP7_75t_L g4551 ( 
.A(n_4436),
.B(n_520),
.Y(n_4551)
);

NOR2xp33_ASAP7_75t_L g4552 ( 
.A(n_4304),
.B(n_520),
.Y(n_4552)
);

INVx1_ASAP7_75t_SL g4553 ( 
.A(n_4324),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4296),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4383),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_4362),
.B(n_521),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4391),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4367),
.B(n_521),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4395),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4407),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4400),
.B(n_522),
.Y(n_4561)
);

INVx2_ASAP7_75t_L g4562 ( 
.A(n_4256),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4410),
.Y(n_4563)
);

OR2x2_ASAP7_75t_L g4564 ( 
.A(n_4356),
.B(n_522),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4423),
.Y(n_4565)
);

OR2x2_ASAP7_75t_L g4566 ( 
.A(n_4271),
.B(n_523),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4401),
.B(n_523),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4435),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4430),
.B(n_524),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4297),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4402),
.B(n_524),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4403),
.B(n_525),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4412),
.B(n_4419),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4317),
.Y(n_4574)
);

OR2x2_ASAP7_75t_L g4575 ( 
.A(n_4321),
.B(n_525),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_4251),
.B(n_526),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4277),
.Y(n_4577)
);

OR2x2_ASAP7_75t_L g4578 ( 
.A(n_4253),
.B(n_526),
.Y(n_4578)
);

OR2x2_ASAP7_75t_L g4579 ( 
.A(n_4350),
.B(n_4352),
.Y(n_4579)
);

INVxp67_ASAP7_75t_SL g4580 ( 
.A(n_4259),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4341),
.B(n_527),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4319),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4261),
.B(n_4249),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4252),
.B(n_527),
.Y(n_4584)
);

AO21x1_ASAP7_75t_L g4585 ( 
.A1(n_4327),
.A2(n_528),
.B(n_529),
.Y(n_4585)
);

INVx2_ASAP7_75t_SL g4586 ( 
.A(n_4231),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4292),
.B(n_4229),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4302),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_4264),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4305),
.Y(n_4590)
);

OR2x2_ASAP7_75t_L g4591 ( 
.A(n_4260),
.B(n_4234),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4449),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4482),
.Y(n_4593)
);

BUFx3_ASAP7_75t_L g4594 ( 
.A(n_4478),
.Y(n_4594)
);

OR2x2_ASAP7_75t_L g4595 ( 
.A(n_4459),
.B(n_4344),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4475),
.Y(n_4596)
);

BUFx2_ASAP7_75t_L g4597 ( 
.A(n_4580),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4553),
.B(n_4355),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4440),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4442),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4444),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4537),
.B(n_4335),
.Y(n_4602)
);

BUFx3_ASAP7_75t_L g4603 ( 
.A(n_4486),
.Y(n_4603)
);

NAND2x1_ASAP7_75t_SL g4604 ( 
.A(n_4468),
.B(n_4278),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4445),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4495),
.B(n_4298),
.Y(n_4606)
);

AOI22xp33_ASAP7_75t_L g4607 ( 
.A1(n_4494),
.A2(n_4280),
.B1(n_4372),
.B2(n_4353),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_4533),
.Y(n_4608)
);

HB1xp67_ASAP7_75t_L g4609 ( 
.A(n_4480),
.Y(n_4609)
);

OR2x2_ASAP7_75t_L g4610 ( 
.A(n_4565),
.B(n_4283),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4474),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4446),
.Y(n_4612)
);

AOI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4501),
.A2(n_4377),
.B1(n_4378),
.B2(n_4337),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4586),
.B(n_4471),
.Y(n_4614)
);

INVxp67_ASAP7_75t_L g4615 ( 
.A(n_4530),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4588),
.B(n_4363),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4589),
.Y(n_4617)
);

INVx2_ASAP7_75t_SL g4618 ( 
.A(n_4531),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4452),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4573),
.B(n_4246),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4579),
.B(n_4334),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4453),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4587),
.B(n_4293),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4488),
.B(n_4291),
.Y(n_4624)
);

OR2x2_ASAP7_75t_L g4625 ( 
.A(n_4577),
.B(n_4299),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4570),
.B(n_4245),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4574),
.B(n_4582),
.Y(n_4627)
);

INVx1_ASAP7_75t_SL g4628 ( 
.A(n_4483),
.Y(n_4628)
);

AOI22xp33_ASAP7_75t_L g4629 ( 
.A1(n_4541),
.A2(n_4424),
.B1(n_4232),
.B2(n_4408),
.Y(n_4629)
);

INVx1_ASAP7_75t_SL g4630 ( 
.A(n_4503),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4454),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4441),
.Y(n_4632)
);

NOR2xp33_ASAP7_75t_L g4633 ( 
.A(n_4447),
.B(n_4316),
.Y(n_4633)
);

AND3x1_ASAP7_75t_L g4634 ( 
.A(n_4443),
.B(n_4247),
.C(n_4562),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4519),
.Y(n_4635)
);

HB1xp67_ASAP7_75t_L g4636 ( 
.A(n_4499),
.Y(n_4636)
);

AND3x1_ASAP7_75t_L g4637 ( 
.A(n_4552),
.B(n_4368),
.C(n_4310),
.Y(n_4637)
);

BUFx2_ASAP7_75t_L g4638 ( 
.A(n_4464),
.Y(n_4638)
);

AOI22xp33_ASAP7_75t_L g4639 ( 
.A1(n_4590),
.A2(n_4422),
.B1(n_4239),
.B2(n_4358),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4522),
.Y(n_4640)
);

INVx3_ASAP7_75t_SL g4641 ( 
.A(n_4503),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4555),
.B(n_4354),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4456),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4450),
.B(n_4312),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4557),
.B(n_4325),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4559),
.B(n_4268),
.Y(n_4646)
);

INVx3_ASAP7_75t_L g4647 ( 
.A(n_4504),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4560),
.B(n_4314),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4457),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4563),
.B(n_4336),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4527),
.Y(n_4651)
);

AOI22xp33_ASAP7_75t_L g4652 ( 
.A1(n_4568),
.A2(n_4375),
.B1(n_4376),
.B2(n_4369),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4462),
.Y(n_4653)
);

AND2x2_ASAP7_75t_L g4654 ( 
.A(n_4493),
.B(n_4554),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4465),
.Y(n_4655)
);

INVx4_ASAP7_75t_L g4656 ( 
.A(n_4448),
.Y(n_4656)
);

OAI21xp33_ASAP7_75t_L g4657 ( 
.A1(n_4508),
.A2(n_4371),
.B(n_4300),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4583),
.B(n_4333),
.Y(n_4658)
);

AND2x4_ASAP7_75t_L g4659 ( 
.A(n_4455),
.B(n_4332),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4463),
.B(n_4340),
.Y(n_4660)
);

INVxp67_ASAP7_75t_SL g4661 ( 
.A(n_4543),
.Y(n_4661)
);

INVx1_ASAP7_75t_SL g4662 ( 
.A(n_4461),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4473),
.B(n_4262),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4591),
.B(n_4311),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4545),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4512),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4524),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4476),
.B(n_4489),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4536),
.Y(n_4669)
);

NAND3xp33_ASAP7_75t_L g4670 ( 
.A(n_4521),
.B(n_4370),
.C(n_4270),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4467),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4509),
.Y(n_4672)
);

AND3x1_ASAP7_75t_L g4673 ( 
.A(n_4472),
.B(n_4266),
.C(n_4269),
.Y(n_4673)
);

HB1xp67_ASAP7_75t_L g4674 ( 
.A(n_4564),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_L g4675 ( 
.A(n_4585),
.B(n_4510),
.Y(n_4675)
);

NOR2xp33_ASAP7_75t_L g4676 ( 
.A(n_4451),
.B(n_4346),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4491),
.B(n_4274),
.Y(n_4677)
);

HB1xp67_ASAP7_75t_L g4678 ( 
.A(n_4513),
.Y(n_4678)
);

INVxp67_ASAP7_75t_L g4679 ( 
.A(n_4515),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4636),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4610),
.Y(n_4681)
);

OAI22xp5_ASAP7_75t_L g4682 ( 
.A1(n_4634),
.A2(n_4514),
.B1(n_4492),
.B2(n_4496),
.Y(n_4682)
);

NAND4xp25_ASAP7_75t_L g4683 ( 
.A(n_4644),
.B(n_4460),
.C(n_4556),
.D(n_4520),
.Y(n_4683)
);

AOI311xp33_ASAP7_75t_L g4684 ( 
.A1(n_4661),
.A2(n_4470),
.A3(n_4481),
.B(n_4479),
.C(n_4477),
.Y(n_4684)
);

AND2x4_ASAP7_75t_L g4685 ( 
.A(n_4594),
.B(n_4484),
.Y(n_4685)
);

OR2x2_ASAP7_75t_L g4686 ( 
.A(n_4675),
.B(n_4502),
.Y(n_4686)
);

AO22x1_ASAP7_75t_L g4687 ( 
.A1(n_4628),
.A2(n_4641),
.B1(n_4651),
.B2(n_4638),
.Y(n_4687)
);

AOI221xp5_ASAP7_75t_L g4688 ( 
.A1(n_4593),
.A2(n_4526),
.B1(n_4529),
.B2(n_4525),
.C(n_4517),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4592),
.Y(n_4689)
);

OAI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4604),
.A2(n_4607),
.B(n_4639),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4603),
.Y(n_4691)
);

OAI22xp5_ASAP7_75t_L g4692 ( 
.A1(n_4629),
.A2(n_4534),
.B1(n_4544),
.B2(n_4538),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4678),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4609),
.Y(n_4694)
);

AND2x4_ASAP7_75t_SL g4695 ( 
.A(n_4659),
.B(n_4275),
.Y(n_4695)
);

XOR2x2_ASAP7_75t_L g4696 ( 
.A(n_4637),
.B(n_4546),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4674),
.Y(n_4697)
);

OAI21xp5_ASAP7_75t_SL g4698 ( 
.A1(n_4613),
.A2(n_4550),
.B(n_4272),
.Y(n_4698)
);

NOR2xp33_ASAP7_75t_L g4699 ( 
.A(n_4656),
.B(n_4458),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4630),
.B(n_4597),
.Y(n_4700)
);

AOI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4615),
.A2(n_4490),
.B1(n_4497),
.B2(n_4485),
.Y(n_4701)
);

AOI221xp5_ASAP7_75t_L g4702 ( 
.A1(n_4679),
.A2(n_4498),
.B1(n_4506),
.B2(n_4505),
.C(n_4500),
.Y(n_4702)
);

XNOR2xp5_ASAP7_75t_L g4703 ( 
.A(n_4673),
.B(n_4584),
.Y(n_4703)
);

AOI21xp5_ASAP7_75t_L g4704 ( 
.A1(n_4614),
.A2(n_4558),
.B(n_4576),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4620),
.B(n_4487),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4670),
.A2(n_4469),
.B1(n_4466),
.B2(n_4566),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4596),
.B(n_4518),
.Y(n_4707)
);

HB1xp67_ASAP7_75t_L g4708 ( 
.A(n_4598),
.Y(n_4708)
);

OAI21xp33_ASAP7_75t_L g4709 ( 
.A1(n_4608),
.A2(n_4511),
.B(n_4507),
.Y(n_4709)
);

NAND4xp25_ASAP7_75t_L g4710 ( 
.A(n_4617),
.B(n_4581),
.C(n_4578),
.D(n_4575),
.Y(n_4710)
);

OAI22xp33_ASAP7_75t_L g4711 ( 
.A1(n_4595),
.A2(n_4523),
.B1(n_4528),
.B2(n_4516),
.Y(n_4711)
);

OAI211xp5_ASAP7_75t_SL g4712 ( 
.A1(n_4657),
.A2(n_4542),
.B(n_4549),
.C(n_4539),
.Y(n_4712)
);

NAND3xp33_ASAP7_75t_L g4713 ( 
.A(n_4611),
.B(n_4535),
.C(n_4532),
.Y(n_4713)
);

OAI211xp5_ASAP7_75t_L g4714 ( 
.A1(n_4627),
.A2(n_4547),
.B(n_4548),
.C(n_4540),
.Y(n_4714)
);

NOR3xp33_ASAP7_75t_L g4715 ( 
.A(n_4633),
.B(n_4561),
.C(n_4551),
.Y(n_4715)
);

OR2x2_ASAP7_75t_L g4716 ( 
.A(n_4662),
.B(n_4567),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_4647),
.B(n_4569),
.Y(n_4717)
);

INVxp67_ASAP7_75t_L g4718 ( 
.A(n_4618),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4602),
.Y(n_4719)
);

AOI21xp33_ASAP7_75t_L g4720 ( 
.A1(n_4625),
.A2(n_4572),
.B(n_4571),
.Y(n_4720)
);

AOI221xp5_ASAP7_75t_L g4721 ( 
.A1(n_4599),
.A2(n_531),
.B1(n_528),
.B2(n_530),
.C(n_532),
.Y(n_4721)
);

AOI21xp33_ASAP7_75t_SL g4722 ( 
.A1(n_4632),
.A2(n_530),
.B(n_531),
.Y(n_4722)
);

NOR2xp33_ASAP7_75t_L g4723 ( 
.A(n_4624),
.B(n_532),
.Y(n_4723)
);

INVxp67_ASAP7_75t_L g4724 ( 
.A(n_4660),
.Y(n_4724)
);

INVxp33_ASAP7_75t_L g4725 ( 
.A(n_4676),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4642),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_4606),
.Y(n_4727)
);

NOR2xp33_ASAP7_75t_L g4728 ( 
.A(n_4672),
.B(n_4668),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4621),
.B(n_533),
.Y(n_4729)
);

O2A1O1Ixp33_ASAP7_75t_L g4730 ( 
.A1(n_4600),
.A2(n_536),
.B(n_534),
.C(n_535),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4623),
.Y(n_4731)
);

INVx2_ASAP7_75t_SL g4732 ( 
.A(n_4663),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4677),
.B(n_534),
.Y(n_4733)
);

AOI211xp5_ASAP7_75t_L g4734 ( 
.A1(n_4658),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4650),
.B(n_4645),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4648),
.A2(n_537),
.B(n_538),
.Y(n_4736)
);

OAI32xp33_ASAP7_75t_L g4737 ( 
.A1(n_4665),
.A2(n_543),
.A3(n_539),
.B1(n_541),
.B2(n_544),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4654),
.B(n_539),
.Y(n_4738)
);

OAI22xp5_ASAP7_75t_L g4739 ( 
.A1(n_4652),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_4646),
.B(n_545),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4635),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4640),
.B(n_546),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_4616),
.Y(n_4743)
);

AOI222xp33_ASAP7_75t_L g4744 ( 
.A1(n_4626),
.A2(n_550),
.B1(n_552),
.B2(n_547),
.C1(n_549),
.C2(n_551),
.Y(n_4744)
);

XNOR2xp5_ASAP7_75t_L g4745 ( 
.A(n_4664),
.B(n_549),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4708),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4718),
.B(n_4666),
.Y(n_4747)
);

INVx2_ASAP7_75t_L g4748 ( 
.A(n_4691),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4703),
.B(n_4667),
.Y(n_4749)
);

INVx3_ASAP7_75t_L g4750 ( 
.A(n_4695),
.Y(n_4750)
);

AOI222xp33_ASAP7_75t_L g4751 ( 
.A1(n_4690),
.A2(n_4619),
.B1(n_4605),
.B2(n_4622),
.C1(n_4612),
.C2(n_4601),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4680),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4707),
.B(n_4669),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_SL g4754 ( 
.A(n_4685),
.B(n_4631),
.Y(n_4754)
);

AND2x4_ASAP7_75t_SL g4755 ( 
.A(n_4685),
.B(n_4643),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4732),
.B(n_4649),
.Y(n_4756)
);

OAI21xp33_ASAP7_75t_L g4757 ( 
.A1(n_4700),
.A2(n_4655),
.B(n_4653),
.Y(n_4757)
);

NOR2xp33_ASAP7_75t_L g4758 ( 
.A(n_4725),
.B(n_4671),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4716),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4686),
.B(n_550),
.Y(n_4760)
);

INVxp67_ASAP7_75t_L g4761 ( 
.A(n_4717),
.Y(n_4761)
);

NOR2xp33_ASAP7_75t_L g4762 ( 
.A(n_4714),
.B(n_553),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4731),
.B(n_553),
.Y(n_4763)
);

INVxp67_ASAP7_75t_L g4764 ( 
.A(n_4728),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4694),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4727),
.B(n_554),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4697),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_SL g4768 ( 
.A(n_4715),
.B(n_554),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4719),
.B(n_555),
.Y(n_4769)
);

INVx1_ASAP7_75t_SL g4770 ( 
.A(n_4687),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4724),
.B(n_4736),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4726),
.B(n_555),
.Y(n_4772)
);

NOR2x1_ASAP7_75t_L g4773 ( 
.A(n_4729),
.B(n_556),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4693),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4681),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4744),
.B(n_556),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4740),
.Y(n_4777)
);

INVx1_ASAP7_75t_SL g4778 ( 
.A(n_4735),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4733),
.Y(n_4779)
);

AOI22xp33_ASAP7_75t_L g4780 ( 
.A1(n_4696),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4689),
.Y(n_4781)
);

NOR2xp33_ASAP7_75t_SL g4782 ( 
.A(n_4699),
.B(n_559),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4710),
.B(n_560),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4723),
.B(n_561),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4704),
.B(n_562),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4683),
.B(n_562),
.Y(n_4786)
);

OR2x2_ASAP7_75t_L g4787 ( 
.A(n_4705),
.B(n_563),
.Y(n_4787)
);

O2A1O1Ixp33_ASAP7_75t_L g4788 ( 
.A1(n_4770),
.A2(n_4722),
.B(n_4739),
.C(n_4682),
.Y(n_4788)
);

AOI221xp5_ASAP7_75t_L g4789 ( 
.A1(n_4757),
.A2(n_4711),
.B1(n_4692),
.B2(n_4712),
.C(n_4702),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_SL g4790 ( 
.A1(n_4785),
.A2(n_4730),
.B(n_4745),
.Y(n_4790)
);

NAND4xp25_ASAP7_75t_L g4791 ( 
.A(n_4749),
.B(n_4684),
.C(n_4701),
.D(n_4741),
.Y(n_4791)
);

AOI211xp5_ASAP7_75t_SL g4792 ( 
.A1(n_4764),
.A2(n_4709),
.B(n_4743),
.C(n_4734),
.Y(n_4792)
);

AOI21xp33_ASAP7_75t_SL g4793 ( 
.A1(n_4746),
.A2(n_4706),
.B(n_4720),
.Y(n_4793)
);

AOI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4762),
.A2(n_4698),
.B1(n_4713),
.B2(n_4688),
.Y(n_4794)
);

AOI221x1_ASAP7_75t_L g4795 ( 
.A1(n_4783),
.A2(n_4742),
.B1(n_4738),
.B2(n_4737),
.C(n_4721),
.Y(n_4795)
);

A2O1A1Ixp33_ASAP7_75t_L g4796 ( 
.A1(n_4780),
.A2(n_565),
.B(n_563),
.C(n_564),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_SL g4797 ( 
.A(n_4750),
.B(n_565),
.Y(n_4797)
);

OAI321xp33_ASAP7_75t_L g4798 ( 
.A1(n_4761),
.A2(n_569),
.A3(n_572),
.B1(n_566),
.B2(n_568),
.C(n_570),
.Y(n_4798)
);

BUFx2_ASAP7_75t_L g4799 ( 
.A(n_4773),
.Y(n_4799)
);

AOI211xp5_ASAP7_75t_L g4800 ( 
.A1(n_4776),
.A2(n_572),
.B(n_566),
.C(n_568),
.Y(n_4800)
);

OAI221xp5_ASAP7_75t_L g4801 ( 
.A1(n_4751),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.C(n_576),
.Y(n_4801)
);

NAND3xp33_ASAP7_75t_L g4802 ( 
.A(n_4754),
.B(n_573),
.C(n_575),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4755),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4748),
.B(n_576),
.Y(n_4804)
);

AOI221xp5_ASAP7_75t_L g4805 ( 
.A1(n_4758),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_4805)
);

NOR3xp33_ASAP7_75t_L g4806 ( 
.A(n_4771),
.B(n_4747),
.C(n_4759),
.Y(n_4806)
);

AOI22xp5_ASAP7_75t_L g4807 ( 
.A1(n_4778),
.A2(n_4768),
.B1(n_4753),
.B2(n_4777),
.Y(n_4807)
);

AOI221xp5_ASAP7_75t_L g4808 ( 
.A1(n_4752),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_4808)
);

AOI22xp5_ASAP7_75t_L g4809 ( 
.A1(n_4775),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_4809)
);

AND4x1_ASAP7_75t_L g4810 ( 
.A(n_4782),
.B(n_583),
.C(n_581),
.D(n_582),
.Y(n_4810)
);

OAI211xp5_ASAP7_75t_L g4811 ( 
.A1(n_4756),
.A2(n_587),
.B(n_585),
.C(n_586),
.Y(n_4811)
);

NOR2xp33_ASAP7_75t_L g4812 ( 
.A(n_4786),
.B(n_586),
.Y(n_4812)
);

OAI211xp5_ASAP7_75t_SL g4813 ( 
.A1(n_4779),
.A2(n_589),
.B(n_587),
.C(n_588),
.Y(n_4813)
);

A2O1A1Ixp33_ASAP7_75t_L g4814 ( 
.A1(n_4760),
.A2(n_590),
.B(n_588),
.C(n_589),
.Y(n_4814)
);

AOI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4784),
.A2(n_590),
.B(n_592),
.Y(n_4815)
);

NOR2x1_ASAP7_75t_L g4816 ( 
.A(n_4766),
.B(n_592),
.Y(n_4816)
);

OAI21xp33_ASAP7_75t_L g4817 ( 
.A1(n_4767),
.A2(n_593),
.B(n_594),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4763),
.Y(n_4818)
);

O2A1O1Ixp33_ASAP7_75t_SL g4819 ( 
.A1(n_4765),
.A2(n_4774),
.B(n_4781),
.C(n_4787),
.Y(n_4819)
);

AOI221x1_ASAP7_75t_L g4820 ( 
.A1(n_4769),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.C(n_596),
.Y(n_4820)
);

NAND4xp25_ASAP7_75t_SL g4821 ( 
.A(n_4772),
.B(n_597),
.C(n_595),
.D(n_596),
.Y(n_4821)
);

OAI321xp33_ASAP7_75t_L g4822 ( 
.A1(n_4749),
.A2(n_599),
.A3(n_602),
.B1(n_597),
.B2(n_598),
.C(n_600),
.Y(n_4822)
);

O2A1O1Ixp33_ASAP7_75t_L g4823 ( 
.A1(n_4770),
.A2(n_602),
.B(n_598),
.C(n_600),
.Y(n_4823)
);

AOI222xp33_ASAP7_75t_L g4824 ( 
.A1(n_4770),
.A2(n_607),
.B1(n_609),
.B2(n_603),
.C1(n_606),
.C2(n_608),
.Y(n_4824)
);

OA21x2_ASAP7_75t_L g4825 ( 
.A1(n_4780),
.A2(n_603),
.B(n_606),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4746),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4750),
.B(n_608),
.Y(n_4827)
);

AOI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4785),
.A2(n_609),
.B(n_611),
.Y(n_4828)
);

AOI22xp33_ASAP7_75t_SL g4829 ( 
.A1(n_4799),
.A2(n_4803),
.B1(n_4801),
.B2(n_4825),
.Y(n_4829)
);

NOR2xp67_ASAP7_75t_L g4830 ( 
.A(n_4807),
.B(n_611),
.Y(n_4830)
);

AOI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_4789),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_4831)
);

OAI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4788),
.A2(n_4823),
.B(n_4792),
.Y(n_4832)
);

AOI21xp33_ASAP7_75t_SL g4833 ( 
.A1(n_4825),
.A2(n_613),
.B(n_614),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4816),
.Y(n_4834)
);

OAI22xp5_ASAP7_75t_L g4835 ( 
.A1(n_4794),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4827),
.B(n_4824),
.Y(n_4836)
);

OAI311xp33_ASAP7_75t_L g4837 ( 
.A1(n_4791),
.A2(n_618),
.A3(n_615),
.B1(n_616),
.C1(n_619),
.Y(n_4837)
);

AOI22xp5_ASAP7_75t_L g4838 ( 
.A1(n_4806),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_4838)
);

OAI221xp5_ASAP7_75t_L g4839 ( 
.A1(n_4793),
.A2(n_623),
.B1(n_620),
.B2(n_621),
.C(n_624),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4818),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4826),
.Y(n_4841)
);

AOI21xp5_ASAP7_75t_L g4842 ( 
.A1(n_4790),
.A2(n_623),
.B(n_624),
.Y(n_4842)
);

OAI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_4800),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4812),
.A2(n_631),
.B1(n_626),
.B2(n_628),
.Y(n_4844)
);

AOI221x1_ASAP7_75t_L g4845 ( 
.A1(n_4828),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.C(n_634),
.Y(n_4845)
);

NOR2xp33_ASAP7_75t_L g4846 ( 
.A(n_4797),
.B(n_632),
.Y(n_4846)
);

NAND2xp33_ASAP7_75t_SL g4847 ( 
.A(n_4804),
.B(n_633),
.Y(n_4847)
);

NOR2x1p5_ASAP7_75t_L g4848 ( 
.A(n_4802),
.B(n_635),
.Y(n_4848)
);

AOI211xp5_ASAP7_75t_L g4849 ( 
.A1(n_4819),
.A2(n_639),
.B(n_636),
.C(n_637),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4815),
.B(n_639),
.Y(n_4850)
);

AOI222xp33_ASAP7_75t_L g4851 ( 
.A1(n_4805),
.A2(n_640),
.B1(n_641),
.B2(n_642),
.C1(n_643),
.C2(n_644),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4810),
.Y(n_4852)
);

OAI211xp5_ASAP7_75t_L g4853 ( 
.A1(n_4795),
.A2(n_642),
.B(n_640),
.C(n_641),
.Y(n_4853)
);

OAI21xp5_ASAP7_75t_L g4854 ( 
.A1(n_4796),
.A2(n_643),
.B(n_644),
.Y(n_4854)
);

CKINVDCx20_ASAP7_75t_R g4855 ( 
.A(n_4809),
.Y(n_4855)
);

NAND2x1_ASAP7_75t_L g4856 ( 
.A(n_4834),
.B(n_4822),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4852),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4829),
.B(n_4820),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4840),
.Y(n_4859)
);

INVx1_ASAP7_75t_SL g4860 ( 
.A(n_4847),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4846),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4841),
.Y(n_4862)
);

INVx3_ASAP7_75t_L g4863 ( 
.A(n_4850),
.Y(n_4863)
);

XNOR2x1_ASAP7_75t_L g4864 ( 
.A(n_4832),
.B(n_4831),
.Y(n_4864)
);

NOR2x1p5_ASAP7_75t_L g4865 ( 
.A(n_4836),
.B(n_4821),
.Y(n_4865)
);

AOI32xp33_ASAP7_75t_L g4866 ( 
.A1(n_4849),
.A2(n_4813),
.A3(n_4798),
.B1(n_4808),
.B2(n_4817),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4833),
.B(n_4814),
.Y(n_4867)
);

AND2x2_ASAP7_75t_L g4868 ( 
.A(n_4848),
.B(n_4811),
.Y(n_4868)
);

NOR2xp33_ASAP7_75t_L g4869 ( 
.A(n_4853),
.B(n_645),
.Y(n_4869)
);

XNOR2x1_ASAP7_75t_L g4870 ( 
.A(n_4864),
.B(n_4865),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4869),
.B(n_4830),
.Y(n_4871)
);

HB1xp67_ASAP7_75t_L g4872 ( 
.A(n_4856),
.Y(n_4872)
);

AOI22xp5_ASAP7_75t_L g4873 ( 
.A1(n_4857),
.A2(n_4855),
.B1(n_4835),
.B2(n_4839),
.Y(n_4873)
);

NOR2xp67_ASAP7_75t_L g4874 ( 
.A(n_4859),
.B(n_4842),
.Y(n_4874)
);

NOR2xp33_ASAP7_75t_R g4875 ( 
.A(n_4863),
.B(n_4844),
.Y(n_4875)
);

OAI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_4858),
.A2(n_4837),
.B(n_4845),
.Y(n_4876)
);

NAND4xp75_ASAP7_75t_L g4877 ( 
.A(n_4874),
.B(n_4862),
.C(n_4861),
.D(n_4867),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4872),
.B(n_4868),
.Y(n_4878)
);

OAI221xp5_ASAP7_75t_L g4879 ( 
.A1(n_4876),
.A2(n_4866),
.B1(n_4860),
.B2(n_4838),
.C(n_4854),
.Y(n_4879)
);

NOR3xp33_ASAP7_75t_L g4880 ( 
.A(n_4879),
.B(n_4871),
.C(n_4873),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_SL g4881 ( 
.A(n_4878),
.B(n_4851),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4877),
.Y(n_4882)
);

BUFx2_ASAP7_75t_L g4883 ( 
.A(n_4882),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4880),
.B(n_4870),
.Y(n_4884)
);

AOI322xp5_ASAP7_75t_L g4885 ( 
.A1(n_4881),
.A2(n_4875),
.A3(n_4843),
.B1(n_647),
.B2(n_648),
.C1(n_649),
.C2(n_650),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4884),
.Y(n_4886)
);

XNOR2x1_ASAP7_75t_L g4887 ( 
.A(n_4885),
.B(n_645),
.Y(n_4887)
);

HB1xp67_ASAP7_75t_L g4888 ( 
.A(n_4883),
.Y(n_4888)
);

AOI22xp5_ASAP7_75t_L g4889 ( 
.A1(n_4888),
.A2(n_649),
.B1(n_646),
.B2(n_648),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_SL g4890 ( 
.A(n_4886),
.B(n_646),
.Y(n_4890)
);

INVxp67_ASAP7_75t_SL g4891 ( 
.A(n_4887),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4888),
.Y(n_4892)
);

NAND3xp33_ASAP7_75t_L g4893 ( 
.A(n_4892),
.B(n_651),
.C(n_652),
.Y(n_4893)
);

AOI21xp33_ASAP7_75t_L g4894 ( 
.A1(n_4891),
.A2(n_651),
.B(n_652),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_SL g4895 ( 
.A(n_4889),
.B(n_654),
.Y(n_4895)
);

OAI22xp5_ASAP7_75t_SL g4896 ( 
.A1(n_4893),
.A2(n_4890),
.B1(n_657),
.B2(n_655),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4895),
.Y(n_4897)
);

AOI221xp5_ASAP7_75t_L g4898 ( 
.A1(n_4896),
.A2(n_4897),
.B1(n_4894),
.B2(n_657),
.C(n_655),
.Y(n_4898)
);

AOI22xp33_ASAP7_75t_R g4899 ( 
.A1(n_4898),
.A2(n_659),
.B1(n_656),
.B2(n_658),
.Y(n_4899)
);

AOI22xp33_ASAP7_75t_L g4900 ( 
.A1(n_4899),
.A2(n_661),
.B1(n_656),
.B2(n_660),
.Y(n_4900)
);

AOI22xp5_ASAP7_75t_L g4901 ( 
.A1(n_4900),
.A2(n_662),
.B1(n_660),
.B2(n_661),
.Y(n_4901)
);

AOI211xp5_ASAP7_75t_L g4902 ( 
.A1(n_4901),
.A2(n_664),
.B(n_662),
.C(n_663),
.Y(n_4902)
);


endmodule