module fake_netlist_6_4608_n_1124 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1124);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1124;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_468;
wire n_372;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_143),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_146),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_41),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_165),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_37),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_106),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_104),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_74),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_26),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_62),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_8),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_132),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_59),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_127),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_88),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_9),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_70),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_126),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_112),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_148),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_142),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_107),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_199),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_200),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_137),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_85),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_2),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_274),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_0),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_206),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_248),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_219),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_266),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_209),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_227),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_206),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_249),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_206),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_210),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_211),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_240),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_228),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_310),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_276),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_287),
.B(n_230),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_284),
.A2(n_273),
.B1(n_214),
.B2(n_217),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_252),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_288),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g350 ( 
.A1(n_285),
.A2(n_261),
.B(n_218),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_270),
.B1(n_269),
.B2(n_264),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_286),
.A2(n_263),
.B1(n_262),
.B2(n_259),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_213),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_240),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_293),
.B(n_220),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_289),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_222),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_231),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_243),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_323),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_320),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_243),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

AO21x2_ASAP7_75t_L g382 ( 
.A1(n_346),
.A2(n_307),
.B(n_306),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_361),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_322),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_308),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_337),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_377),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_342),
.A2(n_313),
.B1(n_309),
.B2(n_304),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

NOR2x1p5_ASAP7_75t_L g417 ( 
.A(n_336),
.B(n_304),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_318),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_330),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_309),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_297),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_324),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_364),
.A2(n_243),
.B(n_233),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_31),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_232),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_352),
.B(n_320),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_234),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_335),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_357),
.B(n_354),
.Y(n_440)
);

AO21x2_ASAP7_75t_L g441 ( 
.A1(n_345),
.A2(n_238),
.B(n_237),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_350),
.A2(n_245),
.B(n_241),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_330),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_341),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_347),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

NOR2x1p5_ASAP7_75t_L g450 ( 
.A(n_339),
.B(n_250),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_368),
.B(n_251),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_339),
.B(n_299),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_337),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_452),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_349),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_371),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

XNOR2x2_ASAP7_75t_L g466 ( 
.A(n_396),
.B(n_377),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

INVx4_ASAP7_75t_SL g470 ( 
.A(n_430),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_449),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_382),
.B(n_350),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_348),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_382),
.B(n_384),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_424),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_382),
.B(n_350),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_398),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_366),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_349),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_432),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_399),
.B(n_280),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_356),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_351),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_420),
.B(n_351),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_366),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_362),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_362),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_410),
.B(n_350),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_417),
.B(n_283),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_393),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_401),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_401),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_386),
.B(n_378),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_386),
.B(n_374),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_452),
.B(n_368),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_399),
.B(n_359),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_421),
.B(n_363),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_441),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_431),
.B(n_368),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_441),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_450),
.B(n_253),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_408),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_408),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_441),
.B(n_359),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_445),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

XOR2x2_ASAP7_75t_L g530 ( 
.A(n_442),
.B(n_359),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_450),
.B(n_367),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_437),
.A2(n_368),
.B(n_380),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_428),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_453),
.B(n_368),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_400),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_437),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_464),
.B(n_412),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_467),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_506),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_412),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

AND2x2_ASAP7_75t_SL g547 ( 
.A(n_525),
.B(n_430),
.Y(n_547)
);

OAI221xp5_ASAP7_75t_L g548 ( 
.A1(n_479),
.A2(n_462),
.B1(n_488),
.B2(n_456),
.C(n_475),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_478),
.A2(n_430),
.B1(n_416),
.B2(n_418),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_412),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_416),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_457),
.B(n_416),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_487),
.B(n_445),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_458),
.B(n_459),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_478),
.A2(n_430),
.B1(n_418),
.B2(n_385),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_496),
.A2(n_430),
.B1(n_452),
.B2(n_418),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_460),
.B(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_487),
.B(n_445),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_471),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_463),
.B(n_394),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_476),
.Y(n_562)
);

AND2x2_ASAP7_75t_SL g563 ( 
.A(n_533),
.B(n_438),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_495),
.B(n_367),
.Y(n_564)
);

OAI221xp5_ASAP7_75t_L g565 ( 
.A1(n_474),
.A2(n_369),
.B1(n_375),
.B2(n_373),
.C(n_254),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_470),
.B(n_445),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_470),
.B(n_448),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_480),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_499),
.A2(n_444),
.B1(n_446),
.B2(n_438),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

NOR3xp33_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_477),
.C(n_531),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_394),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_466),
.B(n_369),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_497),
.A2(n_446),
.B1(n_447),
.B2(n_444),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_489),
.B(n_394),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_497),
.B(n_375),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_500),
.B(n_394),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_501),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_395),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_470),
.B(n_448),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_503),
.A2(n_442),
.B1(n_451),
.B2(n_447),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_484),
.B(n_448),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_484),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_516),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_414),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_473),
.B(n_448),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_532),
.B(n_395),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_516),
.B(n_395),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_541),
.B(n_395),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_473),
.B(n_414),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_490),
.B(n_517),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_481),
.B(n_454),
.Y(n_594)
);

NOR2x1p5_ASAP7_75t_L g595 ( 
.A(n_481),
.B(n_255),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

NOR2x1p5_ASAP7_75t_L g597 ( 
.A(n_505),
.B(n_257),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_504),
.B(n_454),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_494),
.B(n_405),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_483),
.Y(n_600)
);

O2A1O1Ixp5_ASAP7_75t_L g601 ( 
.A1(n_518),
.A2(n_429),
.B(n_436),
.C(n_451),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_482),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_493),
.A2(n_376),
.B1(n_383),
.B2(n_385),
.C(n_390),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_504),
.B(n_454),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_539),
.B(n_405),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_521),
.B(n_376),
.Y(n_608)
);

NAND2x1p5_ASAP7_75t_L g609 ( 
.A(n_507),
.B(n_409),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_546),
.B(n_509),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_569),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

CKINVDCx14_ASAP7_75t_R g614 ( 
.A(n_602),
.Y(n_614)
);

NOR2x1_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_498),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_548),
.B(n_522),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_547),
.A2(n_513),
.B1(n_519),
.B2(n_514),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_520),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_586),
.B(n_523),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_585),
.B(n_530),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_564),
.B(n_578),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_577),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_524),
.Y(n_624)
);

NOR2x2_ASAP7_75t_L g625 ( 
.A(n_543),
.B(n_436),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_461),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_610),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_SL g629 ( 
.A(n_593),
.B(n_536),
.C(n_535),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_574),
.B(n_526),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_549),
.B(n_528),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_608),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_529),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_596),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_580),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_554),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_547),
.B(n_534),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_556),
.B(n_537),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_597),
.B(n_372),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_542),
.B(n_538),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_609),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_545),
.B(n_512),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_550),
.B(n_512),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_572),
.B(n_405),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_560),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_600),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_609),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_562),
.A2(n_429),
.B1(n_376),
.B2(n_414),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_552),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_604),
.B(n_376),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_595),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_568),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_603),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_606),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_587),
.B(n_589),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_591),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_565),
.A2(n_397),
.B(n_383),
.C(n_390),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_599),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_SL g664 ( 
.A(n_555),
.B(n_392),
.C(n_391),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_573),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_391),
.B1(n_392),
.B2(n_397),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_579),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_584),
.B(n_414),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_647),
.A2(n_583),
.B(n_588),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_637),
.B(n_590),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_L g674 ( 
.A(n_616),
.B(n_584),
.C(n_551),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_647),
.A2(n_594),
.B(n_588),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_660),
.A2(n_601),
.B(n_598),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_660),
.A2(n_663),
.B(n_645),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_632),
.A2(n_555),
.B1(n_570),
.B2(n_575),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_630),
.A2(n_607),
.B(n_605),
.C(n_598),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_631),
.A2(n_592),
.B(n_594),
.Y(n_680)
);

OAI21x1_ASAP7_75t_SL g681 ( 
.A1(n_617),
.A2(n_400),
.B(n_409),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_663),
.A2(n_605),
.B(n_559),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_644),
.A2(n_559),
.B(n_553),
.Y(n_683)
);

AO31x2_ASAP7_75t_L g684 ( 
.A1(n_644),
.A2(n_400),
.A3(n_413),
.B(n_409),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_613),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_645),
.A2(n_553),
.B(n_566),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_643),
.A2(n_567),
.B(n_566),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_617),
.A2(n_653),
.B(n_633),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_642),
.A2(n_582),
.B(n_567),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_629),
.A2(n_582),
.B(n_405),
.C(n_434),
.Y(n_690)
);

AO21x1_ASAP7_75t_L g691 ( 
.A1(n_651),
.A2(n_413),
.B(n_409),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_643),
.A2(n_434),
.B(n_419),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_622),
.B(n_0),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_652),
.A2(n_434),
.B(n_419),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_623),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_625),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_618),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_632),
.B(n_454),
.Y(n_698)
);

NOR2x1_ASAP7_75t_L g699 ( 
.A(n_650),
.B(n_419),
.Y(n_699)
);

NOR2x1_ASAP7_75t_SL g700 ( 
.A(n_669),
.B(n_388),
.Y(n_700)
);

AO221x1_ASAP7_75t_L g701 ( 
.A1(n_665),
.A2(n_666),
.B1(n_650),
.B2(n_640),
.C(n_648),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_419),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_646),
.B(n_640),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_642),
.A2(n_414),
.B(n_413),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_626),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_638),
.A2(n_413),
.B(n_406),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_434),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_668),
.A2(n_406),
.B(n_388),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_640),
.B(n_388),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_648),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_670),
.B(n_2),
.Y(n_711)
);

BUFx4_ASAP7_75t_SL g712 ( 
.A(n_654),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_614),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_661),
.A2(n_406),
.B(n_388),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_662),
.A2(n_406),
.B(n_388),
.C(n_5),
.Y(n_715)
);

AO31x2_ASAP7_75t_L g716 ( 
.A1(n_634),
.A2(n_365),
.A3(n_406),
.B(n_388),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_661),
.A2(n_406),
.B(n_33),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_SL g718 ( 
.A1(n_620),
.A2(n_655),
.B(n_656),
.C(n_657),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_620),
.B(n_3),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_619),
.A2(n_34),
.B(n_32),
.Y(n_720)
);

OAI21x1_ASAP7_75t_SL g721 ( 
.A1(n_634),
.A2(n_39),
.B(n_36),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_627),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_619),
.A2(n_43),
.B(n_40),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_615),
.B(n_3),
.Y(n_724)
);

AOI222xp33_ASAP7_75t_L g725 ( 
.A1(n_621),
.A2(n_365),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_628),
.A2(n_365),
.A3(n_10),
.B(n_11),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_667),
.A2(n_45),
.B(n_44),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_646),
.B(n_659),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_635),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_674),
.A2(n_641),
.B(n_626),
.C(n_648),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_677),
.A2(n_664),
.B(n_667),
.Y(n_731)
);

AO31x2_ASAP7_75t_L g732 ( 
.A1(n_691),
.A2(n_649),
.A3(n_639),
.B(n_669),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_728),
.B(n_665),
.Y(n_733)
);

OAI22x1_ASAP7_75t_L g734 ( 
.A1(n_696),
.A2(n_658),
.B1(n_639),
.B2(n_665),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_685),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_666),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_703),
.B(n_666),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_639),
.Y(n_738)
);

AOI221xp5_ASAP7_75t_L g739 ( 
.A1(n_688),
.A2(n_4),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_697),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_722),
.B(n_669),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_719),
.B(n_711),
.Y(n_742)
);

AOI22x1_ASAP7_75t_L g743 ( 
.A1(n_725),
.A2(n_639),
.B1(n_611),
.B2(n_13),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_679),
.A2(n_680),
.B(n_689),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_729),
.B(n_47),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_704),
.A2(n_611),
.B(n_365),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_683),
.A2(n_611),
.B(n_365),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_696),
.B(n_611),
.Y(n_748)
);

AOI221x1_ASAP7_75t_L g749 ( 
.A1(n_715),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_672),
.Y(n_750)
);

AO31x2_ASAP7_75t_L g751 ( 
.A1(n_690),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_695),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_SL g753 ( 
.A(n_698),
.B(n_15),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_724),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_754)
);

AO31x2_ASAP7_75t_L g755 ( 
.A1(n_700),
.A2(n_17),
.A3(n_18),
.B(n_19),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_718),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_722),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_714),
.A2(n_49),
.B(n_48),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_705),
.B(n_702),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_710),
.Y(n_760)
);

AO31x2_ASAP7_75t_L g761 ( 
.A1(n_708),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_676),
.A2(n_671),
.B(n_682),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_706),
.A2(n_51),
.B(n_50),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_705),
.B(n_20),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_678),
.A2(n_675),
.B(n_694),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_678),
.A2(n_205),
.B(n_123),
.Y(n_766)
);

OAI22x1_ASAP7_75t_L g767 ( 
.A1(n_709),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_707),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_701),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_717),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_710),
.B(n_24),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_699),
.B(n_27),
.Y(n_772)
);

AO32x2_ASAP7_75t_L g773 ( 
.A1(n_726),
.A2(n_27),
.A3(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_773)
);

AOI21xp33_ASAP7_75t_L g774 ( 
.A1(n_681),
.A2(n_28),
.B(n_30),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_686),
.A2(n_52),
.B(n_56),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_726),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_699),
.B(n_57),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_720),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_726),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_712),
.B1(n_721),
.B2(n_687),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_727),
.A2(n_692),
.B(n_723),
.Y(n_781)
);

BUFx2_ASAP7_75t_SL g782 ( 
.A(n_716),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_684),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_684),
.B(n_204),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_684),
.A2(n_58),
.B(n_60),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_716),
.A2(n_61),
.B(n_63),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_L g787 ( 
.A1(n_716),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_677),
.A2(n_68),
.B(n_69),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_674),
.B(n_72),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

AO31x2_ASAP7_75t_L g791 ( 
.A1(n_691),
.A2(n_73),
.A3(n_75),
.B(n_76),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_685),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_679),
.A2(n_203),
.B(n_78),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_790),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_743),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_760),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_736),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_752),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_739),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_742),
.B(n_84),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_735),
.Y(n_803)
);

BUFx4f_ASAP7_75t_SL g804 ( 
.A(n_737),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_792),
.Y(n_805)
);

CKINVDCx11_ASAP7_75t_R g806 ( 
.A(n_780),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_730),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_SL g808 ( 
.A1(n_766),
.A2(n_794),
.B1(n_775),
.B2(n_744),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_741),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_SL g810 ( 
.A1(n_789),
.A2(n_90),
.B(n_91),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_793),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_740),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_SL g813 ( 
.A1(n_765),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_757),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_753),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_815)
);

CKINVDCx11_ASAP7_75t_R g816 ( 
.A(n_769),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_734),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_776),
.Y(n_818)
);

BUFx4f_ASAP7_75t_SL g819 ( 
.A(n_771),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_733),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_768),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_754),
.A2(n_767),
.B1(n_738),
.B2(n_774),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_745),
.A2(n_103),
.B1(n_105),
.B2(n_108),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_748),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_764),
.Y(n_825)
);

INVx6_ASAP7_75t_L g826 ( 
.A(n_759),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_770),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_827)
);

BUFx4f_ASAP7_75t_SL g828 ( 
.A(n_778),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_779),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_772),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_830)
);

INVx3_ASAP7_75t_SL g831 ( 
.A(n_781),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_777),
.A2(n_763),
.B1(n_756),
.B2(n_784),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_749),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_761),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_755),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_751),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_781),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_773),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_788),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_782),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_747),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_751),
.Y(n_842)
);

CKINVDCx6p67_ASAP7_75t_R g843 ( 
.A(n_755),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_761),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_746),
.A2(n_785),
.B1(n_731),
.B2(n_758),
.Y(n_845)
);

INVx8_ASAP7_75t_L g846 ( 
.A(n_755),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_786),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_783),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_761),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_762),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_773),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_773),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_791),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_787),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_796),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_828),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_837),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_795),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_829),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_803),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_811),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_834),
.Y(n_866)
);

CKINVDCx6p67_ASAP7_75t_R g867 ( 
.A(n_816),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_795),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_820),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_809),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_844),
.A2(n_853),
.B(n_836),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_809),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_826),
.Y(n_873)
);

CKINVDCx11_ASAP7_75t_R g874 ( 
.A(n_814),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_835),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_795),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_826),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_825),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_820),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_842),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_820),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_824),
.B(n_732),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_842),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_852),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_845),
.A2(n_732),
.B(n_141),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_831),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_846),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_846),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_847),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_843),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_833),
.A2(n_808),
.B1(n_827),
.B2(n_841),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_849),
.B(n_851),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_799),
.B(n_140),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_838),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_838),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_798),
.B(n_147),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_812),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

AO21x2_ASAP7_75t_L g899 ( 
.A1(n_848),
.A2(n_149),
.B(n_150),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_884),
.B(n_840),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_855),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_886),
.B(n_854),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_892),
.A2(n_806),
.B1(n_801),
.B2(n_813),
.Y(n_903)
);

OA21x2_ASAP7_75t_L g904 ( 
.A1(n_871),
.A2(n_832),
.B(n_822),
.Y(n_904)
);

AO21x2_ASAP7_75t_L g905 ( 
.A1(n_871),
.A2(n_817),
.B(n_807),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_886),
.B(n_854),
.Y(n_906)
);

CKINVDCx6p67_ASAP7_75t_R g907 ( 
.A(n_867),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_878),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_870),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_870),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_859),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_866),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_884),
.B(n_840),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_890),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_866),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_858),
.B(n_847),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_888),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_859),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_855),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_858),
.B(n_894),
.Y(n_920)
);

AO21x2_ASAP7_75t_L g921 ( 
.A1(n_880),
.A2(n_802),
.B(n_823),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_861),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_861),
.Y(n_923)
);

AND2x2_ASAP7_75t_SL g924 ( 
.A(n_892),
.B(n_797),
.Y(n_924)
);

OAI211xp5_ASAP7_75t_SL g925 ( 
.A1(n_891),
.A2(n_815),
.B(n_830),
.C(n_810),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_880),
.A2(n_839),
.B(n_804),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_883),
.A2(n_850),
.B(n_819),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_882),
.B(n_151),
.Y(n_928)
);

CKINVDCx8_ASAP7_75t_R g929 ( 
.A(n_907),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_912),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_920),
.B(n_894),
.Y(n_931)
);

OAI211xp5_ASAP7_75t_L g932 ( 
.A1(n_903),
.A2(n_895),
.B(n_885),
.C(n_890),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_920),
.B(n_908),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_914),
.B(n_888),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_902),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_919),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_918),
.B(n_872),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_919),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_912),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_914),
.B(n_885),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_924),
.A2(n_899),
.B1(n_881),
.B2(n_873),
.Y(n_942)
);

NOR2x1_ASAP7_75t_L g943 ( 
.A(n_902),
.B(n_868),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_909),
.B(n_885),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_910),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_923),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_917),
.B(n_885),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_911),
.B(n_856),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_917),
.B(n_883),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_923),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_923),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_917),
.B(n_887),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_930),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_937),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_943),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_929),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_934),
.B(n_902),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_937),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_941),
.A2(n_898),
.B(n_915),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_950),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_934),
.B(n_902),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_930),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_948),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_931),
.B(n_941),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_931),
.B(n_936),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_948),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_936),
.B(n_902),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_950),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_963),
.B(n_938),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_956),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_956),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_966),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_964),
.B(n_933),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_959),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_964),
.B(n_953),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_957),
.B(n_935),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_957),
.B(n_935),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_955),
.B(n_947),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_953),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_962),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_971),
.B(n_959),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_970),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

NAND2x1_ASAP7_75t_SL g984 ( 
.A(n_978),
.B(n_967),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_976),
.B(n_961),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_979),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_965),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_969),
.B(n_965),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_983),
.B(n_977),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_907),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_982),
.B(n_929),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_986),
.Y(n_992)
);

OAI22xp33_ASAP7_75t_L g993 ( 
.A1(n_988),
.A2(n_955),
.B1(n_975),
.B2(n_973),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_987),
.B(n_975),
.Y(n_994)
);

AO221x2_ASAP7_75t_L g995 ( 
.A1(n_984),
.A2(n_981),
.B1(n_867),
.B2(n_980),
.C(n_974),
.Y(n_995)
);

AO221x2_ASAP7_75t_L g996 ( 
.A1(n_981),
.A2(n_974),
.B1(n_973),
.B2(n_874),
.C(n_860),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_992),
.B(n_985),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_989),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_990),
.B(n_978),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_994),
.B(n_978),
.Y(n_1000)
);

INVxp67_ASAP7_75t_SL g1001 ( 
.A(n_993),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_991),
.B(n_967),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_995),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_996),
.B(n_961),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_992),
.B(n_959),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_990),
.B(n_868),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_990),
.B(n_857),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_942),
.B1(n_932),
.B2(n_897),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_997),
.A2(n_897),
.B(n_924),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_998),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_1003),
.B(n_860),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_998),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1000),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_1002),
.B(n_928),
.C(n_925),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_1007),
.B(n_893),
.C(n_876),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_1005),
.A2(n_1004),
.B1(n_999),
.B2(n_1006),
.C(n_944),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1010),
.Y(n_1018)
);

AOI211xp5_ASAP7_75t_SL g1019 ( 
.A1(n_1012),
.A2(n_1008),
.B(n_1009),
.C(n_1015),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_1011),
.Y(n_1020)
);

OAI322xp33_ASAP7_75t_L g1021 ( 
.A1(n_1014),
.A2(n_928),
.A3(n_924),
.B1(n_999),
.B2(n_944),
.C1(n_962),
.C2(n_954),
.Y(n_1021)
);

OAI321xp33_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_925),
.A3(n_906),
.B1(n_916),
.B2(n_877),
.C(n_887),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1013),
.B(n_945),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_1013),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1013),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1020),
.B(n_857),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_L g1027 ( 
.A(n_1017),
.B(n_857),
.C(n_896),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_SL g1028 ( 
.A1(n_1025),
.A2(n_906),
.B1(n_916),
.B2(n_877),
.C(n_947),
.Y(n_1028)
);

AOI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1024),
.A2(n_899),
.B(n_896),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_1018),
.A2(n_899),
.B(n_896),
.Y(n_1030)
);

AOI322xp5_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_900),
.A3(n_913),
.B1(n_952),
.B2(n_954),
.C1(n_958),
.C2(n_968),
.Y(n_1031)
);

INVxp67_ASAP7_75t_SL g1032 ( 
.A(n_1019),
.Y(n_1032)
);

OAI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1021),
.A2(n_904),
.B1(n_906),
.B2(n_958),
.C(n_960),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_1021),
.A2(n_926),
.B1(n_968),
.B2(n_960),
.C(n_905),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_1032),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1026),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1027),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1033),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1034),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1029),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1030),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1031),
.Y(n_1043)
);

CKINVDCx6p67_ASAP7_75t_R g1044 ( 
.A(n_1026),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1044),
.B(n_1022),
.Y(n_1045)
);

NOR3x1_ASAP7_75t_L g1046 ( 
.A(n_1043),
.B(n_911),
.C(n_898),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1035),
.B(n_939),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1035),
.B(n_946),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_1040),
.B(n_869),
.C(n_879),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1036),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1038),
.B(n_869),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1039),
.B(n_1037),
.C(n_1042),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_1052),
.B(n_1050),
.C(n_1049),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1045),
.A2(n_1041),
.B(n_926),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_1051),
.B(n_869),
.Y(n_1055)
);

XNOR2x1_ASAP7_75t_L g1056 ( 
.A(n_1047),
.B(n_153),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_1048),
.B(n_926),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_1046),
.A2(n_952),
.B(n_940),
.C(n_951),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_1050),
.B(n_900),
.C(n_913),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1053),
.B(n_879),
.C(n_869),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_1055),
.B(n_869),
.Y(n_1061)
);

AOI32xp33_ASAP7_75t_L g1062 ( 
.A1(n_1056),
.A2(n_917),
.A3(n_949),
.B1(n_940),
.B2(n_889),
.Y(n_1062)
);

AOI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_1054),
.A2(n_926),
.B1(n_879),
.B2(n_905),
.C(n_918),
.Y(n_1063)
);

OAI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_1059),
.A2(n_906),
.B1(n_904),
.B2(n_879),
.C(n_889),
.Y(n_1064)
);

NAND5xp2_ASAP7_75t_L g1065 ( 
.A(n_1058),
.B(n_949),
.C(n_922),
.D(n_901),
.E(n_927),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_1057),
.B(n_154),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1053),
.A2(n_879),
.B1(n_905),
.B2(n_922),
.C(n_901),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1056),
.B(n_921),
.Y(n_1068)
);

NAND5xp2_ASAP7_75t_L g1069 ( 
.A(n_1053),
.B(n_927),
.C(n_156),
.D(n_157),
.E(n_158),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1066),
.A2(n_906),
.B(n_921),
.Y(n_1070)
);

CKINVDCx12_ASAP7_75t_R g1071 ( 
.A(n_1069),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1060),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1061),
.B(n_865),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1065),
.B(n_904),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_1062),
.B(n_155),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_L g1077 ( 
.A(n_1064),
.B(n_927),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1067),
.B(n_921),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1074),
.A2(n_1063),
.B(n_921),
.Y(n_1079)
);

NAND4xp75_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_904),
.C(n_161),
.D(n_162),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1077),
.B(n_865),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1076),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1071),
.Y(n_1083)
);

XNOR2x1_ASAP7_75t_L g1084 ( 
.A(n_1075),
.B(n_160),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1073),
.B(n_927),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1078),
.Y(n_1086)
);

NOR3x1_ASAP7_75t_L g1087 ( 
.A(n_1070),
.B(n_164),
.C(n_167),
.Y(n_1087)
);

XOR2x1_ASAP7_75t_SL g1088 ( 
.A(n_1071),
.B(n_168),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1072),
.B(n_863),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1072),
.B(n_905),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_SL g1091 ( 
.A(n_1072),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1091),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1083),
.Y(n_1093)
);

NOR4xp25_ASAP7_75t_L g1094 ( 
.A(n_1082),
.B(n_169),
.C(n_171),
.D(n_172),
.Y(n_1094)
);

XNOR2xp5_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_174),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1087),
.Y(n_1096)
);

XNOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1088),
.B(n_176),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1089),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1086),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1081),
.B(n_864),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1093),
.Y(n_1101)
);

OR3x1_ASAP7_75t_L g1102 ( 
.A(n_1098),
.B(n_1079),
.C(n_1080),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1092),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1096),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_1097),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1099),
.A2(n_1085),
.B1(n_1090),
.B2(n_862),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1095),
.Y(n_1107)
);

XOR2xp5_ASAP7_75t_L g1108 ( 
.A(n_1103),
.B(n_1094),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1101),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1104),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_1110),
.A2(n_1107),
.B(n_1105),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1111),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1112),
.B(n_1109),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_1108),
.B(n_1106),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_1102),
.B1(n_1100),
.B2(n_862),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1114),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1113),
.A2(n_864),
.B1(n_863),
.B2(n_915),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_182),
.B(n_183),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_185),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1117),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_915),
.B1(n_912),
.B2(n_875),
.Y(n_1121)
);

AO221x2_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1122),
.A2(n_1118),
.B1(n_190),
.B2(n_192),
.Y(n_1123)
);

AOI211xp5_ASAP7_75t_L g1124 ( 
.A1(n_1123),
.A2(n_1121),
.B(n_193),
.C(n_196),
.Y(n_1124)
);


endmodule