module fake_jpeg_31926_n_424 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_424);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_424;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_62),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_56),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_14),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_19),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_26),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_42),
.B1(n_39),
.B2(n_34),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_121),
.B1(n_39),
.B2(n_31),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_58),
.B1(n_82),
.B2(n_80),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_65),
.B1(n_77),
.B2(n_76),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_21),
.B(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_99),
.B(n_26),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_48),
.A2(n_36),
.B1(n_38),
.B2(n_27),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_117),
.B(n_26),
.C(n_70),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_124),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_63),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_46),
.A2(n_26),
.B1(n_20),
.B2(n_35),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_55),
.B(n_26),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_45),
.B(n_42),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_123),
.B1(n_122),
.B2(n_112),
.Y(n_170)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_143),
.B1(n_152),
.B2(n_153),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_150),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_36),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_28),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_28),
.B1(n_24),
.B2(n_25),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_66),
.B1(n_75),
.B2(n_74),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_44),
.B1(n_67),
.B2(n_72),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_98),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_25),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_105),
.B1(n_51),
.B2(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_160),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.Y(n_177)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_118),
.B1(n_93),
.B2(n_52),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_25),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_122),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_172),
.B1(n_180),
.B2(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_117),
.B1(n_103),
.B2(n_123),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_117),
.B1(n_90),
.B2(n_116),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_35),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_142),
.C(n_40),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_202),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_134),
.A3(n_151),
.B1(n_136),
.B2(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_151),
.B1(n_90),
.B2(n_81),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_208),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_113),
.B1(n_116),
.B2(n_59),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_139),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_148),
.B(n_128),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_176),
.B(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_147),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_164),
.B(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_183),
.B1(n_165),
.B2(n_168),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_218),
.B1(n_228),
.B2(n_235),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_165),
.B1(n_170),
.B2(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_186),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_208),
.C(n_211),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_188),
.B(n_205),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_185),
.B1(n_167),
.B2(n_176),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_179),
.B(n_167),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_225),
.B(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_192),
.B1(n_206),
.B2(n_197),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_197),
.B1(n_198),
.B2(n_212),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_220),
.B1(n_234),
.B2(n_230),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_238),
.B(n_227),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_195),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_239),
.A2(n_245),
.B(n_254),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_198),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_246),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_208),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_252),
.C(n_262),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_248),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_215),
.B(n_192),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_244),
.B(n_233),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_198),
.B1(n_209),
.B2(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_259),
.Y(n_263)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_256),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_188),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_226),
.C(n_232),
.Y(n_252)
);

OAI221xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_202),
.B1(n_199),
.B2(n_196),
.C(n_40),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_203),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_182),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_181),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_237),
.B1(n_239),
.B2(n_254),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_228),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_268),
.Y(n_308)
);

AOI22x1_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_218),
.B1(n_235),
.B2(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_216),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_272),
.B(n_154),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_217),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_218),
.C(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_283),
.C(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_281),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_227),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_290),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_233),
.C(n_227),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_236),
.C(n_245),
.Y(n_287)
);

AO22x1_ASAP7_75t_L g288 ( 
.A1(n_248),
.A2(n_227),
.B1(n_146),
.B2(n_207),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_288),
.A2(n_119),
.B(n_107),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_240),
.C(n_236),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_207),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_169),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_304),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_274),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_295),
.A2(n_296),
.B1(n_302),
.B2(n_309),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_260),
.B1(n_246),
.B2(n_258),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_263),
.A2(n_249),
.B1(n_253),
.B2(n_250),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_299),
.B1(n_277),
.B2(n_284),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_250),
.B1(n_181),
.B2(n_205),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_169),
.B(n_145),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_301),
.A2(n_312),
.B(n_316),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_189),
.B1(n_175),
.B2(n_169),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_153),
.C(n_171),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_289),
.C(n_272),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_189),
.B1(n_131),
.B2(n_20),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_307),
.A2(n_286),
.B1(n_265),
.B2(n_280),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_311),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_171),
.B1(n_107),
.B2(n_158),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_269),
.B(n_138),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_94),
.B(n_119),
.Y(n_312)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_145),
.B(n_115),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_278),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_338),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_319),
.A2(n_334),
.B1(n_340),
.B2(n_271),
.Y(n_350)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_300),
.B1(n_297),
.B2(n_294),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_331),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_281),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_326),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_328),
.C(n_335),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_283),
.C(n_285),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_302),
.B1(n_131),
.B2(n_138),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_298),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_279),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_14),
.B(n_13),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_266),
.C(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_336),
.A2(n_270),
.B1(n_299),
.B2(n_316),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_305),
.B(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_145),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_275),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_282),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_340),
.C(n_315),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_266),
.C(n_290),
.Y(n_340)
);

AO221x1_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_297),
.B1(n_280),
.B2(n_270),
.C(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_314),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_339),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_294),
.B1(n_271),
.B2(n_314),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_357),
.B1(n_320),
.B2(n_157),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_320),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_350),
.A2(n_352),
.B1(n_353),
.B2(n_338),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_319),
.A2(n_161),
.B1(n_159),
.B2(n_135),
.Y(n_353)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_152),
.B1(n_149),
.B2(n_129),
.Y(n_355)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_356),
.B(n_346),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_113),
.B1(n_20),
.B2(n_69),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_358),
.B(n_322),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_364),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_318),
.C(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_347),
.C(n_345),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_346),
.B(n_327),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_372),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_371),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_325),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_14),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_360),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_359),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_376),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_156),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_385),
.C(n_371),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_363),
.A2(n_345),
.B(n_351),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_378),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_350),
.C(n_348),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_380),
.B(n_383),
.Y(n_390)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_351),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_344),
.C(n_353),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_386),
.B(n_31),
.Y(n_396)
);

AOI31xp67_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_360),
.A3(n_365),
.B(n_344),
.Y(n_389)
);

AOI322xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_95),
.A3(n_73),
.B1(n_64),
.B2(n_120),
.C1(n_109),
.C2(n_5),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_369),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_393),
.C(n_0),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_376),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_395),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_384),
.A2(n_375),
.B1(n_366),
.B2(n_101),
.Y(n_395)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_377),
.B(n_387),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_397),
.A2(n_398),
.B(n_388),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_95),
.B(n_50),
.Y(n_398)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_400),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_390),
.A2(n_384),
.B(n_120),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_401),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_403),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_399),
.A2(n_109),
.B1(n_1),
.B2(n_2),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_22),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_406),
.C(n_3),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_394),
.A2(n_0),
.B(n_2),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_405),
.A2(n_3),
.B(n_5),
.Y(n_409)
);

AOI322xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_413),
.A3(n_408),
.B1(n_404),
.B2(n_393),
.C1(n_7),
.C2(n_8),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_407),
.A2(n_391),
.B(n_398),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_7),
.C(n_9),
.Y(n_418)
);

AOI21x1_ASAP7_75t_L g420 ( 
.A1(n_415),
.A2(n_416),
.B(n_417),
.Y(n_420)
);

AOI322xp5_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_416)
);

AOI322xp5_ASAP7_75t_L g417 ( 
.A1(n_412),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_411),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_419),
.A2(n_9),
.B(n_10),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_420),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_10),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_423),
.A2(n_10),
.B1(n_11),
.B2(n_346),
.Y(n_424)
);


endmodule