module fake_jpeg_4312_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_51)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_18),
.B1(n_16),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_46),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_14),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_44),
.C(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_42),
.C(n_41),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_8),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_20),
.B1(n_14),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_63),
.B1(n_27),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_61),
.B1(n_25),
.B2(n_27),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_22),
.B1(n_28),
.B2(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_67),
.Y(n_96)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_78),
.Y(n_120)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_50),
.B1(n_48),
.B2(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_98),
.B1(n_56),
.B2(n_49),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_35),
.B(n_41),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_73),
.B(n_52),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_47),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_56),
.B1(n_10),
.B2(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_5),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_60),
.B1(n_73),
.B2(n_72),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_113),
.B(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_62),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_115),
.B1(n_98),
.B2(n_82),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_71),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_12),
.C(n_11),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_75),
.B1(n_54),
.B2(n_53),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_96),
.C(n_90),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_133),
.B1(n_136),
.B2(n_120),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_102),
.C(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_96),
.C(n_77),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_79),
.B1(n_115),
.B2(n_111),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_94),
.B(n_82),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_141),
.B(n_143),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_101),
.B(n_120),
.C(n_119),
.D(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_108),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_123),
.C(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_118),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_146),
.B(n_148),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_117),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_121),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_106),
.A3(n_104),
.B1(n_92),
.B2(n_88),
.C1(n_80),
.C2(n_105),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_121),
.C(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_122),
.B1(n_130),
.B2(n_80),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_157),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_152),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_156),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_154),
.B(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_149),
.C(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_155),
.C(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_137),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_167),
.C1(n_165),
.C2(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);


endmodule