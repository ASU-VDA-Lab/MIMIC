module fake_jpeg_26263_n_222 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_33),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_62),
.B1(n_30),
.B2(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_24),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_35),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_75),
.B(n_80),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_95),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_45),
.B1(n_38),
.B2(n_43),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_63),
.B1(n_26),
.B2(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_90),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_57),
.B1(n_25),
.B2(n_26),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_18),
.B1(n_17),
.B2(n_26),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_57),
.B1(n_44),
.B2(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_75),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_36),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_18),
.C(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_35),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_10),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_103),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_114),
.B1(n_89),
.B2(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_122),
.C(n_73),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_29),
.CI(n_18),
.CON(n_112),
.SN(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_71),
.B(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_73),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_80),
.C(n_79),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_130),
.B(n_113),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_72),
.B(n_89),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_131),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_129),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_83),
.C(n_81),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_110),
.C(n_104),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_81),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_9),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_146),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_87),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_133),
.B(n_107),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_149),
.B(n_153),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_117),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_136),
.B(n_139),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_111),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_132),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_112),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_137),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_131),
.B1(n_130),
.B2(n_108),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_142),
.B1(n_126),
.B2(n_105),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_169),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_155),
.A3(n_160),
.B1(n_149),
.B2(n_153),
.C(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_159),
.C(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_165),
.Y(n_188)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_156),
.B1(n_141),
.B2(n_105),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_135),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_179),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_105),
.A3(n_135),
.B1(n_112),
.B2(n_128),
.C1(n_145),
.C2(n_115),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_192),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_148),
.C(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_171),
.B1(n_168),
.B2(n_13),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_101),
.C(n_163),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_116),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_180),
.B(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_182),
.B(n_184),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_197),
.B(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_183),
.B1(n_188),
.B2(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_189),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_212),
.B(n_213),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_193),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_189),
.A3(n_8),
.B(n_13),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_7),
.C(n_14),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_202),
.C(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_16),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_208),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_215),
.C(n_203),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_204),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);


endmodule