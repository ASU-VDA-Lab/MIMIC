module fake_jpeg_29320_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_23),
.B1(n_4),
.B2(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_22),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_17),
.B1(n_19),
.B2(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_10),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_28),
.B1(n_22),
.B2(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_47),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_12),
.A3(n_15),
.B1(n_20),
.B2(n_21),
.C1(n_25),
.C2(n_24),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_21),
.A3(n_25),
.B1(n_15),
.B2(n_33),
.C1(n_44),
.C2(n_16),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_38),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_16),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_48),
.C(n_6),
.Y(n_51)
);


endmodule