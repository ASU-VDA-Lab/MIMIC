module real_aes_7862_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_241;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_1), .A2(n_159), .B(n_162), .C(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_2), .A2(n_188), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g488 ( .A(n_3), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_4), .B(n_218), .Y(n_217) );
AOI21xp33_ASAP7_75t_L g471 ( .A1(n_5), .A2(n_188), .B(n_472), .Y(n_471) );
AND2x6_ASAP7_75t_L g159 ( .A(n_6), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g255 ( .A(n_7), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_41), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_8), .B(n_41), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_9), .A2(n_187), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_10), .B(n_171), .Y(n_244) );
INVx1_ASAP7_75t_L g476 ( .A(n_11), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_12), .B(n_212), .Y(n_511) );
INVx1_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
INVx1_ASAP7_75t_L g523 ( .A(n_14), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_15), .A2(n_78), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_15), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_16), .A2(n_196), .B(n_277), .C(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_17), .B(n_218), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_18), .B(n_454), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_19), .B(n_188), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_20), .B(n_202), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_21), .A2(n_212), .B(n_263), .C(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_22), .B(n_218), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_23), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_24), .A2(n_198), .B(n_279), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_25), .B(n_171), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_26), .Y(n_153) );
INVx1_ASAP7_75t_L g225 ( .A(n_27), .Y(n_225) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_28), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_29), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_30), .B(n_171), .Y(n_489) );
INVx1_ASAP7_75t_L g194 ( .A(n_31), .Y(n_194) );
INVx1_ASAP7_75t_L g466 ( .A(n_32), .Y(n_466) );
INVx2_ASAP7_75t_L g157 ( .A(n_33), .Y(n_157) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_34), .A2(n_130), .B1(n_133), .B2(n_726), .C1(n_727), .C2(n_729), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_35), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_36), .A2(n_212), .B(n_213), .C(n_215), .Y(n_211) );
INVxp67_ASAP7_75t_L g197 ( .A(n_37), .Y(n_197) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_38), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_39), .A2(n_162), .B(n_224), .C(n_228), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_40), .A2(n_159), .B(n_162), .C(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g465 ( .A(n_42), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_43), .A2(n_173), .B(n_253), .C(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_44), .B(n_171), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_45), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_46), .Y(n_190) );
INVx1_ASAP7_75t_L g261 ( .A(n_47), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_48), .Y(n_467) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_49), .A2(n_59), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_49), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_50), .B(n_188), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_51), .A2(n_162), .B1(n_265), .B2(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_52), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g485 ( .A(n_53), .Y(n_485) );
CKINVDCx14_ASAP7_75t_R g251 ( .A(n_54), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_55), .A2(n_215), .B(n_253), .C(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_56), .Y(n_128) );
INVx1_ASAP7_75t_L g473 ( .A(n_57), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_58), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_59), .Y(n_739) );
INVx1_ASAP7_75t_L g160 ( .A(n_60), .Y(n_160) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
INVx1_ASAP7_75t_SL g214 ( .A(n_62), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_64), .B(n_218), .Y(n_267) );
INVx1_ASAP7_75t_L g166 ( .A(n_65), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_SL g453 ( .A1(n_66), .A2(n_215), .B(n_454), .C(n_455), .Y(n_453) );
INVxp67_ASAP7_75t_L g456 ( .A(n_67), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_68), .A2(n_102), .B1(n_115), .B2(n_742), .Y(n_101) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_70), .A2(n_188), .B(n_250), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_71), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_72), .A2(n_188), .B(n_274), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_73), .Y(n_469) );
INVx1_ASAP7_75t_L g529 ( .A(n_74), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_75), .A2(n_187), .B(n_189), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g222 ( .A(n_76), .Y(n_222) );
INVx1_ASAP7_75t_L g275 ( .A(n_77), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_78), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_79), .A2(n_159), .B(n_162), .C(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_80), .A2(n_188), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g278 ( .A(n_81), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_82), .B(n_195), .Y(n_500) );
INVx2_ASAP7_75t_L g148 ( .A(n_83), .Y(n_148) );
INVx1_ASAP7_75t_L g243 ( .A(n_84), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_85), .B(n_454), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_86), .A2(n_159), .B(n_162), .C(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
OR2x2_ASAP7_75t_L g124 ( .A(n_87), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g441 ( .A(n_87), .B(n_126), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_88), .A2(n_162), .B(n_165), .C(n_175), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_89), .B(n_180), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_90), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_91), .A2(n_159), .B(n_162), .C(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_92), .Y(n_515) );
INVx1_ASAP7_75t_L g452 ( .A(n_93), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_94), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_95), .B(n_195), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_96), .B(n_146), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_97), .B(n_146), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g264 ( .A(n_99), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_100), .A2(n_188), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g743 ( .A(n_105), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g126 ( .A(n_110), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g725 ( .A(n_111), .B(n_126), .Y(n_725) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_111), .B(n_125), .Y(n_731) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_129), .B1(n_732), .B2(n_734), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g733 ( .A(n_119), .Y(n_733) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_121), .A2(n_735), .B(n_740), .Y(n_734) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_128), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g741 ( .A(n_124), .Y(n_741) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g726 ( .A(n_130), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_441), .B1(n_442), .B2(n_723), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_134), .A2(n_135), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_135), .A2(n_441), .B1(n_723), .B2(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_375), .Y(n_135) );
NAND5xp2_ASAP7_75t_L g136 ( .A(n_137), .B(n_304), .C(n_334), .D(n_355), .E(n_361), .Y(n_136) );
AOI221xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_234), .B1(n_268), .B2(n_270), .C(n_281), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_231), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_203), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_SL g355 ( .A1(n_142), .A2(n_219), .B(n_356), .C(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g425 ( .A(n_142), .B(n_220), .Y(n_425) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_181), .Y(n_142) );
AND2x2_ASAP7_75t_L g283 ( .A(n_143), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g287 ( .A(n_143), .B(n_284), .Y(n_287) );
OR2x2_ASAP7_75t_L g313 ( .A(n_143), .B(n_220), .Y(n_313) );
AND2x2_ASAP7_75t_L g315 ( .A(n_143), .B(n_206), .Y(n_315) );
AND2x2_ASAP7_75t_L g333 ( .A(n_143), .B(n_205), .Y(n_333) );
INVx1_ASAP7_75t_L g366 ( .A(n_143), .Y(n_366) );
INVx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
BUFx2_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
AND2x2_ASAP7_75t_L g269 ( .A(n_144), .B(n_206), .Y(n_269) );
AND2x2_ASAP7_75t_L g422 ( .A(n_144), .B(n_220), .Y(n_422) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_152), .B(n_177), .Y(n_144) );
INVx3_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_145), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_145), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_SL g502 ( .A(n_145), .B(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_146), .A2(n_450), .B(n_457), .Y(n_449) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_148), .B(n_149), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_161), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_154), .A2(n_180), .B(n_222), .C(n_223), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_154), .A2(n_240), .B(n_241), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_154), .A2(n_176), .B1(n_463), .B2(n_467), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_154), .A2(n_485), .B(n_486), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_154), .A2(n_529), .B(n_530), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
AND2x4_ASAP7_75t_L g188 ( .A(n_155), .B(n_159), .Y(n_188) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g199 ( .A(n_156), .Y(n_199) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
INVx1_ASAP7_75t_L g266 ( .A(n_157), .Y(n_266) );
INVx1_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_158), .Y(n_169) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
INVx3_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx1_ASAP7_75t_L g454 ( .A(n_158), .Y(n_454) );
INVx4_ASAP7_75t_SL g176 ( .A(n_159), .Y(n_176) );
BUFx3_ASAP7_75t_L g228 ( .A(n_159), .Y(n_228) );
INVx5_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
AND2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx3_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_170), .C(n_172), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_172), .B(n_243), .C(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_168), .A2(n_169), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
INVx4_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
INVx2_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_172), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_172), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g279 ( .A(n_174), .Y(n_279) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_176), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_191), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_176), .A2(n_191), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_176), .A2(n_191), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_SL g274 ( .A1(n_176), .A2(n_191), .B(n_275), .C(n_276), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_176), .A2(n_191), .B(n_452), .C(n_453), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_176), .A2(n_191), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_176), .A2(n_191), .B(n_520), .C(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_179), .A2(n_507), .B(n_514), .Y(n_506) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g238 ( .A(n_180), .Y(n_238) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_180), .A2(n_249), .B(n_256), .Y(n_248) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_180), .A2(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g303 ( .A(n_181), .B(n_204), .Y(n_303) );
OR2x2_ASAP7_75t_L g307 ( .A(n_181), .B(n_220), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_181), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g379 ( .A(n_181), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_181), .B(n_341), .Y(n_427) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_185), .B(n_200), .Y(n_181) );
INVx1_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_182), .A2(n_528), .B(n_534), .Y(n_527) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_SL g496 ( .A1(n_183), .A2(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_184), .A2(n_462), .B(n_468), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_184), .B(n_469), .Y(n_468) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_184), .A2(n_484), .B(n_491), .Y(n_483) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_186), .A2(n_201), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_193), .B(n_199), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B1(n_197), .B2(n_198), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_195), .A2(n_225), .B(n_226), .C(n_227), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_195), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
INVx5_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_196), .B(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_196), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_196), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_198), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_198), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_198), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OAI322xp33_ASAP7_75t_L g428 ( .A1(n_203), .A2(n_364), .A3(n_387), .B1(n_408), .B2(n_429), .C1(n_431), .C2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_204), .B(n_284), .Y(n_431) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_219), .Y(n_204) );
AND2x2_ASAP7_75t_L g232 ( .A(n_205), .B(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g300 ( .A(n_205), .B(n_220), .Y(n_300) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g341 ( .A(n_206), .B(n_220), .Y(n_341) );
AND2x2_ASAP7_75t_L g385 ( .A(n_206), .B(n_219), .Y(n_385) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_217), .Y(n_206) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_207), .A2(n_259), .B(n_267), .Y(n_258) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_207), .A2(n_273), .B(n_280), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_212), .B(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_216), .Y(n_512) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_218), .A2(n_471), .B(n_477), .Y(n_470) );
AND2x2_ASAP7_75t_L g268 ( .A(n_219), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g286 ( .A(n_219), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_219), .B(n_315), .Y(n_439) );
INVx3_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g231 ( .A(n_220), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_220), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g353 ( .A(n_220), .B(n_284), .Y(n_353) );
AND2x2_ASAP7_75t_L g380 ( .A(n_220), .B(n_315), .Y(n_380) );
OR2x2_ASAP7_75t_L g436 ( .A(n_220), .B(n_287), .Y(n_436) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_229), .Y(n_220) );
INVx1_ASAP7_75t_SL g322 ( .A(n_231), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_232), .B(n_353), .Y(n_354) );
AND2x2_ASAP7_75t_L g388 ( .A(n_232), .B(n_378), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_232), .B(n_311), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_232), .B(n_433), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_234), .A2(n_268), .A3(n_407), .B(n_409), .Y(n_406) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_235), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g389 ( .A(n_235), .B(n_324), .Y(n_389) );
OR2x2_ASAP7_75t_L g396 ( .A(n_235), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g408 ( .A(n_235), .B(n_297), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g342 ( .A(n_236), .B(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g270 ( .A(n_237), .B(n_271), .Y(n_270) );
INVx4_ASAP7_75t_L g291 ( .A(n_237), .Y(n_291) );
AND2x2_ASAP7_75t_L g328 ( .A(n_237), .B(n_272), .Y(n_328) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_245), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_238), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_238), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_238), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g327 ( .A(n_247), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g397 ( .A(n_247), .Y(n_397) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_257), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_248), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g297 ( .A(n_248), .B(n_258), .Y(n_297) );
INVx2_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_248), .B(n_258), .Y(n_331) );
AND2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_294), .Y(n_338) );
BUFx3_ASAP7_75t_L g348 ( .A(n_248), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_248), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_257), .B(n_291), .Y(n_301) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g271 ( .A(n_258), .B(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_258), .Y(n_325) );
INVx2_ASAP7_75t_L g490 ( .A(n_265), .Y(n_490) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g308 ( .A(n_269), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_269), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_269), .B(n_378), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_270), .B(n_348), .Y(n_401) );
INVx1_ASAP7_75t_SL g435 ( .A(n_270), .Y(n_435) );
INVx1_ASAP7_75t_SL g343 ( .A(n_271), .Y(n_343) );
INVx1_ASAP7_75t_SL g294 ( .A(n_272), .Y(n_294) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_272), .Y(n_305) );
OR2x2_ASAP7_75t_L g316 ( .A(n_272), .B(n_291), .Y(n_316) );
AND2x2_ASAP7_75t_L g330 ( .A(n_272), .B(n_291), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_272), .B(n_320), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_286), .B(n_288), .C(n_299), .Y(n_281) );
AOI31xp33_ASAP7_75t_L g398 ( .A1(n_282), .A2(n_399), .A3(n_400), .B(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g371 ( .A(n_283), .B(n_300), .Y(n_371) );
BUFx3_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_284), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g347 ( .A(n_284), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_284), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g302 ( .A(n_287), .Y(n_302) );
OAI222xp33_ASAP7_75t_L g411 ( .A1(n_287), .A2(n_412), .B1(n_415), .B2(n_416), .C1(n_417), .C2(n_418), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_295), .Y(n_288) );
INVx1_ASAP7_75t_L g417 ( .A(n_289), .Y(n_417) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_291), .B(n_294), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_291), .B(n_317), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_291), .B(n_292), .Y(n_387) );
INVx1_ASAP7_75t_L g438 ( .A(n_291), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_292), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g440 ( .A(n_292), .Y(n_440) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g320 ( .A(n_293), .Y(n_320) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g299 ( .A1(n_295), .A2(n_300), .A3(n_301), .B1(n_302), .B2(n_303), .Y(n_299) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_297), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g374 ( .A(n_297), .Y(n_374) );
OR2x2_ASAP7_75t_L g415 ( .A(n_297), .B(n_316), .Y(n_415) );
INVx1_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_300), .B(n_311), .Y(n_336) );
INVx3_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
AOI322xp5_ASAP7_75t_L g361 ( .A1(n_300), .A2(n_345), .A3(n_362), .B1(n_364), .B2(n_367), .C1(n_371), .C2(n_372), .Y(n_361) );
AND2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_L g414 ( .A(n_301), .Y(n_414) );
A2O1A1O1Ixp25_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B(n_309), .C(n_317), .D(n_318), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_305), .B(n_348), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_307), .A2(n_319), .B1(n_322), .B2(n_323), .C(n_326), .Y(n_318) );
INVx1_ASAP7_75t_SL g433 ( .A(n_307), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B(n_316), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_311), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_313), .A2(n_397), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_403) );
OAI222xp33_ASAP7_75t_L g434 ( .A1(n_314), .A2(n_435), .B1(n_436), .B2(n_437), .C1(n_439), .C2(n_440), .Y(n_434) );
AND2x2_ASAP7_75t_L g392 ( .A(n_315), .B(n_378), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_315), .A2(n_330), .B(n_377), .Y(n_404) );
INVx1_ASAP7_75t_L g418 ( .A(n_315), .Y(n_418) );
INVx2_ASAP7_75t_SL g321 ( .A(n_316), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_317), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_SL g358 ( .A(n_320), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_320), .B(n_330), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_321), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_321), .B(n_331), .Y(n_360) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI21xp5_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B(n_332), .Y(n_326) );
INVx1_ASAP7_75t_SL g344 ( .A(n_328), .Y(n_344) );
AND2x2_ASAP7_75t_L g391 ( .A(n_328), .B(n_374), .Y(n_391) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g430 ( .A(n_330), .B(n_348), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_331), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g416 ( .A(n_332), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_339), .B2(n_346), .C(n_349), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_344), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_343), .A2(n_350), .B1(n_352), .B2(n_354), .Y(n_349) );
OR2x2_ASAP7_75t_L g420 ( .A(n_344), .B(n_348), .Y(n_420) );
OR2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_358), .Y(n_423) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_365), .A2(n_420), .B1(n_421), .B2(n_423), .C(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND3xp33_ASAP7_75t_SL g375 ( .A(n_376), .B(n_390), .C(n_402), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_383), .B2(n_386), .C1(n_388), .C2(n_389), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_378), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g405 ( .A(n_391), .Y(n_405) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g424 ( .A1(n_395), .A2(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
NOR5xp2_ASAP7_75t_L g402 ( .A(n_403), .B(n_411), .C(n_419), .D(n_428), .E(n_434), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g728 ( .A(n_442), .Y(n_728) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_443), .B(n_660), .Y(n_442) );
NOR4xp25_ASAP7_75t_L g443 ( .A(n_444), .B(n_590), .C(n_621), .D(n_640), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_548), .C(n_563), .D(n_581), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_493), .B1(n_525), .B2(n_536), .C1(n_541), .C2(n_543), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_478), .Y(n_446) );
INVx1_ASAP7_75t_L g604 ( .A(n_447), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_458), .Y(n_447) );
AND2x2_ASAP7_75t_L g479 ( .A(n_448), .B(n_470), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_448), .B(n_482), .Y(n_633) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g540 ( .A(n_449), .B(n_460), .Y(n_540) );
AND2x2_ASAP7_75t_L g549 ( .A(n_449), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g575 ( .A(n_449), .Y(n_575) );
AND2x2_ASAP7_75t_L g596 ( .A(n_449), .B(n_460), .Y(n_596) );
BUFx2_ASAP7_75t_L g619 ( .A(n_449), .Y(n_619) );
AND2x2_ASAP7_75t_L g643 ( .A(n_449), .B(n_461), .Y(n_643) );
AND2x2_ASAP7_75t_L g707 ( .A(n_449), .B(n_470), .Y(n_707) );
AND2x2_ASAP7_75t_L g608 ( .A(n_458), .B(n_539), .Y(n_608) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_459), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .Y(n_459) );
OR2x2_ASAP7_75t_L g568 ( .A(n_460), .B(n_483), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_460), .B(n_539), .Y(n_580) );
BUFx2_ASAP7_75t_L g712 ( .A(n_460), .Y(n_712) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g481 ( .A(n_461), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g562 ( .A(n_461), .B(n_483), .Y(n_562) );
AND2x2_ASAP7_75t_L g615 ( .A(n_461), .B(n_470), .Y(n_615) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_461), .Y(n_651) );
AND2x2_ASAP7_75t_L g538 ( .A(n_470), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_SL g550 ( .A(n_470), .Y(n_550) );
INVx2_ASAP7_75t_L g561 ( .A(n_470), .Y(n_561) );
BUFx2_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_470), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AOI332xp33_ASAP7_75t_L g563 ( .A1(n_479), .A2(n_564), .A3(n_568), .B1(n_569), .B2(n_573), .B3(n_576), .C1(n_577), .C2(n_579), .Y(n_563) );
NAND2x1_ASAP7_75t_L g648 ( .A(n_479), .B(n_539), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_479), .B(n_553), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_SL g581 ( .A1(n_480), .A2(n_582), .B(n_585), .C(n_586), .Y(n_581) );
AND2x2_ASAP7_75t_L g720 ( .A(n_480), .B(n_561), .Y(n_720) );
INVx3_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g617 ( .A(n_481), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g622 ( .A(n_481), .B(n_619), .Y(n_622) );
INVx1_ASAP7_75t_L g553 ( .A(n_482), .Y(n_553) );
AND2x2_ASAP7_75t_L g656 ( .A(n_482), .B(n_615), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_482), .B(n_596), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_482), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_482), .B(n_574), .Y(n_682) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
OAI31xp33_ASAP7_75t_L g721 ( .A1(n_493), .A2(n_642), .A3(n_649), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
AND2x2_ASAP7_75t_L g525 ( .A(n_494), .B(n_526), .Y(n_525) );
NAND2x1_ASAP7_75t_SL g544 ( .A(n_494), .B(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_494), .Y(n_631) );
AND2x2_ASAP7_75t_L g636 ( .A(n_494), .B(n_547), .Y(n_636) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_495), .A2(n_549), .B(n_551), .C(n_554), .Y(n_548) );
OR2x2_ASAP7_75t_L g565 ( .A(n_495), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g578 ( .A(n_495), .Y(n_578) );
AND2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_527), .Y(n_584) );
INVx2_ASAP7_75t_L g602 ( .A(n_495), .Y(n_602) );
AND2x2_ASAP7_75t_L g613 ( .A(n_495), .B(n_567), .Y(n_613) );
AND2x2_ASAP7_75t_L g645 ( .A(n_495), .B(n_603), .Y(n_645) );
AND2x2_ASAP7_75t_L g649 ( .A(n_495), .B(n_572), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_495), .B(n_504), .Y(n_654) );
AND2x2_ASAP7_75t_L g688 ( .A(n_495), .B(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_495), .B(n_591), .Y(n_722) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g630 ( .A(n_504), .Y(n_630) );
AND2x2_ASAP7_75t_L g692 ( .A(n_504), .B(n_613), .Y(n_692) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
OR2x2_ASAP7_75t_L g546 ( .A(n_505), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g556 ( .A(n_505), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_505), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g664 ( .A(n_505), .Y(n_664) );
AND2x2_ASAP7_75t_L g681 ( .A(n_505), .B(n_527), .Y(n_681) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g572 ( .A(n_506), .B(n_516), .Y(n_572) );
AND2x2_ASAP7_75t_L g601 ( .A(n_506), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g612 ( .A(n_506), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_506), .B(n_567), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g526 ( .A(n_517), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g547 ( .A(n_517), .Y(n_547) );
AND2x2_ASAP7_75t_L g603 ( .A(n_517), .B(n_567), .Y(n_603) );
INVx1_ASAP7_75t_L g705 ( .A(n_525), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_526), .Y(n_709) );
INVx2_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_538), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_538), .B(n_643), .Y(n_701) );
OR2x2_ASAP7_75t_L g542 ( .A(n_539), .B(n_540), .Y(n_542) );
INVx1_ASAP7_75t_SL g594 ( .A(n_539), .Y(n_594) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_545), .A2(n_598), .B1(n_600), .B2(n_604), .C(n_605), .Y(n_597) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g625 ( .A(n_546), .B(n_589), .Y(n_625) );
INVx2_ASAP7_75t_L g557 ( .A(n_547), .Y(n_557) );
INVx1_ASAP7_75t_L g583 ( .A(n_547), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_547), .B(n_567), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_547), .B(n_570), .Y(n_677) );
INVx1_ASAP7_75t_L g685 ( .A(n_547), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_549), .B(n_553), .Y(n_599) );
AND2x4_ASAP7_75t_L g574 ( .A(n_550), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g687 ( .A(n_553), .B(n_643), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_556), .B(n_588), .Y(n_587) );
INVxp67_ASAP7_75t_L g695 ( .A(n_557), .Y(n_695) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g595 ( .A(n_561), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g667 ( .A(n_561), .B(n_643), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_561), .B(n_580), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g627 ( .A1(n_562), .A2(n_596), .A3(n_603), .B1(n_628), .B2(n_631), .C1(n_632), .C2(n_634), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_562), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g693 ( .A(n_565), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
INVx2_ASAP7_75t_L g570 ( .A(n_567), .Y(n_570) );
INVx1_ASAP7_75t_L g629 ( .A(n_567), .Y(n_629) );
CKINVDCx16_ASAP7_75t_R g576 ( .A(n_568), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_L g665 ( .A(n_570), .B(n_578), .Y(n_665) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g577 ( .A(n_572), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g620 ( .A(n_572), .B(n_613), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_572), .B(n_584), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g634 ( .A1(n_573), .A2(n_635), .B(n_637), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_573), .A2(n_705), .B1(n_706), .B2(n_708), .Y(n_704) );
INVx3_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_574), .B(n_594), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_576), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g716 ( .A(n_583), .Y(n_716) );
INVx4_ASAP7_75t_L g589 ( .A(n_584), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_584), .B(n_611), .Y(n_659) );
INVx1_ASAP7_75t_SL g671 ( .A(n_585), .Y(n_671) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_589), .B(n_685), .Y(n_684) );
OAI211xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B(n_597), .C(n_614), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g710 ( .A1(n_592), .A2(n_630), .B1(n_709), .B2(n_711), .C(n_713), .Y(n_710) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_594), .B(n_707), .Y(n_706) );
OAI31xp33_ASAP7_75t_L g686 ( .A1(n_595), .A2(n_672), .A3(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g626 ( .A(n_596), .Y(n_626) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g676 ( .A(n_601), .Y(n_676) );
AND2x2_ASAP7_75t_L g689 ( .A(n_603), .B(n_612), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_609), .Y(n_605) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_613), .B(n_716), .Y(n_715) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B1(n_625), .B2(n_626), .C(n_627), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_622), .A2(n_691), .B(n_693), .C(n_696), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_625), .B(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g652 ( .A(n_633), .Y(n_652) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g638 ( .A(n_636), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g680 ( .A(n_636), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B(n_646), .C(n_655), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_644), .A2(n_654), .B1(n_718), .B2(n_719), .C(n_721), .Y(n_717) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_650), .B2(n_653), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_657), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_SL g718 ( .A(n_657), .Y(n_718) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_690), .C(n_710), .D(n_717), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_666), .B(n_668), .C(n_686), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_674), .C(n_678), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g697 ( .A(n_675), .Y(n_697) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OR2x2_ASAP7_75t_L g708 ( .A(n_676), .B(n_709), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B(n_683), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_702), .C(n_704), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_707), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
endmodule