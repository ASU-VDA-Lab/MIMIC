module fake_jpeg_14058_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_49),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_50),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_54),
.Y(n_104)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_53),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_56),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_73),
.Y(n_101)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_72),
.Y(n_107)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_17),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_4),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_87),
.Y(n_119)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_85),
.Y(n_130)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_92),
.Y(n_139)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_5),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_22),
.B(n_14),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_21),
.B1(n_47),
.B2(n_44),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_103),
.A2(n_106),
.B1(n_112),
.B2(n_131),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_99),
.B1(n_95),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_45),
.B1(n_41),
.B2(n_29),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_126),
.Y(n_156)
);

CKINVDCx12_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_125),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_24),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_62),
.A2(n_41),
.B1(n_24),
.B2(n_35),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_23),
.B1(n_38),
.B2(n_36),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_145),
.B1(n_117),
.B2(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_50),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_49),
.B(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_143),
.B(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_63),
.B(n_23),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_105),
.A2(n_50),
.B(n_38),
.C(n_39),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_153),
.A2(n_164),
.B(n_166),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_6),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_161),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_171),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.C(n_131),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_104),
.B(n_140),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_181),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_183),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_190),
.Y(n_209)
);

OR2x2_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_106),
.B(n_117),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_185),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_187),
.B1(n_142),
.B2(n_189),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_135),
.B1(n_147),
.B2(n_100),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_116),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_100),
.B1(n_111),
.B2(n_134),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_204),
.B1(n_207),
.B2(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_103),
.B1(n_111),
.B2(n_114),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_162),
.B1(n_174),
.B2(n_182),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_116),
.B1(n_138),
.B2(n_121),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_154),
.A2(n_138),
.B1(n_121),
.B2(n_120),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_179),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_208),
.C(n_224),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_120),
.B1(n_142),
.B2(n_152),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_219),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_180),
.B(n_178),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_220),
.A2(n_164),
.B(n_173),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_153),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_175),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_156),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_228),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_157),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_232),
.Y(n_250)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_161),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_233),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_238),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_248),
.B(n_207),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_222),
.Y(n_241)
);

NOR2x1_ASAP7_75t_R g262 ( 
.A(n_241),
.B(n_247),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_170),
.B1(n_159),
.B2(n_163),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_245),
.B1(n_218),
.B2(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_193),
.B1(n_168),
.B2(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_212),
.B1(n_196),
.B2(n_223),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_177),
.C(n_192),
.Y(n_247)
);

AOI221xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_158),
.B1(n_220),
.B2(n_208),
.C(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_203),
.B1(n_198),
.B2(n_225),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_257),
.B1(n_239),
.B2(n_242),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_215),
.B1(n_209),
.B2(n_204),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_212),
.B(n_223),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_237),
.B(n_241),
.Y(n_272)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_235),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_268),
.B1(n_270),
.B2(n_260),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_237),
.B1(n_243),
.B2(n_234),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_279),
.B1(n_257),
.B2(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_255),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_231),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_233),
.C(n_247),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_262),
.C(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_245),
.A3(n_243),
.B1(n_232),
.B2(n_205),
.C1(n_221),
.C2(n_201),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_260),
.C(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.C(n_287),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_249),
.B1(n_269),
.B2(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_279),
.B1(n_276),
.B2(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_262),
.C(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_299),
.B1(n_277),
.B2(n_261),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_267),
.B(n_266),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_283),
.C(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_277),
.B1(n_265),
.B2(n_201),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_293),
.B(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_281),
.B1(n_290),
.B2(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_297),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_298),
.C(n_301),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_298),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_309),
.B1(n_295),
.B2(n_305),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_196),
.A3(n_205),
.B1(n_282),
.B2(n_296),
.C1(n_311),
.C2(n_315),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_318),
.Y(n_320)
);


endmodule