module real_aes_1926_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_793, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_793;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_0), .B(n_143), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_1), .A2(n_152), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_2), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_3), .B(n_143), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_4), .B(n_159), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_5), .B(n_159), .Y(n_222) );
INVx1_ASAP7_75t_L g150 ( .A(n_6), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_7), .B(n_159), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g788 ( .A(n_8), .Y(n_788) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_9), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g474 ( .A(n_10), .B(n_169), .Y(n_474) );
AND2x2_ASAP7_75t_L g534 ( .A(n_11), .B(n_138), .Y(n_534) );
INVx2_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
AOI221x1_ASAP7_75t_L g238 ( .A1(n_13), .A2(n_24), .B1(n_143), .B2(n_152), .C(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_14), .B(n_159), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_15), .B(n_787), .C(n_789), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_16), .B(n_143), .Y(n_142) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_17), .A2(n_138), .B(n_141), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_18), .B(n_177), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_19), .B(n_159), .Y(n_186) );
AO21x1_ASAP7_75t_L g217 ( .A1(n_20), .A2(n_143), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_21), .B(n_143), .Y(n_539) );
INVx1_ASAP7_75t_L g118 ( .A(n_22), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_23), .A2(n_89), .B1(n_143), .B2(n_479), .Y(n_478) );
NAND2x1_ASAP7_75t_L g208 ( .A(n_25), .B(n_159), .Y(n_208) );
NAND2x1_ASAP7_75t_L g196 ( .A(n_26), .B(n_161), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_27), .Y(n_766) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_28), .A2(n_86), .B(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g164 ( .A(n_28), .B(n_86), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_29), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_30), .B(n_161), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_31), .B(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_32), .A2(n_169), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_33), .B(n_161), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_34), .A2(n_152), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_35), .B(n_159), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_36), .A2(n_152), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g149 ( .A(n_37), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g153 ( .A(n_37), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g487 ( .A(n_37), .Y(n_487) );
OR2x6_ASAP7_75t_L g116 ( .A(n_38), .B(n_117), .Y(n_116) );
INVxp67_ASAP7_75t_L g789 ( .A(n_38), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_39), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_40), .B(n_143), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_41), .B(n_159), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_42), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_43), .B(n_161), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_44), .B(n_143), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_45), .A2(n_152), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_46), .A2(n_152), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_47), .B(n_161), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_48), .B(n_161), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_49), .B(n_143), .Y(n_505) );
INVx1_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_50), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_51), .B(n_159), .Y(n_472) );
AND2x2_ASAP7_75t_L g494 ( .A(n_52), .B(n_177), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_53), .B(n_161), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_54), .B(n_159), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_55), .B(n_161), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_56), .A2(n_152), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_57), .B(n_143), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_58), .B(n_143), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_59), .A2(n_152), .B(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_60), .A2(n_98), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
AO21x1_ASAP7_75t_L g219 ( .A1(n_61), .A2(n_152), .B(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g545 ( .A(n_62), .B(n_178), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_63), .B(n_143), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_64), .B(n_161), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_65), .B(n_143), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_66), .A2(n_78), .B1(n_776), .B2(n_777), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_66), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_67), .B(n_161), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_68), .A2(n_93), .B1(n_152), .B2(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g232 ( .A(n_69), .B(n_178), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_70), .B(n_159), .Y(n_542) );
INVx1_ASAP7_75t_L g148 ( .A(n_71), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_71), .Y(n_154) );
AND2x2_ASAP7_75t_L g200 ( .A(n_72), .B(n_169), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_73), .B(n_161), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_74), .A2(n_152), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_75), .A2(n_152), .B(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_76), .A2(n_152), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g517 ( .A(n_77), .B(n_178), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_78), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_79), .B(n_177), .Y(n_476) );
INVx1_ASAP7_75t_L g119 ( .A(n_80), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_80), .B(n_118), .Y(n_785) );
AND2x2_ASAP7_75t_L g168 ( .A(n_81), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_82), .B(n_143), .Y(n_188) );
AND2x2_ASAP7_75t_L g465 ( .A(n_83), .B(n_138), .Y(n_465) );
INVxp33_ASAP7_75t_L g791 ( .A(n_84), .Y(n_791) );
AND2x2_ASAP7_75t_L g218 ( .A(n_85), .B(n_163), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_87), .B(n_161), .Y(n_187) );
AND2x2_ASAP7_75t_L g212 ( .A(n_88), .B(n_169), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_90), .B(n_159), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_91), .A2(n_152), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_92), .B(n_161), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_94), .A2(n_152), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_95), .B(n_159), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_96), .B(n_159), .Y(n_175) );
BUFx2_ASAP7_75t_L g544 ( .A(n_97), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_98), .Y(n_123) );
BUFx2_ASAP7_75t_L g106 ( .A(n_99), .Y(n_106) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_99), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_100), .A2(n_152), .B(n_157), .Y(n_151) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_782), .B(n_790), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_121), .B(n_770), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_108), .A2(n_774), .B(n_779), .Y(n_773) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g781 ( .A(n_113), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g130 ( .A(n_114), .B(n_115), .Y(n_130) );
AND2x6_ASAP7_75t_SL g759 ( .A(n_114), .B(n_116), .Y(n_759) );
OR2x2_ASAP7_75t_L g769 ( .A(n_114), .B(n_116), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_760), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_122), .A2(n_761), .B(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_131), .B1(n_453), .B2(n_756), .Y(n_126) );
BUFx4f_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
OAI22x1_ASAP7_75t_L g761 ( .A1(n_128), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
CKINVDCx11_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g762 ( .A(n_131), .Y(n_762) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_374), .Y(n_131) );
NOR3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_286), .C(n_326), .Y(n_132) );
OAI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_201), .B1(n_250), .B2(n_265), .C(n_268), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_165), .Y(n_135) );
INVx2_ASAP7_75t_L g283 ( .A(n_136), .Y(n_283) );
AND2x2_ASAP7_75t_L g313 ( .A(n_136), .B(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g251 ( .A(n_137), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g258 ( .A(n_137), .B(n_191), .Y(n_258) );
INVx2_ASAP7_75t_L g264 ( .A(n_137), .Y(n_264) );
AND2x2_ASAP7_75t_L g273 ( .A(n_137), .B(n_167), .Y(n_273) );
INVx1_ASAP7_75t_L g289 ( .A(n_137), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_137), .B(n_335), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_138), .A2(n_539), .B(n_540), .Y(n_538) );
BUFx4f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x4_ASAP7_75t_L g163 ( .A(n_140), .B(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_140), .B(n_164), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_151), .B(n_163), .Y(n_141) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
AND2x6_ASAP7_75t_L g161 ( .A(n_145), .B(n_154), .Y(n_161) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g159 ( .A(n_147), .B(n_156), .Y(n_159) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
AND2x2_ASAP7_75t_L g155 ( .A(n_150), .B(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_150), .Y(n_482) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
BUFx3_ASAP7_75t_L g483 ( .A(n_153), .Y(n_483) );
INVx2_ASAP7_75t_L g489 ( .A(n_154), .Y(n_489) );
AND2x4_ASAP7_75t_L g485 ( .A(n_155), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g481 ( .A(n_156), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_161), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_162), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_162), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_162), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_162), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_162), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_162), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_162), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_162), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_162), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_162), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_162), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_162), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_162), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_SL g182 ( .A(n_163), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_163), .B(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_163), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_163), .A2(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_179), .Y(n_165) );
INVx4_ASAP7_75t_L g254 ( .A(n_166), .Y(n_254) );
AND2x2_ASAP7_75t_L g285 ( .A(n_166), .B(n_192), .Y(n_285) );
AND2x2_ASAP7_75t_L g361 ( .A(n_166), .B(n_335), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_166), .B(n_191), .Y(n_403) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_167), .B(n_191), .Y(n_290) );
AND2x2_ASAP7_75t_L g314 ( .A(n_167), .B(n_192), .Y(n_314) );
BUFx2_ASAP7_75t_L g330 ( .A(n_167), .Y(n_330) );
NOR2x1_ASAP7_75t_SL g433 ( .A(n_167), .B(n_335), .Y(n_433) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_171), .Y(n_167) );
INVx3_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_170), .A2(n_468), .B(n_474), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_177), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_177), .Y(n_199) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_177), .A2(n_238), .B(n_242), .Y(n_237) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_177), .A2(n_238), .B(n_242), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_177), .A2(n_460), .B(n_461), .Y(n_459) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_177), .A2(n_478), .B(n_484), .Y(n_477) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_179), .A2(n_377), .B1(n_379), .B2(n_381), .C(n_386), .Y(n_376) );
AND2x2_ASAP7_75t_L g396 ( .A(n_179), .B(n_289), .Y(n_396) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_191), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
INVx1_ASAP7_75t_L g305 ( .A(n_181), .Y(n_305) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_182), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g335 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_191), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g274 ( .A(n_191), .B(n_262), .Y(n_274) );
INVx2_ASAP7_75t_L g316 ( .A(n_191), .Y(n_316) );
AND2x2_ASAP7_75t_L g449 ( .A(n_191), .B(n_264), .Y(n_449) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_192), .Y(n_306) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_199), .B(n_200), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_198), .Y(n_193) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_199), .A2(n_528), .B(n_534), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_233), .C(n_248), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_213), .Y(n_202) );
INVx2_ASAP7_75t_L g363 ( .A(n_203), .Y(n_363) );
AND2x2_ASAP7_75t_L g408 ( .A(n_203), .B(n_285), .Y(n_408) );
BUFx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g353 ( .A(n_204), .Y(n_353) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_204), .B(n_280), .Y(n_368) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_204) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_211), .A2(n_226), .B(n_232), .Y(n_225) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_211), .A2(n_226), .B(n_232), .Y(n_245) );
AO21x1_ASAP7_75t_SL g510 ( .A1(n_211), .A2(n_511), .B(n_517), .Y(n_510) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_211), .A2(n_511), .B(n_517), .Y(n_568) );
INVx2_ASAP7_75t_L g322 ( .A(n_213), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_213), .B(n_352), .Y(n_378) );
AND2x4_ASAP7_75t_L g411 ( .A(n_213), .B(n_358), .Y(n_411) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
AND2x2_ASAP7_75t_L g249 ( .A(n_214), .B(n_244), .Y(n_249) );
OR2x2_ASAP7_75t_L g279 ( .A(n_214), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_214), .B(n_300), .Y(n_348) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g293 ( .A(n_215), .Y(n_293) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g267 ( .A(n_216), .Y(n_267) );
OAI21x1_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_219), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_218), .Y(n_224) );
INVx2_ASAP7_75t_L g280 ( .A(n_225), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_231), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_233), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_243), .Y(n_234) );
AND2x2_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g321 ( .A(n_235), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g406 ( .A(n_235), .Y(n_406) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g266 ( .A(n_236), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g385 ( .A(n_236), .B(n_245), .Y(n_385) );
AND2x2_ASAP7_75t_L g389 ( .A(n_236), .B(n_255), .Y(n_389) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g358 ( .A(n_237), .Y(n_358) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_237), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_243), .B(n_266), .Y(n_342) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_244), .B(n_267), .Y(n_452) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g256 ( .A(n_245), .B(n_247), .Y(n_256) );
AND2x2_ASAP7_75t_L g338 ( .A(n_245), .B(n_300), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_245), .B(n_246), .Y(n_357) );
BUFx2_ASAP7_75t_L g278 ( .A(n_246), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_246), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx3_ASAP7_75t_L g255 ( .A(n_247), .Y(n_255) );
INVxp67_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
INVx1_ASAP7_75t_L g271 ( .A(n_249), .Y(n_271) );
AND2x2_ASAP7_75t_L g307 ( .A(n_249), .B(n_278), .Y(n_307) );
NAND2xp33_ASAP7_75t_L g388 ( .A(n_249), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g425 ( .A(n_249), .B(n_426), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B1(n_256), .B2(n_257), .C(n_259), .Y(n_250) );
AND2x2_ASAP7_75t_L g354 ( .A(n_251), .B(n_254), .Y(n_354) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_251), .B(n_314), .Y(n_373) );
AND2x2_ASAP7_75t_L g391 ( .A(n_251), .B(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g446 ( .A(n_251), .B(n_285), .Y(n_446) );
INVx1_ASAP7_75t_L g262 ( .A(n_252), .Y(n_262) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_252), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_253), .Y(n_398) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_254), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_254), .B(n_305), .Y(n_380) );
AND2x2_ASAP7_75t_L g347 ( .A(n_255), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g383 ( .A(n_255), .Y(n_383) );
AND2x2_ASAP7_75t_L g292 ( .A(n_256), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_256), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g434 ( .A(n_256), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_256), .B(n_358), .Y(n_444) );
AND2x4_ASAP7_75t_L g360 ( .A(n_257), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g431 ( .A(n_258), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
OR2x2_ASAP7_75t_L g302 ( .A(n_263), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g309 ( .A(n_264), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g340 ( .A(n_264), .B(n_314), .Y(n_340) );
AND2x2_ASAP7_75t_L g414 ( .A(n_264), .B(n_335), .Y(n_414) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g362 ( .A(n_266), .B(n_363), .Y(n_362) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_266), .A2(n_428), .A3(n_430), .B1(n_431), .B2(n_434), .Y(n_427) );
AND2x4_ASAP7_75t_L g299 ( .A(n_267), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g397 ( .A(n_267), .B(n_300), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B1(n_275), .B2(n_281), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_SL g386 ( .A1(n_270), .A2(n_284), .B(n_387), .C(n_388), .Y(n_386) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g370 ( .A(n_271), .B(n_298), .Y(n_370) );
INVx1_ASAP7_75t_SL g441 ( .A(n_272), .Y(n_441) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x4_ASAP7_75t_L g344 ( .A(n_274), .B(n_283), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_274), .A2(n_423), .B1(n_424), .B2(n_425), .C(n_427), .Y(n_422) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_279), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_282), .A2(n_312), .B1(n_365), .B2(n_366), .Y(n_364) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_283), .A2(n_401), .B(n_409), .C(n_422), .Y(n_400) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g320 ( .A(n_285), .B(n_289), .Y(n_320) );
OAI211xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_291), .B(n_294), .C(n_323), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g317 ( .A(n_289), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g437 ( .A(n_289), .B(n_433), .Y(n_437) );
OAI32xp33_ASAP7_75t_L g394 ( .A1(n_290), .A2(n_395), .A3(n_397), .B1(n_398), .B2(n_399), .Y(n_394) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_293), .B(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_301), .B1(n_307), .B2(n_308), .C(n_311), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g451 ( .A(n_298), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_299), .B(n_363), .Y(n_365) );
A2O1A1O1Ixp25_ASAP7_75t_L g436 ( .A1(n_299), .A2(n_368), .B(n_384), .C(n_430), .D(n_437), .Y(n_436) );
AOI31xp33_ASAP7_75t_L g438 ( .A1(n_299), .A2(n_320), .A3(n_430), .B(n_437), .Y(n_438) );
AND2x2_ASAP7_75t_L g352 ( .A(n_300), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_302), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_L g429 ( .A(n_304), .Y(n_429) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g424 ( .A(n_305), .B(n_316), .Y(n_424) );
INVx1_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
AND2x2_ASAP7_75t_L g324 ( .A(n_308), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AOI31xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .A3(n_319), .B(n_321), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_314), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g447 ( .A(n_314), .B(n_393), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g392 ( .A(n_316), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g418 ( .A(n_316), .Y(n_418) );
INVxp67_ASAP7_75t_L g387 ( .A(n_317), .Y(n_387) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g325 ( .A(n_321), .Y(n_325) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND3xp33_ASAP7_75t_SL g326 ( .A(n_327), .B(n_343), .C(n_359), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_336), .B1(n_340), .B2(n_341), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g413 ( .A(n_330), .Y(n_413) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_334), .Y(n_393) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_334), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_334), .B(n_403), .Y(n_420) );
NAND2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B1(n_354), .B2(n_355), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_352), .A2(n_357), .B1(n_391), .B2(n_392), .C(n_394), .Y(n_390) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
AND2x2_ASAP7_75t_L g367 ( .A(n_358), .B(n_368), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_SL g415 ( .A1(n_358), .A2(n_416), .B(n_420), .C(n_421), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_364), .C(n_369), .Y(n_359) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g421 ( .A(n_368), .Y(n_421) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B(n_372), .Y(n_369) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_400), .C(n_435), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_376), .B(n_390), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
INVxp67_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g407 ( .A(n_397), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_407), .B2(n_408), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_415), .Y(n_409) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g448 ( .A(n_433), .B(n_449), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_439), .B2(n_442), .C(n_445), .Y(n_435) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI31xp33_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_447), .A3(n_448), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_SL g763 ( .A(n_453), .Y(n_763) );
OAI22xp5_ASAP7_75t_SL g774 ( .A1(n_453), .A2(n_763), .B1(n_775), .B2(n_778), .Y(n_774) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_454), .B(n_652), .Y(n_453) );
NOR3xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_561), .C(n_593), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_490), .B1(n_518), .B2(n_535), .C(n_546), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g524 ( .A(n_458), .B(n_467), .Y(n_524) );
INVx4_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_458), .B(n_526), .Y(n_592) );
BUFx2_ASAP7_75t_L g602 ( .A(n_458), .Y(n_602) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_458), .B(n_607), .Y(n_668) );
AND2x2_ASAP7_75t_L g677 ( .A(n_458), .B(n_605), .Y(n_677) );
OR2x2_ASAP7_75t_L g685 ( .A(n_458), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g711 ( .A(n_458), .B(n_550), .Y(n_711) );
AND2x4_ASAP7_75t_L g730 ( .A(n_458), .B(n_731), .Y(n_730) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
INVx2_ASAP7_75t_SL g643 ( .A(n_466), .Y(n_643) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_527), .Y(n_550) );
INVx2_ASAP7_75t_L g577 ( .A(n_467), .Y(n_577) );
INVx2_ASAP7_75t_L g607 ( .A(n_467), .Y(n_607) );
AND2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_526), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
AND2x2_ASAP7_75t_L g551 ( .A(n_475), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g574 ( .A(n_475), .Y(n_574) );
BUFx3_ASAP7_75t_L g588 ( .A(n_475), .Y(n_588) );
AND2x2_ASAP7_75t_L g617 ( .A(n_475), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x4_ASAP7_75t_L g522 ( .A(n_476), .B(n_477), .Y(n_522) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NOR2x1p5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g623 ( .A(n_490), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
OR2x2_ASAP7_75t_L g734 ( .A(n_491), .B(n_535), .Y(n_734) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g590 ( .A(n_492), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_492), .B(n_501), .Y(n_651) );
OR2x2_ASAP7_75t_L g749 ( .A(n_492), .B(n_671), .Y(n_749) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_536), .Y(n_560) );
OR2x2_ASAP7_75t_SL g570 ( .A(n_493), .B(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_493), .Y(n_632) );
NAND2x1_ASAP7_75t_L g638 ( .A(n_493), .B(n_537), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_493), .B(n_503), .Y(n_663) );
OR2x2_ASAP7_75t_L g684 ( .A(n_493), .B(n_567), .Y(n_684) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g579 ( .A(n_501), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_501), .A2(n_673), .B(n_676), .C(n_678), .Y(n_672) );
AND2x2_ASAP7_75t_L g745 ( .A(n_501), .B(n_521), .Y(n_745) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
INVx1_ASAP7_75t_L g612 ( .A(n_502), .Y(n_612) );
AND2x2_ASAP7_75t_L g682 ( .A(n_502), .B(n_537), .Y(n_682) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
OR2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_537), .Y(n_571) );
INVx1_ASAP7_75t_L g587 ( .A(n_503), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_503), .B(n_510), .Y(n_599) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_503), .Y(n_705) );
NOR2x1_ASAP7_75t_SL g536 ( .A(n_510), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
OR2x2_ASAP7_75t_L g669 ( .A(n_520), .B(n_604), .Y(n_669) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_521), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g751 ( .A(n_521), .B(n_648), .Y(n_751) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g596 ( .A(n_522), .B(n_577), .Y(n_596) );
AND2x2_ASAP7_75t_L g692 ( .A(n_522), .B(n_605), .Y(n_692) );
INVx1_ASAP7_75t_L g609 ( .A(n_523), .Y(n_609) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g659 ( .A(n_524), .Y(n_659) );
INVx2_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g606 ( .A(n_526), .Y(n_606) );
INVx1_ASAP7_75t_L g731 ( .A(n_526), .Y(n_731) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_527), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
OR2x2_ASAP7_75t_L g702 ( .A(n_535), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g557 ( .A(n_537), .Y(n_557) );
OR2x2_ASAP7_75t_L g580 ( .A(n_537), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g591 ( .A(n_537), .B(n_567), .Y(n_591) );
AND2x2_ASAP7_75t_L g665 ( .A(n_537), .B(n_581), .Y(n_665) );
BUFx2_ASAP7_75t_L g748 ( .A(n_537), .Y(n_748) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_545), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_553), .B(n_558), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g700 ( .A(n_549), .B(n_622), .Y(n_700) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g559 ( .A(n_550), .B(n_552), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_551), .B(n_621), .Y(n_722) );
INVx1_ASAP7_75t_L g752 ( .A(n_551), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_552), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_552), .B(n_688), .Y(n_725) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
AND2x4_ASAP7_75t_SL g589 ( .A(n_555), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_555), .B(n_583), .Y(n_736) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_556), .B(n_638), .Y(n_694) );
AND2x2_ASAP7_75t_L g712 ( .A(n_556), .B(n_665), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_557), .B(n_599), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_557), .A2(n_603), .B(n_645), .C(n_650), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_559), .A2(n_632), .B1(n_740), .B2(n_746), .C(n_750), .Y(n_739) );
INVx1_ASAP7_75t_SL g727 ( .A(n_560), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_572), .B1(n_578), .B2(n_582), .C(n_793), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g637 ( .A(n_566), .Y(n_637) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g642 ( .A(n_567), .B(n_587), .Y(n_642) );
INVx2_ASAP7_75t_L g675 ( .A(n_567), .Y(n_675) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI32xp33_ASAP7_75t_L g726 ( .A1(n_570), .A2(n_617), .A3(n_648), .B1(n_727), .B2(n_728), .Y(n_726) );
OR2x2_ASAP7_75t_L g697 ( .A(n_571), .B(n_684), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_572), .Y(n_707) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
AND2x2_ASAP7_75t_L g693 ( .A(n_573), .B(n_668), .Y(n_693) );
OR2x2_ASAP7_75t_L g724 ( .A(n_573), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_574), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g618 ( .A(n_577), .Y(n_618) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_SL g583 ( .A(n_580), .Y(n_583) );
OR2x2_ASAP7_75t_L g670 ( .A(n_580), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_581), .B(n_599), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_581), .B(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g717 ( .A(n_581), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_589), .C(n_592), .Y(n_582) );
AND2x2_ASAP7_75t_L g732 ( .A(n_584), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g658 ( .A(n_588), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_588), .B(n_592), .Y(n_679) );
AND2x2_ASAP7_75t_L g710 ( .A(n_588), .B(n_711), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_590), .A2(n_721), .B(n_723), .C(n_726), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g594 ( .A1(n_591), .A2(n_595), .B1(n_597), .B2(n_600), .C1(n_608), .C2(n_610), .Y(n_594) );
AND2x2_ASAP7_75t_L g662 ( .A(n_591), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g595 ( .A(n_592), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g616 ( .A(n_592), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_613), .C(n_634), .D(n_644), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_596), .B(n_602), .Y(n_656) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g664 ( .A(n_599), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_SL g671 ( .A(n_599), .Y(n_671) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_601), .A2(n_635), .B(n_639), .C(n_643), .Y(n_634) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_602), .B(n_617), .Y(n_738) );
OR2x2_ASAP7_75t_L g742 ( .A(n_602), .B(n_628), .Y(n_742) );
INVx1_ASAP7_75t_L g715 ( .A(n_603), .Y(n_715) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g649 ( .A(n_606), .Y(n_649) );
INVx1_ASAP7_75t_L g629 ( .A(n_607), .Y(n_629) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_609), .B(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g633 ( .A(n_611), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .A3(n_617), .B1(n_619), .B2(n_623), .C1(n_624), .C2(n_630), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_SL g695 ( .A1(n_616), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g718 ( .A(n_617), .Y(n_718) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g676 ( .A(n_622), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_628), .Y(n_698) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx3_ASAP7_75t_L g641 ( .A(n_638), .Y(n_641) );
OR2x2_ASAP7_75t_L g709 ( .A(n_638), .B(n_671), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_638), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_SL g741 ( .A(n_642), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_643), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g746 ( .A(n_651), .B(n_747), .C(n_749), .Y(n_746) );
NOR3xp33_ASAP7_75t_SL g652 ( .A(n_653), .B(n_690), .C(n_719), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_672), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_666), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g699 ( .A1(n_655), .A2(n_677), .A3(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx2_ASAP7_75t_L g714 ( .A(n_662), .Y(n_714) );
INVx1_ASAP7_75t_L g689 ( .A(n_664), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g716 ( .A(n_674), .B(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g755 ( .A(n_675), .Y(n_755) );
OAI22xp33_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B1(n_685), .B2(n_689), .Y(n_678) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_684), .Y(n_696) );
OR2x2_ASAP7_75t_L g747 ( .A(n_684), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_699), .C(n_706), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B(n_694), .C(n_695), .Y(n_691) );
INVx2_ASAP7_75t_L g728 ( .A(n_692), .Y(n_728) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_716), .B2(n_718), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_729), .C(n_739), .Y(n_719) );
INVxp33_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_735), .B2(n_737), .Y(n_729) );
INVx2_ASAP7_75t_L g743 ( .A(n_730), .Y(n_743) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp33_ASAP7_75t_SL g750 ( .A1(n_749), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx4_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
CKINVDCx6p67_ASAP7_75t_R g764 ( .A(n_757), .Y(n_764) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_775), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_784), .B(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_SL g784 ( .A(n_785), .B(n_786), .Y(n_784) );
endmodule