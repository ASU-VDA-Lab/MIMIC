module real_aes_1343_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g237 ( .A(n_0), .B(n_159), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_1), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g152 ( .A(n_2), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_3), .B(n_165), .Y(n_178) );
NAND2xp33_ASAP7_75t_SL g229 ( .A(n_4), .B(n_163), .Y(n_229) );
INVx1_ASAP7_75t_L g210 ( .A(n_5), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_6), .B(n_183), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_7), .A2(n_127), .B1(n_128), .B2(n_130), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_7), .Y(n_127) );
INVx1_ASAP7_75t_L g536 ( .A(n_8), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_9), .Y(n_121) );
AND2x2_ASAP7_75t_L g176 ( .A(n_10), .B(n_169), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_11), .Y(n_503) );
INVx2_ASAP7_75t_L g170 ( .A(n_12), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_13), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_14), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_14), .B(n_27), .Y(n_732) );
INVx1_ASAP7_75t_L g564 ( .A(n_15), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_16), .A2(n_27), .B1(n_786), .B2(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_16), .Y(n_818) );
AOI221x1_ASAP7_75t_L g223 ( .A1(n_17), .A2(n_147), .B1(n_224), .B2(n_226), .C(n_228), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_18), .B(n_165), .Y(n_198) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g562 ( .A(n_20), .Y(n_562) );
INVx1_ASAP7_75t_SL g485 ( .A(n_21), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_22), .B(n_166), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_23), .A2(n_147), .B(n_180), .Y(n_179) );
AOI221xp5_ASAP7_75t_SL g190 ( .A1(n_24), .A2(n_40), .B1(n_147), .B2(n_165), .C(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_25), .B(n_159), .Y(n_181) );
AOI33xp33_ASAP7_75t_L g522 ( .A1(n_26), .A2(n_54), .A3(n_213), .B1(n_219), .B2(n_523), .B3(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g786 ( .A(n_27), .Y(n_786) );
INVx1_ASAP7_75t_L g496 ( .A(n_28), .Y(n_496) );
OR2x2_ASAP7_75t_L g171 ( .A(n_29), .B(n_94), .Y(n_171) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_29), .A2(n_94), .B(n_170), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_30), .B(n_155), .Y(n_202) );
INVxp67_ASAP7_75t_L g222 ( .A(n_31), .Y(n_222) );
AND2x2_ASAP7_75t_L g253 ( .A(n_32), .B(n_168), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_33), .B(n_211), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_34), .A2(n_147), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_35), .B(n_155), .Y(n_192) );
AND2x2_ASAP7_75t_L g148 ( .A(n_36), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g163 ( .A(n_36), .B(n_152), .Y(n_163) );
INVx1_ASAP7_75t_L g218 ( .A(n_36), .Y(n_218) );
OR2x6_ASAP7_75t_L g115 ( .A(n_37), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_38), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_39), .B(n_211), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_41), .A2(n_183), .B1(n_227), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_42), .B(n_554), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_43), .A2(n_84), .B1(n_147), .B2(n_216), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_44), .B(n_166), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_45), .B(n_159), .Y(n_251) );
INVx1_ASAP7_75t_L g794 ( .A(n_46), .Y(n_794) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_47), .B(n_88), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_48), .B(n_203), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_49), .B(n_166), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_50), .Y(n_549) );
AND2x2_ASAP7_75t_L g240 ( .A(n_51), .B(n_168), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_52), .B(n_168), .Y(n_194) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_52), .B(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_53), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_55), .B(n_166), .Y(n_514) );
INVx1_ASAP7_75t_L g151 ( .A(n_56), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_56), .Y(n_161) );
AND2x2_ASAP7_75t_L g515 ( .A(n_57), .B(n_168), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_58), .A2(n_77), .B1(n_211), .B2(n_216), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_59), .B(n_211), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_60), .B(n_165), .Y(n_252) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_61), .A2(n_126), .B1(n_131), .B2(n_132), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_61), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_62), .B(n_227), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g474 ( .A1(n_63), .A2(n_216), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g172 ( .A(n_64), .B(n_168), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_65), .B(n_155), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_66), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_67), .B(n_169), .Y(n_205) );
INVx1_ASAP7_75t_L g559 ( .A(n_68), .Y(n_559) );
XNOR2xp5_ASAP7_75t_L g128 ( .A(n_69), .B(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_70), .A2(n_147), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g513 ( .A(n_71), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_72), .B(n_155), .Y(n_182) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_73), .B(n_203), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_74), .A2(n_216), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g149 ( .A(n_75), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_75), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_76), .B(n_211), .Y(n_525) );
AND2x2_ASAP7_75t_L g487 ( .A(n_78), .B(n_226), .Y(n_487) );
INVx1_ASAP7_75t_L g560 ( .A(n_79), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_80), .A2(n_216), .B(n_484), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_81), .A2(n_216), .B(n_286), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_82), .B(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_83), .A2(n_87), .B1(n_165), .B2(n_211), .Y(n_288) );
INVx1_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_86), .B(n_226), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_89), .A2(n_216), .B1(n_520), .B2(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_90), .B(n_159), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_91), .B(n_159), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_92), .B(n_797), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_93), .A2(n_147), .B(n_153), .Y(n_146) );
INVx1_ASAP7_75t_L g476 ( .A(n_95), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_96), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g526 ( .A(n_97), .B(n_226), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_98), .A2(n_494), .B(n_495), .C(n_497), .Y(n_493) );
INVxp67_ASAP7_75t_L g225 ( .A(n_99), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_100), .B(n_165), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_101), .B(n_155), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_102), .A2(n_147), .B(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_SL g792 ( .A(n_103), .Y(n_792) );
BUFx2_ASAP7_75t_L g804 ( .A(n_103), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_104), .B(n_166), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_122), .B(n_829), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_108), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_119), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g798 ( .A(n_112), .Y(n_798) );
NOR2x1_ASAP7_75t_R g803 ( .A(n_112), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_113), .Y(n_787) );
OR2x2_ASAP7_75t_L g795 ( .A(n_113), .B(n_115), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
OAI32xp33_ASAP7_75t_L g799 ( .A1(n_115), .A2(n_800), .A3(n_801), .B1(n_802), .B2(n_833), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_805), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_788), .B(n_799), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_133), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_125), .Y(n_828) );
INVxp33_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
INVx1_ASAP7_75t_L g130 ( .A(n_128), .Y(n_130) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_134), .Y(n_827) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_462), .Y(n_134) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_401), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_294), .C(n_345), .Y(n_137) );
OAI211xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_184), .B(n_241), .C(n_272), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_173), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_143), .B(n_246), .Y(n_409) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g254 ( .A(n_144), .B(n_175), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_144), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g271 ( .A(n_144), .B(n_261), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_144), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_144), .B(n_284), .Y(n_308) );
INVx2_ASAP7_75t_L g334 ( .A(n_144), .Y(n_334) );
AND2x4_ASAP7_75t_L g343 ( .A(n_144), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g448 ( .A(n_144), .B(n_315), .Y(n_448) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_167), .B(n_172), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_164), .Y(n_145) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
AND2x6_ASAP7_75t_L g159 ( .A(n_149), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
AND2x4_ASAP7_75t_L g216 ( .A(n_150), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x4_ASAP7_75t_L g155 ( .A(n_151), .B(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_158), .B(n_162), .Y(n_153) );
INVxp67_ASAP7_75t_L g565 ( .A(n_155), .Y(n_565) );
AND2x4_ASAP7_75t_L g166 ( .A(n_156), .B(n_160), .Y(n_166) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVxp67_ASAP7_75t_L g563 ( .A(n_159), .Y(n_563) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_162), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_162), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_162), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_162), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_162), .A2(n_250), .B(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_162), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_162), .A2(n_477), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_162), .A2(n_477), .B(n_513), .C(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g520 ( .A(n_162), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_162), .A2(n_477), .B(n_536), .C(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_162), .A2(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_162), .B(n_183), .Y(n_566) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g165 ( .A(n_163), .B(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_163), .Y(n_497) );
INVx1_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_167), .A2(n_247), .B(n_253), .Y(n_246) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_167), .A2(n_247), .B(n_253), .Y(n_261) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_167), .A2(n_481), .B(n_487), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_168), .A2(n_190), .B(n_194), .Y(n_189) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_170), .B(n_171), .Y(n_169) );
AND2x4_ASAP7_75t_L g183 ( .A(n_170), .B(n_171), .Y(n_183) );
AND2x2_ASAP7_75t_L g332 ( .A(n_173), .B(n_333), .Y(n_332) );
OAI32xp33_ASAP7_75t_L g415 ( .A1(n_173), .A2(n_337), .A3(n_341), .B1(n_348), .B2(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_173), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g269 ( .A(n_174), .B(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_174), .B(n_264), .C(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g368 ( .A(n_174), .B(n_271), .Y(n_368) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
INVx5_ASAP7_75t_L g293 ( .A(n_175), .Y(n_293) );
AND2x4_ASAP7_75t_L g349 ( .A(n_175), .B(n_261), .Y(n_349) );
OR2x2_ASAP7_75t_L g364 ( .A(n_175), .B(n_284), .Y(n_364) );
OR2x2_ASAP7_75t_L g390 ( .A(n_175), .B(n_246), .Y(n_390) );
AND2x2_ASAP7_75t_L g398 ( .A(n_175), .B(n_344), .Y(n_398) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_175), .B(n_343), .Y(n_423) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_183), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_183), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_183), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_183), .B(n_225), .Y(n_224) );
NOR3xp33_ASAP7_75t_L g228 ( .A(n_183), .B(n_229), .C(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_183), .A2(n_474), .B(n_479), .Y(n_473) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_185), .B(n_343), .Y(n_419) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_186), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OR2x6_ASAP7_75t_SL g243 ( .A(n_187), .B(n_244), .Y(n_243) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g268 ( .A(n_188), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_188), .B(n_303), .Y(n_321) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_188), .Y(n_459) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
AND2x2_ASAP7_75t_L g301 ( .A(n_189), .B(n_232), .Y(n_301) );
INVx2_ASAP7_75t_L g329 ( .A(n_189), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_189), .B(n_196), .Y(n_370) );
BUFx3_ASAP7_75t_L g394 ( .A(n_189), .Y(n_394) );
OR2x2_ASAP7_75t_L g406 ( .A(n_189), .B(n_196), .Y(n_406) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_189), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_195), .A2(n_437), .B1(n_440), .B2(n_441), .Y(n_436) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
INVx1_ASAP7_75t_L g264 ( .A(n_196), .Y(n_264) );
OR2x2_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_196), .B(n_207), .Y(n_299) );
AND2x4_ASAP7_75t_L g304 ( .A(n_196), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g313 ( .A(n_196), .Y(n_313) );
OR2x2_ASAP7_75t_L g319 ( .A(n_196), .B(n_207), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_196), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_196), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_196), .B(n_301), .Y(n_435) );
OR2x2_ASAP7_75t_L g451 ( .A(n_196), .B(n_354), .Y(n_451) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_205), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_203), .Y(n_197) );
INVx2_ASAP7_75t_SL g286 ( .A(n_203), .Y(n_286) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_203), .A2(n_534), .B(n_538), .Y(n_533) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g227 ( .A(n_204), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_206), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g277 ( .A(n_206), .Y(n_277) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_206), .B(n_268), .Y(n_384) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_231), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_207), .B(n_232), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_207), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_207), .B(n_276), .Y(n_280) );
INVx3_ASAP7_75t_L g305 ( .A(n_207), .Y(n_305) );
INVx1_ASAP7_75t_L g338 ( .A(n_207), .Y(n_338) );
AND2x2_ASAP7_75t_L g418 ( .A(n_207), .B(n_282), .Y(n_418) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_223), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B1(n_216), .B2(n_221), .Y(n_208) );
INVx1_ASAP7_75t_L g506 ( .A(n_211), .Y(n_506) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g547 ( .A(n_212), .Y(n_547) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
OR2x6_ASAP7_75t_L g477 ( .A(n_213), .B(n_220), .Y(n_477) );
INVxp33_ASAP7_75t_L g523 ( .A(n_213), .Y(n_523) );
INVx1_ASAP7_75t_L g548 ( .A(n_215), .Y(n_548) );
INVxp67_ASAP7_75t_L g504 ( .A(n_216), .Y(n_504) );
NOR2x1p5_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g524 ( .A(n_219), .Y(n_524) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_226), .A2(n_493), .B1(n_498), .B2(n_499), .Y(n_492) );
INVx3_ASAP7_75t_L g499 ( .A(n_226), .Y(n_499) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_227), .A2(n_234), .B(n_240), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_227), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_230), .B(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_230), .A2(n_477), .B1(n_559), .B2(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_232), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g303 ( .A(n_232), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_232), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g354 ( .A(n_232), .B(n_276), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_232), .B(n_305), .Y(n_371) );
INVx1_ASAP7_75t_L g377 ( .A(n_232), .Y(n_377) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_239), .Y(n_234) );
AOI222xp33_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_245), .B1(n_255), .B2(n_262), .C1(n_265), .C2(n_269), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_254), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_246), .B(n_315), .Y(n_366) );
AND2x4_ASAP7_75t_L g382 ( .A(n_246), .B(n_293), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_252), .Y(n_247) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g307 ( .A(n_258), .B(n_308), .Y(n_307) );
AOI222xp33_ASAP7_75t_L g272 ( .A1(n_259), .A2(n_273), .B1(n_278), .B2(n_283), .C1(n_291), .C2(n_832), .Y(n_272) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g411 ( .A(n_260), .B(n_315), .Y(n_411) );
OR2x2_ASAP7_75t_L g454 ( .A(n_260), .B(n_360), .Y(n_454) );
AND2x2_ASAP7_75t_L g283 ( .A(n_261), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_261), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_262), .A2(n_373), .B(n_378), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g400 ( .A(n_264), .Y(n_400) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g330 ( .A(n_269), .Y(n_330) );
AND2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g323 ( .A(n_270), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI31xp33_ASAP7_75t_L g365 ( .A1(n_273), .A2(n_291), .A3(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_274), .A2(n_324), .B(n_368), .C(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
OR2x2_ASAP7_75t_L g356 ( .A(n_275), .B(n_305), .Y(n_356) );
INVx2_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
BUFx2_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_284), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_290), .Y(n_285) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_286), .A2(n_518), .B(n_526), .Y(n_517) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_286), .A2(n_518), .B(n_526), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_293), .B(n_350), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_306), .B(n_309), .C(n_331), .Y(n_294) );
INVxp33_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_302), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g335 ( .A(n_299), .B(n_328), .Y(n_335) );
OR2x2_ASAP7_75t_L g311 ( .A(n_300), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g341 ( .A(n_300), .B(n_315), .Y(n_341) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g417 ( .A(n_301), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g440 ( .A(n_302), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_304), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_304), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g452 ( .A(n_304), .B(n_328), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_304), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g395 ( .A(n_305), .B(n_377), .Y(n_395) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AOI322xp5_ASAP7_75t_L g449 ( .A1(n_308), .A2(n_328), .A3(n_382), .B1(n_407), .B2(n_450), .C1(n_452), .C2(n_453), .Y(n_449) );
AOI211xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_314), .B(n_316), .C(n_325), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_312), .B(n_340), .Y(n_362) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g327 ( .A(n_313), .B(n_328), .Y(n_327) );
NOR2x1p5_ASAP7_75t_L g393 ( .A(n_313), .B(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_313), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_314), .A2(n_332), .B(n_335), .C(n_336), .Y(n_331) );
AND2x4_ASAP7_75t_L g350 ( .A(n_315), .B(n_334), .Y(n_350) );
INVx2_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_315), .B(n_349), .Y(n_380) );
AND2x2_ASAP7_75t_L g422 ( .A(n_315), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_315), .B(n_439), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_315), .B(n_343), .Y(n_461) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B(n_322), .Y(n_316) );
AND2x2_ASAP7_75t_L g412 ( .A(n_318), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_333), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g427 ( .A(n_333), .Y(n_427) );
O2A1O1Ixp33_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_341), .C(n_342), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_340), .Y(n_424) );
INVx3_ASAP7_75t_SL g439 ( .A(n_343), .Y(n_439) );
NAND5xp2_ASAP7_75t_L g345 ( .A(n_346), .B(n_365), .C(n_372), .D(n_385), .E(n_396), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_351), .B1(n_355), .B2(n_357), .C1(n_361), .C2(n_363), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_348), .A2(n_429), .B1(n_433), .B2(n_434), .Y(n_428) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_350), .Y(n_378) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_359), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_360), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g397 ( .A(n_360), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g408 ( .A(n_360), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g438 ( .A(n_364), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_371), .Y(n_386) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B(n_383), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_382), .A2(n_386), .B1(n_387), .B2(n_391), .Y(n_385) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g399 ( .A(n_384), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g404 ( .A(n_386), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_SL g432 ( .A(n_395), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_420), .C(n_443), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_403), .B(n_419), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g444 ( .A(n_406), .B(n_432), .Y(n_444) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OAI321xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .A3(n_425), .B1(n_427), .B2(n_428), .C(n_436), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_434), .A2(n_456), .B1(n_460), .B2(n_461), .Y(n_455) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_445), .B(n_449), .C(n_455), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_783), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_733), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_673), .B(n_732), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_465), .B(n_734), .C(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g823 ( .A(n_465), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_637), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_578), .C(n_607), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_468), .B(n_567), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_488), .B1(n_527), .B2(n_539), .Y(n_468) );
NAND2x1_ASAP7_75t_L g769 ( .A(n_469), .B(n_568), .Y(n_769) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
INVx2_ASAP7_75t_L g541 ( .A(n_471), .Y(n_541) );
INVx4_ASAP7_75t_L g583 ( .A(n_471), .Y(n_583) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_471), .Y(n_603) );
AND2x4_ASAP7_75t_L g614 ( .A(n_471), .B(n_582), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_471), .B(n_544), .Y(n_620) );
NOR2x1_ASAP7_75t_SL g693 ( .A(n_471), .B(n_555), .Y(n_693) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVxp67_ASAP7_75t_L g494 ( .A(n_477), .Y(n_494) );
INVx2_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
INVx2_ASAP7_75t_L g586 ( .A(n_480), .Y(n_586) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_480), .Y(n_600) );
INVx1_ASAP7_75t_L g611 ( .A(n_480), .Y(n_611) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_480), .Y(n_623) );
AND2x2_ASAP7_75t_L g655 ( .A(n_480), .B(n_555), .Y(n_655) );
INVx1_ASAP7_75t_L g681 ( .A(n_480), .Y(n_681) );
AND2x2_ASAP7_75t_L g743 ( .A(n_480), .B(n_571), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_507), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g636 ( .A(n_490), .B(n_575), .Y(n_636) );
INVx2_ASAP7_75t_L g678 ( .A(n_490), .Y(n_678) );
AND2x2_ASAP7_75t_L g780 ( .A(n_490), .B(n_507), .Y(n_780) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_491), .B(n_530), .Y(n_574) );
INVx2_ASAP7_75t_L g595 ( .A(n_491), .Y(n_595) );
AND2x4_ASAP7_75t_L g617 ( .A(n_491), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g652 ( .A(n_491), .Y(n_652) );
AND2x2_ASAP7_75t_L g776 ( .A(n_491), .B(n_533), .Y(n_776) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_499), .A2(n_509), .B(n_515), .Y(n_508) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_499), .A2(n_509), .B(n_515), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g750 ( .A(n_507), .Y(n_750) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
NOR2xp67_ASAP7_75t_L g625 ( .A(n_508), .B(n_595), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_508), .B(n_595), .Y(n_630) );
INVx2_ASAP7_75t_L g643 ( .A(n_508), .Y(n_643) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_508), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AND2x4_ASAP7_75t_L g616 ( .A(n_516), .B(n_529), .Y(n_616) );
AND2x2_ASAP7_75t_L g631 ( .A(n_516), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g686 ( .A(n_516), .Y(n_686) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_517), .B(n_533), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_517), .B(n_530), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVxp33_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx3_ASAP7_75t_L g592 ( .A(n_529), .Y(n_592) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
AND2x2_ASAP7_75t_L g704 ( .A(n_530), .B(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g647 ( .A(n_531), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_531), .B(n_686), .Y(n_727) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g594 ( .A(n_532), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g575 ( .A(n_533), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
INVxp67_ASAP7_75t_L g632 ( .A(n_533), .Y(n_632) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_533), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_533), .Y(n_709) );
INVx1_ASAP7_75t_L g687 ( .A(n_539), .Y(n_687) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_540), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g729 ( .A(n_541), .B(n_570), .Y(n_729) );
OR2x2_ASAP7_75t_L g781 ( .A(n_542), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g680 ( .A(n_543), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g716 ( .A(n_543), .B(n_603), .Y(n_716) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x4_ASAP7_75t_L g570 ( .A(n_544), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
INVx2_ASAP7_75t_L g599 ( .A(n_544), .Y(n_599) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_544), .Y(n_725) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVx3_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx2_ASAP7_75t_L g665 ( .A(n_555), .Y(n_665) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_566), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_569), .B(n_645), .Y(n_662) );
NOR2x1_ASAP7_75t_L g754 ( .A(n_569), .B(n_583), .Y(n_754) );
INVx4_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_570), .B(n_645), .Y(n_731) );
AND2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g612 ( .A(n_571), .Y(n_612) );
AOI22xp5_ASAP7_75t_SL g660 ( .A1(n_572), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_573), .B(n_631), .Y(n_657) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g765 ( .A(n_574), .B(n_606), .Y(n_765) );
AND2x2_ASAP7_75t_L g588 ( .A(n_575), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g624 ( .A(n_575), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g767 ( .A(n_575), .B(n_678), .Y(n_767) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g642 ( .A(n_577), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g668 ( .A(n_577), .Y(n_668) );
AND2x2_ASAP7_75t_L g703 ( .A(n_577), .B(n_595), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_587), .B1(n_591), .B2(n_596), .C(n_601), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_581), .B(n_655), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_581), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NOR2xp67_ASAP7_75t_SL g627 ( .A(n_583), .B(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
AND2x4_ASAP7_75t_SL g724 ( .A(n_583), .B(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g771 ( .A(n_583), .B(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g645 ( .A(n_585), .Y(n_645) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_586), .Y(n_782) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221x1_ASAP7_75t_L g735 ( .A1(n_588), .A2(n_736), .B1(n_738), .B2(n_739), .C(n_741), .Y(n_735) );
AND2x2_ASAP7_75t_L g661 ( .A(n_589), .B(n_617), .Y(n_661) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g604 ( .A(n_592), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_592), .B(n_594), .Y(n_778) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_598), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_598), .B(n_611), .Y(n_628) );
INVx2_ASAP7_75t_L g635 ( .A(n_598), .Y(n_635) );
INVx1_ASAP7_75t_L g697 ( .A(n_599), .Y(n_697) );
BUFx2_ASAP7_75t_L g717 ( .A(n_600), .Y(n_717) );
NAND2xp33_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
OR2x6_ASAP7_75t_L g634 ( .A(n_603), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g763 ( .A(n_603), .B(n_655), .Y(n_763) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_626), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_615), .B1(n_619), .B2(n_624), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
AND2x2_ASAP7_75t_SL g672 ( .A(n_610), .B(n_614), .Y(n_672) );
AND2x4_ASAP7_75t_L g738 ( .A(n_610), .B(n_696), .Y(n_738) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_611), .B(n_612), .Y(n_610) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_611), .Y(n_753) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_614), .B(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_614), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_614), .B(n_645), .Y(n_737) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g758 ( .A(n_616), .B(n_677), .Y(n_758) );
INVx3_ASAP7_75t_L g669 ( .A(n_617), .Y(n_669) );
AND2x2_ASAP7_75t_L g690 ( .A(n_617), .B(n_642), .Y(n_690) );
NAND2x1_ASAP7_75t_SL g761 ( .A(n_617), .B(n_668), .Y(n_761) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_633), .B2(n_636), .Y(n_626) );
BUFx2_ASAP7_75t_L g682 ( .A(n_628), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_629), .A2(n_720), .B1(n_729), .B2(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_630), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g650 ( .A(n_631), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_635), .B(n_715), .C(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
AOI211x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_646), .B(n_648), .C(n_666), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_641), .B(n_729), .Y(n_748) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_642), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g720 ( .A(n_642), .B(n_678), .Y(n_720) );
AND2x2_ASAP7_75t_L g775 ( .A(n_642), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g698 ( .A(n_645), .Y(n_698) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g740 ( .A(n_647), .B(n_685), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_660), .Y(n_648) );
AOI22xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B1(n_656), .B2(n_658), .Y(n_649) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g713 ( .A(n_652), .B(n_708), .Y(n_713) );
INVx1_ASAP7_75t_SL g755 ( .A(n_652), .Y(n_755) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_655), .B(n_724), .Y(n_723) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g759 ( .A(n_664), .B(n_681), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B(n_671), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_668), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g683 ( .A(n_669), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_673), .Y(n_825) );
NAND3x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_710), .C(n_718), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g784 ( .A(n_674), .B(n_710), .C(n_718), .D(n_785), .Y(n_784) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_688), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_682), .B2(n_683), .C1(n_685), .C2(n_687), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g762 ( .A1(n_680), .A2(n_763), .B(n_764), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_681), .B(n_696), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_684), .A2(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_699), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_692), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_696), .B(n_698), .Y(n_701) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_706), .B2(n_707), .Y(n_699) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g707 ( .A(n_703), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g744 ( .A(n_713), .Y(n_744) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_728), .Y(n_718) );
AOI22xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_721), .B1(n_723), .B2(n_726), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp33_ASAP7_75t_L g733 ( .A(n_732), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g824 ( .A(n_734), .Y(n_824) );
NAND3x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_746), .C(n_766), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_738), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_757) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g772 ( .A(n_743), .Y(n_772) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_756), .Y(n_746) );
AOI21xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_749), .B(n_755), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_762), .Y(n_756) );
INVx2_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_761), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_770), .B2(n_773), .C(n_777), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_789), .B(n_827), .C(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_796), .Y(n_789) );
INVxp33_ASAP7_75t_L g801 ( .A(n_790), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
CKINVDCx8_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_796), .Y(n_800) );
INVx1_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_800), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_804), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_812), .B(n_826), .Y(n_805) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_815), .B1(n_821), .B2(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AND3x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .C(n_825), .Y(n_822) );
endmodule