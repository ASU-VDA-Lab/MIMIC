module fake_jpeg_27798_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx11_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_12),
.B1(n_18),
.B2(n_15),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_19),
.B1(n_16),
.B2(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_11),
.C(n_14),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_23),
.C(n_10),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_31),
.B(n_2),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_46),
.B(n_1),
.Y(n_52)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_55),
.B1(n_41),
.B2(n_26),
.Y(n_61)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_8),
.C(n_7),
.D(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

OAI22x1_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_30),
.B1(n_10),
.B2(n_14),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.C(n_11),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_30),
.B(n_10),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_63),
.C(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_48),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_4),
.C(n_6),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_48),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_14),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.C(n_1),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_24),
.C(n_20),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_75),
.B(n_2),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_24),
.Y(n_78)
);


endmodule