module fake_netlist_1_12672_n_717 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_717, n_716);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_717;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_SL g107 ( .A(n_91), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_36), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_60), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_106), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_65), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_67), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_71), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_103), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_0), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_9), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_42), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_74), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_75), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_96), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
OR2x2_ASAP7_75t_L g124 ( .A(n_29), .B(n_16), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_32), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_23), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_2), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_34), .Y(n_129) );
INVxp33_ASAP7_75t_SL g130 ( .A(n_27), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_21), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_73), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_35), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_33), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_43), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_50), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_47), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_24), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_6), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_17), .Y(n_140) );
BUFx5_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_54), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_62), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_11), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_53), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_87), .Y(n_146) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_1), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_15), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_78), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_143), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_150), .B(n_1), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_112), .A2(n_51), .B(n_104), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_107), .B(n_2), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_118), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_107), .B(n_3), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_125), .B(n_4), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_122), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_157), .B(n_130), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_171), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_165), .B(n_119), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_157), .B(n_110), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_171), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_171), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_152), .B(n_112), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_165), .B(n_110), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_152), .B(n_144), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_152), .B(n_133), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_170), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_166), .B(n_108), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_154), .A2(n_117), .B1(n_127), .B2(n_148), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_163), .B(n_140), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_158), .B(n_121), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_171), .B(n_133), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_168), .B(n_109), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_195), .A2(n_163), .B1(n_166), .B2(n_146), .Y(n_199) );
AO22x1_ASAP7_75t_L g200 ( .A1(n_193), .A2(n_130), .B1(n_160), .B2(n_151), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_183), .B(n_154), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_190), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_173), .B(n_111), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_193), .A2(n_160), .B1(n_168), .B2(n_169), .Y(n_205) );
BUFx12f_ASAP7_75t_L g206 ( .A(n_195), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_193), .A2(n_168), .B1(n_169), .B2(n_164), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_186), .B(n_111), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_193), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_136), .B(n_115), .C(n_123), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_192), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_193), .B(n_176), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_194), .B(n_132), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_177), .B(n_132), .Y(n_215) );
NOR2xp67_ASAP7_75t_L g216 ( .A(n_185), .B(n_155), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_193), .B(n_151), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_172), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_193), .B(n_155), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_193), .B(n_155), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_198), .B(n_155), .Y(n_222) );
AND2x6_ASAP7_75t_L g223 ( .A(n_174), .B(n_113), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_198), .B(n_162), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_174), .B(n_162), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_195), .B(n_147), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_169), .B(n_164), .C(n_161), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_195), .A2(n_122), .B1(n_146), .B2(n_126), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
AND2x6_ASAP7_75t_SL g230 ( .A(n_185), .B(n_116), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_167), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_180), .B(n_167), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_174), .B(n_162), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_209), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
NOR2x1_ASAP7_75t_L g236 ( .A(n_226), .B(n_126), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_204), .B(n_181), .Y(n_238) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_228), .A2(n_156), .A3(n_158), .B1(n_191), .B2(n_162), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_197), .B(n_191), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_211), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_229), .B(n_181), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_209), .B(n_181), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_213), .A2(n_181), .B(n_187), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_187), .B(n_196), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_233), .A2(n_187), .B(n_188), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_214), .B(n_187), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_203), .A2(n_179), .B(n_188), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_226), .A2(n_114), .B1(n_184), .B2(n_179), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_201), .A2(n_184), .B(n_178), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_223), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_218), .B(n_172), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_201), .B(n_178), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_189), .B(n_182), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
NAND3xp33_ASAP7_75t_SL g260 ( .A(n_212), .B(n_128), .C(n_124), .Y(n_260) );
CKINVDCx8_ASAP7_75t_R g261 ( .A(n_212), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_202), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_206), .A2(n_189), .B1(n_182), .B2(n_164), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_221), .Y(n_264) );
NAND3x1_ASAP7_75t_L g265 ( .A(n_236), .B(n_199), .C(n_230), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_240), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_264), .A2(n_220), .B(n_219), .C(n_224), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_256), .B(n_222), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_257), .A2(n_232), .A3(n_231), .B(n_189), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_250), .A2(n_210), .B(n_216), .C(n_205), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_254), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_217), .B(n_200), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_246), .A2(n_207), .B(n_156), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_250), .A2(n_215), .B(n_156), .C(n_208), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_255), .A2(n_182), .B(n_142), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_247), .A2(n_145), .B(n_129), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_242), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_264), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_248), .A2(n_134), .B(n_149), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_254), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_244), .B(n_223), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_138), .B(n_135), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_251), .A2(n_158), .B(n_120), .Y(n_284) );
INVx5_ASAP7_75t_L g285 ( .A(n_243), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_261), .B(n_206), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_158), .B(n_223), .C(n_137), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_260), .A2(n_223), .B1(n_131), .B2(n_158), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_240), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_273), .A2(n_262), .B(n_252), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_282), .B(n_259), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_275), .A2(n_273), .B(n_283), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_268), .B(n_262), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_284), .A2(n_258), .B(n_249), .Y(n_294) );
AOI21x1_ASAP7_75t_L g295 ( .A1(n_284), .A2(n_237), .B(n_263), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_279), .B(n_239), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_282), .B(n_244), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_289), .A2(n_243), .B(n_245), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_267), .A2(n_243), .B(n_245), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_274), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_266), .B(n_243), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_285), .B(n_238), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_269), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_239), .B(n_238), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_276), .A2(n_234), .B(n_239), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_277), .A2(n_234), .B(n_158), .Y(n_307) );
AND2x6_ASAP7_75t_L g308 ( .A(n_285), .B(n_239), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_265), .A2(n_223), .B1(n_158), .B2(n_7), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_285), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_294), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_300), .B(n_269), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_311), .B(n_281), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_301), .B(n_285), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_311), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_280), .Y(n_318) );
OR2x6_ASAP7_75t_L g319 ( .A(n_296), .B(n_281), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_304), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_304), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_309), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_290), .A2(n_272), .B(n_280), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_271), .Y(n_327) );
BUFx2_ASAP7_75t_SL g328 ( .A(n_308), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_291), .B(n_270), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_308), .B(n_223), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_306), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_307), .A2(n_287), .B(n_288), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
BUFx4f_ASAP7_75t_L g339 ( .A(n_319), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_331), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_335), .B(n_305), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_335), .B(n_292), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_331), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_325), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_332), .B(n_308), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_325), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_332), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_314), .B(n_292), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_305), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_320), .B(n_305), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_321), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_324), .B(n_337), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_337), .A2(n_306), .B(n_295), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_324), .B(n_308), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_337), .B(n_295), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_332), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_336), .B(n_291), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_291), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_332), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_312), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_338), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_329), .A2(n_310), .B1(n_297), .B2(n_303), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_327), .B(n_286), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_312), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_5), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_322), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_323), .B(n_297), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_318), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_338), .B(n_299), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_359), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_382), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_378), .B(n_330), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_378), .B(n_330), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_339), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_351), .B(n_328), .Y(n_389) );
AND2x4_ASAP7_75t_SL g390 ( .A(n_371), .B(n_319), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_351), .B(n_328), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_370), .B(n_327), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_379), .B(n_319), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_351), .B(n_338), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_348), .B(n_338), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_379), .B(n_329), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_348), .B(n_333), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_345), .B(n_319), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_341), .B(n_317), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_348), .B(n_329), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_352), .B(n_329), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_352), .B(n_342), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_373), .B(n_317), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_341), .B(n_326), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_352), .B(n_326), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_342), .B(n_326), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_342), .B(n_316), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_341), .B(n_316), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_359), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_355), .B(n_334), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_344), .B(n_315), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_354), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_373), .B(n_315), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_354), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_345), .B(n_315), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_360), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_360), .B(n_315), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_339), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_367), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_355), .B(n_6), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_339), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_344), .B(n_7), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_355), .B(n_8), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_377), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_362), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_359), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_339), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_357), .B(n_8), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_370), .B(n_9), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_344), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_344), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_357), .B(n_10), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_346), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_357), .B(n_10), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_359), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_377), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_346), .B(n_11), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_363), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_388), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_346), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_414), .B(n_350), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_388), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_390), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_393), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_393), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_441), .A2(n_339), .B(n_359), .C(n_371), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_406), .B(n_350), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_390), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_408), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_350), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_402), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_389), .B(n_363), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_387), .B(n_345), .Y(n_467) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_387), .B(n_345), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_389), .B(n_364), .Y(n_469) );
NOR2xp67_ASAP7_75t_SL g470 ( .A(n_396), .B(n_359), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_391), .B(n_397), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_410), .B(n_358), .Y(n_472) );
NAND2x1_ASAP7_75t_L g473 ( .A(n_427), .B(n_345), .Y(n_473) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_415), .B(n_359), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_392), .A2(n_369), .B1(n_373), .B2(n_375), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_429), .B(n_12), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_402), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_394), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_401), .B(n_347), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_410), .B(n_412), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_401), .B(n_347), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_399), .B(n_375), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_399), .B(n_375), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_412), .B(n_358), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_416), .B(n_358), .Y(n_486) );
NAND2xp67_ASAP7_75t_L g487 ( .A(n_390), .B(n_364), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_391), .B(n_364), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_397), .B(n_347), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_394), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_384), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_416), .B(n_361), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_404), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_401), .B(n_361), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_404), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_443), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_418), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_398), .B(n_361), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_385), .B(n_365), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_420), .B(n_365), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_429), .B(n_12), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_420), .B(n_365), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_438), .B(n_340), .Y(n_505) );
NOR2x1p5_ASAP7_75t_SL g506 ( .A(n_408), .B(n_366), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_422), .B(n_366), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_445), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_433), .B(n_13), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_440), .B(n_369), .C(n_340), .D(n_343), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_385), .B(n_372), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_422), .B(n_372), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_419), .B(n_374), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_430), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_405), .B(n_374), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_438), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_398), .B(n_368), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_405), .B(n_368), .Y(n_519) );
INVxp67_ASAP7_75t_SL g520 ( .A(n_384), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_430), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_403), .B(n_368), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_437), .B(n_356), .Y(n_523) );
BUFx2_ASAP7_75t_SL g524 ( .A(n_427), .Y(n_524) );
NOR2xp67_ASAP7_75t_L g525 ( .A(n_401), .B(n_340), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_403), .B(n_376), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_421), .B(n_376), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_421), .B(n_376), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_437), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_423), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_386), .B(n_376), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_481), .B(n_400), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_530), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_511), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_452), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_456), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_517), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_462), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_463), .B(n_386), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_474), .B(n_431), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_463), .B(n_384), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_455), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_457), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_459), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_471), .B(n_421), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_450), .B(n_421), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_451), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_479), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_527), .B(n_383), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_486), .B(n_409), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_497), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_528), .B(n_447), .Y(n_554) );
AOI21xp33_ASAP7_75t_SL g555 ( .A1(n_460), .A2(n_431), .B(n_439), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_519), .B(n_447), .Y(n_556) );
NAND2x1_ASAP7_75t_L g557 ( .A(n_470), .B(n_439), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_476), .B(n_395), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_490), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_502), .B(n_395), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_522), .B(n_526), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_486), .B(n_409), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_472), .B(n_409), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_472), .B(n_411), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_509), .B(n_423), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_485), .B(n_407), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_465), .B(n_440), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_495), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_510), .B(n_433), .C(n_446), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_485), .B(n_411), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_453), .B(n_411), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_461), .B(n_424), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_477), .B(n_444), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_489), .B(n_444), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_454), .B(n_424), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_499), .B(n_446), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_492), .B(n_432), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_498), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_464), .B(n_424), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_510), .A2(n_449), .B1(n_343), .B2(n_340), .Y(n_582) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_475), .B(n_449), .C(n_432), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_514), .B(n_434), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_475), .A2(n_343), .B1(n_380), .B2(n_376), .Y(n_585) );
INVxp33_ASAP7_75t_L g586 ( .A(n_467), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_466), .B(n_381), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_525), .B(n_343), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_521), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_469), .B(n_381), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_492), .B(n_14), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_515), .B(n_434), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_381), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_529), .B(n_434), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_513), .B(n_14), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_458), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_500), .Y(n_597) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_480), .B(n_381), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_483), .B(n_435), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_523), .B(n_435), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_518), .B(n_381), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_523), .B(n_435), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_480), .B(n_380), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_524), .Y(n_605) );
AOI32xp33_ASAP7_75t_L g606 ( .A1(n_605), .A2(n_482), .A3(n_494), .B1(n_487), .B2(n_505), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_484), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_570), .A2(n_482), .B1(n_494), .B2(n_468), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_547), .B(n_473), .Y(n_609) );
OAI211xp5_ASAP7_75t_SL g610 ( .A1(n_605), .A2(n_501), .B(n_504), .C(n_531), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_600), .Y(n_611) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_540), .B(n_503), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_596), .B(n_504), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_546), .B(n_491), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g615 ( .A1(n_586), .A2(n_520), .A3(n_516), .B1(n_508), .B2(n_506), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_532), .B(n_520), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_533), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_535), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_538), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_541), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_542), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_543), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
AOI211xp5_ASAP7_75t_SL g624 ( .A1(n_595), .A2(n_507), .B(n_512), .C(n_380), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_550), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_591), .A2(n_507), .B(n_512), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_555), .B(n_436), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_583), .A2(n_380), .B1(n_448), .B2(n_436), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_539), .B(n_436), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_559), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_548), .B(n_562), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_536), .B(n_15), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_582), .B(n_448), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_549), .A2(n_448), .B(n_428), .C(n_426), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_566), .B(n_380), .C(n_426), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_537), .Y(n_637) );
AOI21xp33_ASAP7_75t_L g638 ( .A1(n_558), .A2(n_16), .B(n_17), .Y(n_638) );
INVxp67_ASAP7_75t_L g639 ( .A(n_597), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_569), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_560), .A2(n_428), .B1(n_425), .B2(n_297), .C(n_356), .Y(n_641) );
OAI32xp33_ASAP7_75t_L g642 ( .A1(n_567), .A2(n_425), .A3(n_19), .B1(n_18), .B2(n_356), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_585), .A2(n_425), .B1(n_298), .B2(n_18), .C(n_19), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_557), .A2(n_356), .B1(n_22), .B2(n_25), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_539), .B(n_356), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_592), .A2(n_20), .A3(n_26), .B1(n_28), .B2(n_30), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_580), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_534), .B(n_105), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_552), .B(n_31), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_589), .Y(n_652) );
OAI322xp33_ASAP7_75t_SL g653 ( .A1(n_552), .A2(n_37), .A3(n_38), .B1(n_39), .B2(n_40), .C1(n_41), .C2(n_44), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_632), .A2(n_541), .B(n_598), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_626), .A2(n_563), .B1(n_568), .B2(n_575), .C(n_579), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_613), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_619), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_606), .B(n_588), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_624), .A2(n_577), .B(n_573), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_638), .A2(n_603), .B(n_601), .C(n_564), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_620), .B(n_563), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_619), .B(n_564), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g663 ( .A1(n_624), .A2(n_604), .B(n_578), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_615), .A2(n_565), .B1(n_577), .B2(n_573), .C(n_576), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_608), .A2(n_565), .B(n_603), .C(n_601), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_627), .B(n_604), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_611), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_610), .A2(n_590), .B1(n_593), .B2(n_587), .C(n_584), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_639), .B(n_544), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_653), .A2(n_594), .B(n_584), .Y(n_671) );
OAI32xp33_ASAP7_75t_L g672 ( .A1(n_616), .A2(n_581), .A3(n_599), .B1(n_556), .B2(n_551), .Y(n_672) );
AOI221xp5_ASAP7_75t_SL g673 ( .A1(n_634), .A2(n_554), .B1(n_602), .B2(n_594), .C(n_553), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_612), .A2(n_45), .B(n_46), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_638), .A2(n_48), .B1(n_49), .B2(n_52), .C(n_55), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_641), .A2(n_56), .B1(n_57), .B2(n_58), .C1(n_61), .C2(n_64), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_646), .A2(n_66), .B1(n_68), .B2(n_69), .C(n_70), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_628), .A2(n_72), .B1(n_76), .B2(n_77), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_609), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_645), .B(n_82), .Y(n_680) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_645), .A2(n_83), .B(n_85), .Y(n_681) );
NAND4xp75_ASAP7_75t_L g682 ( .A(n_650), .B(n_614), .C(n_617), .D(n_652), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_635), .A2(n_88), .B(n_89), .Y(n_683) );
NAND2xp67_ASAP7_75t_SL g684 ( .A(n_631), .B(n_92), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_621), .B(n_93), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_637), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_637), .A2(n_94), .B1(n_95), .B2(n_97), .Y(n_687) );
OAI322xp33_ASAP7_75t_SL g688 ( .A1(n_647), .A2(n_98), .A3(n_99), .B1(n_100), .B2(n_101), .C1(n_102), .C2(n_633), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_643), .A2(n_636), .B(n_642), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_651), .B(n_630), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_622), .B(n_623), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_625), .A2(n_640), .B1(n_644), .B2(n_649), .C(n_629), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_607), .A2(n_606), .B(n_624), .C(n_615), .Y(n_693) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_681), .B(n_675), .C(n_693), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_658), .A2(n_663), .B1(n_664), .B2(n_657), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_675), .B(n_689), .C(n_660), .Y(n_696) );
NOR3x1_ASAP7_75t_L g697 ( .A(n_682), .B(n_659), .C(n_666), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_676), .B(n_673), .C(n_671), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_687), .B(n_679), .C(n_665), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_692), .B(n_655), .Y(n_700) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_694), .B(n_684), .Y(n_701) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_695), .B(n_662), .Y(n_702) );
AND4x1_ASAP7_75t_L g703 ( .A(n_698), .B(n_674), .C(n_690), .D(n_683), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_700), .B(n_680), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_701), .B(n_696), .C(n_699), .Y(n_705) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_702), .B(n_697), .C(n_654), .D(n_677), .Y(n_706) );
XNOR2xp5_ASAP7_75t_L g707 ( .A(n_703), .B(n_686), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_705), .B(n_704), .C(n_685), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_707), .B(n_669), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_708), .A2(n_706), .B1(n_656), .B2(n_670), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_709), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_711), .B(n_668), .C(n_667), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_710), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_672), .B(n_688), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_712), .B1(n_661), .B2(n_678), .Y(n_715) );
UNKNOWN g716 ( );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_691), .B(n_648), .Y(n_717) );
endmodule