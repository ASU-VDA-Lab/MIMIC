module fake_jpeg_16496_n_45 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_5),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_16),
.A2(n_24),
.B1(n_8),
.B2(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_12),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_14),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_3),
.C(n_4),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_13),
.C(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_7),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_10),
.B(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_32),
.B1(n_19),
.B2(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_22),
.C(n_30),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_16),
.B(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.C(n_39),
.Y(n_41)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_33),
.B(n_28),
.C(n_25),
.D(n_26),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_37),
.C(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_26),
.A3(n_35),
.B1(n_38),
.B2(n_42),
.C1(n_41),
.C2(n_37),
.Y(n_44)
);


endmodule