module fake_jpeg_8076_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_30),
.B1(n_22),
.B2(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_49),
.B(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_32),
.B1(n_24),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_71),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_24),
.B1(n_40),
.B2(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_41),
.B1(n_37),
.B2(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_65),
.B1(n_72),
.B2(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_35),
.B1(n_34),
.B2(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_41),
.B1(n_45),
.B2(n_36),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_25),
.Y(n_87)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_34),
.B1(n_17),
.B2(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_31),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_85),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_20),
.Y(n_82)
);

NOR2x1_ASAP7_75t_SL g140 ( 
.A(n_82),
.B(n_102),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_96),
.B1(n_70),
.B2(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_87),
.B(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_93),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_41),
.B1(n_38),
.B2(n_45),
.Y(n_89)
);

OAI22x1_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_70),
.B1(n_61),
.B2(n_67),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_41),
.C(n_25),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_63),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_12),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_33),
.B1(n_18),
.B2(n_63),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_100),
.Y(n_129)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NOR4xp25_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_11),
.C(n_16),
.D(n_15),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_123),
.B1(n_128),
.B2(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_127),
.B1(n_113),
.B2(n_85),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_134),
.B(n_18),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_67),
.B1(n_27),
.B2(n_21),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_21),
.B1(n_17),
.B2(n_33),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_100),
.B1(n_109),
.B2(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_83),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_146),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_165),
.B1(n_172),
.B2(n_167),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_111),
.B(n_81),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_149),
.B(n_155),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_90),
.C(n_103),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_151),
.C(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_150),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_111),
.B(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_76),
.C(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_153),
.B1(n_113),
.B2(n_121),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_116),
.B(n_87),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_157),
.B(n_158),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_102),
.B(n_86),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_86),
.B(n_98),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_2),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_4),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_97),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_161),
.B1(n_75),
.B2(n_3),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_107),
.B(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_107),
.B1(n_88),
.B2(n_33),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_79),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_186),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_191),
.C(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_134),
.B1(n_125),
.B2(n_130),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_185),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_125),
.B1(n_128),
.B2(n_126),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_161),
.A3(n_173),
.B1(n_154),
.B2(n_162),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_120),
.B1(n_133),
.B2(n_119),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_170),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_119),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_133),
.B1(n_138),
.B2(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_18),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_124),
.B1(n_59),
.B2(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_79),
.C(n_124),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_203),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_141),
.A2(n_124),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_201),
.B(n_164),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_10),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2x1_ASAP7_75t_R g201 ( 
.A(n_170),
.B(n_10),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_75),
.C(n_3),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_217),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_214),
.B(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_157),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_222),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_155),
.B(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_162),
.B1(n_155),
.B2(n_164),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_154),
.B(n_148),
.C(n_159),
.D(n_161),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_15),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_191),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_226),
.B1(n_190),
.B2(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_204),
.Y(n_243)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_5),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_233),
.B(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_218),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_249),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_178),
.B1(n_186),
.B2(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_250),
.B1(n_228),
.B2(n_216),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_176),
.C(n_196),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_247),
.C(n_255),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_198),
.CI(n_185),
.CON(n_241),
.SN(n_241)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_232),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_179),
.B1(n_204),
.B2(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_197),
.B(n_195),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_214),
.B(n_221),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_206),
.A3(n_182),
.B1(n_205),
.B2(n_203),
.C1(n_14),
.C2(n_7),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_206),
.C(n_9),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_15),
.C(n_16),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_242),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_210),
.B(n_221),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_262),
.B(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_209),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_209),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_269),
.B(n_274),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_215),
.C(n_224),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_215),
.C(n_237),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_226),
.B(n_208),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_241),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_228),
.B1(n_231),
.B2(n_220),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_250),
.B1(n_254),
.B2(n_240),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_286),
.C(n_257),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_249),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_245),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_288),
.B(n_289),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_262),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_251),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_256),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_270),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_295),
.C(n_297),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_260),
.B(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_294),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_235),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_217),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_260),
.C(n_265),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_264),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_257),
.C(n_258),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_259),
.B1(n_277),
.B2(n_269),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_313),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_259),
.B1(n_282),
.B2(n_272),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_293),
.B(n_223),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_281),
.B1(n_279),
.B2(n_274),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_311),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_283),
.B(n_261),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_252),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_263),
.B1(n_273),
.B2(n_241),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_273),
.B1(n_286),
.B2(n_252),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_300),
.B(n_295),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_319),
.A3(n_320),
.B1(n_305),
.B2(n_311),
.C1(n_313),
.C2(n_304),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_219),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_219),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_291),
.B(n_255),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_323),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_247),
.CI(n_219),
.CON(n_323),
.SN(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_325),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_323),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_314),
.Y(n_329)
);


endmodule