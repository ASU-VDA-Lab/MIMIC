module fake_jpeg_18211_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_19),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_21),
.B(n_1),
.Y(n_25)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_1),
.B1(n_6),
.B2(n_9),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_17),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_7),
.B(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_33),
.B(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_11),
.B1(n_16),
.B2(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_1),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_14),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_34),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_37),
.B(n_36),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_45),
.B(n_38),
.Y(n_48)
);


endmodule