module fake_jpeg_3188_n_637 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_637);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_637;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_60),
.B(n_75),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_18),
.C(n_1),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_61),
.B(n_12),
.C(n_13),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_71),
.Y(n_153)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_72),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_73),
.Y(n_192)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_15),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_78),
.B(n_119),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_79),
.B(n_82),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_80),
.Y(n_212)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_0),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_91),
.Y(n_132)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_88),
.A2(n_112),
.B1(n_25),
.B2(n_41),
.Y(n_193)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_90),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_22),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_107),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_102),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_105),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx11_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_3),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_3),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_29),
.Y(n_150)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_26),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_113),
.Y(n_225)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_21),
.B(n_4),
.Y(n_119)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_21),
.B(n_15),
.CON(n_121),
.SN(n_121)
);

HAxp5_ASAP7_75t_SL g221 ( 
.A(n_121),
.B(n_126),
.CON(n_221),
.SN(n_221)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_26),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_122),
.A2(n_34),
.B1(n_37),
.B2(n_128),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_123),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_20),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_128),
.Y(n_184)
);

HAxp5_ASAP7_75t_SL g126 ( 
.A(n_27),
.B(n_5),
.CON(n_126),
.SN(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_31),
.Y(n_127)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_130),
.Y(n_194)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_53),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_51),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_139),
.B(n_141),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_51),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_33),
.B1(n_55),
.B2(n_53),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g263 ( 
.A1(n_142),
.A2(n_212),
.B1(n_175),
.B2(n_219),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_150),
.B(n_152),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_66),
.B(n_47),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_77),
.B(n_55),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_SL g261 ( 
.A(n_156),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_77),
.B(n_47),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_157),
.B(n_164),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_63),
.A2(n_37),
.B1(n_55),
.B2(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_161),
.A2(n_193),
.B1(n_215),
.B2(n_14),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_163),
.A2(n_197),
.B1(n_202),
.B2(n_227),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_29),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_85),
.B(n_28),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_166),
.B(n_167),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_70),
.B(n_28),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_106),
.B(n_50),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_171),
.B(n_172),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_27),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_50),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_181),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_102),
.A2(n_55),
.B1(n_53),
.B2(n_37),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_215),
.B1(n_211),
.B2(n_180),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_44),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_214),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_25),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_182),
.B(n_191),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_64),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_123),
.A2(n_42),
.B1(n_57),
.B2(n_34),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_118),
.B(n_20),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_198),
.B(n_203),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_199),
.B(n_201),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_118),
.B(n_20),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_125),
.A2(n_25),
.B1(n_41),
.B2(n_38),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_41),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_59),
.B(n_57),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_204),
.B(n_207),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_74),
.B(n_110),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_89),
.B(n_38),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_100),
.B(n_38),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_131),
.B(n_34),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_37),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_216),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_69),
.B(n_15),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_217),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_126),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_83),
.B1(n_90),
.B2(n_95),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_108),
.B(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_212),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_73),
.B(n_12),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_226),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_111),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_141),
.A2(n_84),
.B1(n_97),
.B2(n_80),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_233),
.B(n_302),
.Y(n_328)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_154),
.Y(n_236)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_238),
.A2(n_303),
.B1(n_306),
.B2(n_178),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_132),
.A2(n_113),
.B1(n_12),
.B2(n_14),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_242),
.A2(n_277),
.B1(n_288),
.B2(n_295),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_246),
.Y(n_353)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_249),
.A2(n_251),
.B1(n_257),
.B2(n_262),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_161),
.B1(n_222),
.B2(n_142),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_250),
.A2(n_233),
.B1(n_249),
.B2(n_232),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_169),
.A2(n_134),
.B1(n_195),
.B2(n_139),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_252),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_218),
.B(n_142),
.C(n_156),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_148),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_255),
.B(n_260),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_186),
.B1(n_142),
.B2(n_211),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g258 ( 
.A(n_146),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_258),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_170),
.A2(n_221),
.B1(n_229),
.B2(n_136),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_263),
.A2(n_269),
.B1(n_317),
.B2(n_253),
.Y(n_372)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_149),
.A2(n_156),
.B(n_184),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_267),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_136),
.A2(n_162),
.B1(n_138),
.B2(n_143),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_149),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_270),
.B(n_273),
.Y(n_336)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_149),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_190),
.A2(n_184),
.B1(n_147),
.B2(n_135),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_190),
.A2(n_184),
.B1(n_147),
.B2(n_174),
.Y(n_277)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g340 ( 
.A(n_278),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_282),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_153),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_283),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_175),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_286),
.B(n_287),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_145),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_135),
.A2(n_174),
.B1(n_224),
.B2(n_185),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_162),
.A2(n_188),
.B(n_165),
.C(n_140),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_290),
.B(n_291),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_145),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_165),
.B(n_188),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_224),
.A2(n_223),
.B1(n_133),
.B2(n_189),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_159),
.Y(n_296)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_159),
.B(n_179),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_133),
.Y(n_299)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_299),
.Y(n_375)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_179),
.Y(n_300)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_196),
.A2(n_225),
.B1(n_205),
.B2(n_189),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_158),
.A2(n_196),
.B1(n_205),
.B2(n_225),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_158),
.B(n_143),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_153),
.Y(n_305)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_155),
.A2(n_200),
.B1(n_137),
.B2(n_220),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_208),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_318),
.Y(n_362)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_309),
.Y(n_335)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_137),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_192),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_310),
.B(n_260),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_213),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_266),
.C(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_168),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_313),
.B(n_314),
.Y(n_351)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_151),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_316),
.Y(n_352)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_160),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_178),
.A2(n_220),
.B1(n_219),
.B2(n_173),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_213),
.A2(n_168),
.B(n_200),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_325),
.B(n_345),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_333),
.A2(n_373),
.B1(n_244),
.B2(n_237),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_289),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_261),
.B(n_151),
.C(n_173),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_350),
.C(n_265),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_259),
.B(n_173),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_347),
.B(n_365),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_261),
.B(n_259),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_256),
.B(n_268),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_355),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_246),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_379),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_292),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_364),
.A2(n_371),
.B(n_305),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_247),
.B(n_240),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_240),
.B(n_285),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_369),
.B(n_280),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_370),
.A2(n_250),
.B1(n_263),
.B2(n_319),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_276),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_290),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_270),
.A2(n_273),
.B1(n_263),
.B2(n_248),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_271),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_265),
.B(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_336),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_409),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_323),
.A2(n_319),
.B1(n_271),
.B2(n_298),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_384),
.A2(n_376),
.B(n_338),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_385),
.B(n_331),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_320),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_387),
.A2(n_328),
.B1(n_333),
.B2(n_321),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_346),
.C(n_359),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_416),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_390),
.B(n_414),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_362),
.A2(n_301),
.B(n_254),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_392),
.A2(n_400),
.B(n_419),
.Y(n_433)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_364),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_394),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_362),
.A2(n_318),
.B(n_234),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_363),
.B(n_366),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_372),
.A2(n_302),
.B1(n_304),
.B2(n_297),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_397),
.A2(n_402),
.B1(n_404),
.B2(n_410),
.Y(n_450)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_324),
.A2(n_236),
.B(n_235),
.Y(n_400)
);

OR2x2_ASAP7_75t_SL g401 ( 
.A(n_327),
.B(n_324),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_413),
.C(n_423),
.Y(n_427)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_326),
.Y(n_403)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_370),
.A2(n_253),
.B1(n_294),
.B2(n_314),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_405),
.Y(n_448)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_407),
.Y(n_465)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_349),
.A2(n_241),
.B1(n_245),
.B2(n_300),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_417),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_354),
.A2(n_316),
.B1(n_296),
.B2(n_299),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_412),
.A2(n_418),
.B1(n_424),
.B2(n_426),
.Y(n_453)
);

OR2x2_ASAP7_75t_SL g413 ( 
.A(n_327),
.B(n_258),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_275),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_SL g415 ( 
.A(n_380),
.B(n_313),
.C(n_307),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_415),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_354),
.A2(n_264),
.B1(n_308),
.B2(n_281),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_343),
.A2(n_309),
.B(n_282),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_284),
.C(n_252),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_352),
.Y(n_438)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_358),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g423 ( 
.A1(n_347),
.A2(n_278),
.B(n_272),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_366),
.A2(n_243),
.B1(n_279),
.B2(n_315),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_425),
.B(n_341),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_329),
.A2(n_328),
.B1(n_320),
.B2(n_323),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_428),
.A2(n_458),
.B(n_384),
.Y(n_489)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_442),
.C(n_446),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_451),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_385),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_401),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_334),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_395),
.A2(n_328),
.B(n_342),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_400),
.B(n_419),
.Y(n_474)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_386),
.B(n_329),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_334),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_459),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_391),
.B(n_365),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_462),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_402),
.B(n_332),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_332),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_463),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_369),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_461),
.B(n_351),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_420),
.B(n_331),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_396),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_464),
.A2(n_381),
.B1(n_399),
.B2(n_393),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_325),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_390),
.B(n_335),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_361),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_436),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_468),
.B(n_432),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_435),
.B(n_392),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_472),
.B(n_475),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_474),
.A2(n_483),
.B(n_489),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_426),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_463),
.A2(n_387),
.B1(n_418),
.B2(n_412),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_477),
.A2(n_495),
.B1(n_497),
.B2(n_498),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_500),
.C(n_432),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_344),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_479),
.B(n_361),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_421),
.C(n_404),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_438),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_428),
.A2(n_397),
.B(n_413),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_434),
.Y(n_484)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_487),
.Y(n_525)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_382),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_493),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_494),
.B(n_496),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_450),
.B1(n_453),
.B2(n_440),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_450),
.A2(n_405),
.B1(n_406),
.B2(n_403),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_453),
.A2(n_422),
.B1(n_425),
.B2(n_409),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_504),
.B1(n_455),
.B2(n_448),
.Y(n_519)
);

NAND4xp25_ASAP7_75t_SL g501 ( 
.A(n_459),
.B(n_376),
.C(n_340),
.D(n_357),
.Y(n_501)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_501),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_407),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_445),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_454),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_445),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_497),
.A2(n_447),
.B1(n_460),
.B2(n_456),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_506),
.A2(n_512),
.B1(n_536),
.B2(n_486),
.Y(n_562)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_509),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_511),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_496),
.A2(n_456),
.B1(n_427),
.B2(n_433),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_457),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_514),
.B(n_515),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_516),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_498),
.A2(n_451),
.B1(n_441),
.B2(n_433),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_517),
.A2(n_527),
.B1(n_495),
.B2(n_473),
.Y(n_543)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_519),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_487),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_520),
.B(n_523),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_489),
.A2(n_462),
.B(n_452),
.Y(n_522)
);

OAI21x1_ASAP7_75t_SL g542 ( 
.A1(n_522),
.A2(n_480),
.B(n_474),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_526),
.B(n_476),
.C(n_521),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_483),
.A2(n_444),
.B1(n_455),
.B2(n_448),
.Y(n_527)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_529),
.Y(n_539)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_530),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_411),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_532),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_534),
.B(n_502),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_480),
.A2(n_429),
.B1(n_465),
.B2(n_430),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_472),
.B(n_465),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_476),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_540),
.B(n_554),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_542),
.A2(n_524),
.B(n_531),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_543),
.B(n_545),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_516),
.A2(n_471),
.B1(n_470),
.B2(n_473),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_544),
.A2(n_551),
.B1(n_564),
.B2(n_565),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_475),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_549),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_510),
.A2(n_471),
.B1(n_499),
.B2(n_470),
.Y(n_551)
);

FAx1_ASAP7_75t_SL g552 ( 
.A(n_527),
.B(n_482),
.CI(n_504),
.CON(n_552),
.SN(n_552)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_536),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_492),
.Y(n_553)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_553),
.Y(n_586)
);

XNOR2x1_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_512),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_556),
.B(n_559),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_505),
.C(n_494),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_518),
.C(n_522),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_485),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_534),
.B(n_484),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_368),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_562),
.A2(n_517),
.B1(n_507),
.B2(n_508),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_525),
.B(n_491),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_563),
.B(n_368),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_506),
.A2(n_490),
.B1(n_430),
.B2(n_431),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_523),
.A2(n_501),
.B1(n_358),
.B2(n_356),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_567),
.A2(n_357),
.B1(n_339),
.B2(n_377),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_547),
.B(n_509),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_568),
.B(n_571),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_546),
.A2(n_507),
.B1(n_538),
.B2(n_535),
.Y(n_572)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_573),
.A2(n_577),
.B(n_552),
.Y(n_599)
);

NAND4xp25_ASAP7_75t_L g574 ( 
.A(n_543),
.B(n_529),
.C(n_513),
.D(n_528),
.Y(n_574)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_574),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_SL g575 ( 
.A1(n_563),
.A2(n_524),
.B(n_544),
.C(n_560),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_584),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_541),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_576),
.A2(n_557),
.B1(n_539),
.B2(n_565),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_531),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_583),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_545),
.B(n_528),
.C(n_367),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_580),
.B(n_585),
.C(n_587),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_560),
.A2(n_356),
.B1(n_408),
.B2(n_341),
.Y(n_582)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_582),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_540),
.B(n_374),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_339),
.C(n_377),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_573),
.A2(n_555),
.B(n_554),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_588),
.A2(n_604),
.B1(n_595),
.B2(n_590),
.Y(n_615)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_553),
.Y(n_594)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_549),
.C(n_561),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_600),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_570),
.A2(n_551),
.B1(n_564),
.B2(n_559),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_598),
.A2(n_567),
.B1(n_575),
.B2(n_566),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_602),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_550),
.C(n_557),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_552),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_601),
.B(n_566),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_571),
.A2(n_348),
.B(n_353),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_608),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_589),
.B(n_569),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_609),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_593),
.B(n_578),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_600),
.B(n_580),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_610),
.B(n_616),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_569),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_615),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_578),
.C(n_583),
.Y(n_616)
);

AOI322xp5_ASAP7_75t_L g618 ( 
.A1(n_614),
.A2(n_595),
.A3(n_594),
.B1(n_603),
.B2(n_601),
.C1(n_599),
.C2(n_590),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_618),
.B(n_623),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_612),
.A2(n_598),
.B1(n_588),
.B2(n_596),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_622),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_616),
.B(n_592),
.C(n_596),
.Y(n_622)
);

AOI322xp5_ASAP7_75t_L g623 ( 
.A1(n_605),
.A2(n_575),
.A3(n_602),
.B1(n_604),
.B2(n_585),
.C1(n_592),
.C2(n_353),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_617),
.A2(n_624),
.B(n_607),
.Y(n_625)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_625),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_619),
.A2(n_613),
.B(n_606),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_628),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_622),
.A2(n_611),
.B(n_613),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_627),
.B(n_621),
.C(n_620),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_629),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_633),
.B(n_634),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_632),
.A2(n_621),
.B(n_609),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_630),
.B(n_575),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_636),
.B(n_348),
.Y(n_637)
);


endmodule