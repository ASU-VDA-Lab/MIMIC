module fake_aes_5650_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
AND2x2_ASAP7_75t_SL g4 ( .A(n_0), .B(n_2), .Y(n_4) );
AND2x4_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
AOI22xp33_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
AOI21xp33_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_6), .B(n_5), .Y(n_8) );
O2A1O1Ixp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_7), .B(n_5), .C(n_2), .Y(n_9) );
OR5x1_ASAP7_75t_L g10 ( .A(n_9), .B(n_1), .C(n_5), .D(n_4), .E(n_2), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
endmodule