module fake_netlist_1_6558_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
AOI22xp33_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_5) );
O2A1O1Ixp33_ASAP7_75t_SL g6 ( .A1(n_3), .A2(n_4), .B(n_1), .C(n_0), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_0), .Y(n_8) );
NAND4xp25_ASAP7_75t_L g9 ( .A(n_8), .B(n_1), .C(n_2), .D(n_7), .Y(n_9) );
NAND2x1p5_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_1), .B1(n_2), .B2(n_7), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
endmodule