module real_jpeg_8324_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_2),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_2),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_25),
.B(n_58),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_79),
.B1(n_92),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_2),
.A2(n_32),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_32),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_2),
.A2(n_44),
.B1(n_84),
.B2(n_145),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_9),
.A2(n_25),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_9),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_11),
.A2(n_36),
.B1(n_92),
.B2(n_115),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_12),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_25),
.B1(n_37),
.B2(n_70),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_70),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_15),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_74),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_86),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_19),
.B(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_63),
.C(n_75),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_20),
.A2(n_21),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_41),
.B1(n_42),
.B2(n_62),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_38),
.B1(n_40),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_24),
.A2(n_30),
.B1(n_35),
.B2(n_78),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_79),
.CON(n_78),
.SN(n_78)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_27),
.B(n_32),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_29),
.A2(n_31),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_32),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_65),
.Y(n_66)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_40),
.B(n_79),
.Y(n_156)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_51),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_46),
.B1(n_84),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_44),
.A2(n_84),
.B1(n_127),
.B2(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_44),
.B(n_79),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_45),
.A2(n_54),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_45),
.B(n_83),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_48),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_47),
.B(n_68),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_47),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_48),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_60),
.C(n_62),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_59),
.B(n_92),
.C(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_79),
.B(n_91),
.C(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_63),
.A2(n_75),
.B1(n_76),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_63),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B(n_71),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_64),
.A2(n_67),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_64),
.A2(n_67),
.B1(n_135),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_158),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_67),
.B(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_77),
.B(n_81),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_129),
.B(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_100),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_173),
.B(n_179),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_162),
.B(n_172),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_152),
.B(n_161),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_141),
.B(n_151),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_130),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_140),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_146),
.B(n_150),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_155),
.B(n_163),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.CI(n_159),
.CON(n_155),
.SN(n_155)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_166),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);


endmodule