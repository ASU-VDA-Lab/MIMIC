module real_aes_6538_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_156;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_0), .A2(n_177), .B(n_552), .C(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_1), .B(n_502), .Y(n_556) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g189 ( .A(n_3), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_4), .B(n_149), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_5), .A2(n_475), .B(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_6), .A2(n_169), .B(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_7), .A2(n_38), .B1(n_143), .B2(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_8), .B(n_169), .Y(n_178) );
AND2x6_ASAP7_75t_L g161 ( .A(n_9), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_10), .A2(n_161), .B(n_480), .C(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_11), .B(n_39), .Y(n_437) );
INVx1_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
INVx1_ASAP7_75t_L g182 ( .A(n_13), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_14), .B(n_147), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_15), .B(n_149), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_16), .B(n_135), .Y(n_253) );
AO32x2_ASAP7_75t_L g195 ( .A1(n_17), .A2(n_134), .A3(n_160), .B1(n_169), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_18), .B(n_143), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_19), .B(n_135), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_20), .A2(n_54), .B1(n_143), .B2(n_198), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_21), .A2(n_81), .B1(n_143), .B2(n_147), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_22), .B(n_143), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_23), .A2(n_160), .B(n_480), .C(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_24), .A2(n_60), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_24), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_25), .A2(n_160), .B(n_480), .C(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_26), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_27), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_28), .B(n_442), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_29), .A2(n_475), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_30), .B(n_164), .Y(n_212) );
INVx2_ASAP7_75t_L g145 ( .A(n_31), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_32), .A2(n_478), .B(n_488), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_33), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_34), .B(n_164), .Y(n_223) );
XNOR2x2_ASAP7_75t_SL g122 ( .A(n_35), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_36), .B(n_219), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_37), .A2(n_85), .B1(n_457), .B2(n_458), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_37), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_40), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_41), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_42), .B(n_149), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_43), .B(n_475), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_44), .A2(n_478), .B(n_482), .C(n_488), .Y(n_477) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_45), .A2(n_122), .A3(n_431), .B1(n_438), .B2(n_439), .C(n_441), .Y(n_121) );
INVx1_ASAP7_75t_L g438 ( .A(n_45), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_46), .B(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g553 ( .A(n_47), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_48), .A2(n_91), .B1(n_198), .B2(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g483 ( .A(n_49), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_50), .B(n_143), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_51), .B(n_143), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_52), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_53), .B(n_155), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_55), .A2(n_61), .B1(n_143), .B2(n_147), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_56), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_57), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_58), .B(n_143), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_59), .B(n_143), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_60), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_60), .A2(n_126), .B1(n_127), .B2(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g162 ( .A(n_62), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_63), .B(n_475), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_64), .B(n_502), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_65), .A2(n_155), .B(n_185), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_66), .B(n_143), .Y(n_190) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_68), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_69), .B(n_149), .Y(n_520) );
AO32x2_ASAP7_75t_L g233 ( .A1(n_70), .A2(n_160), .A3(n_169), .B1(n_234), .B2(n_238), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_71), .B(n_150), .Y(n_566) );
INVx1_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
INVx1_ASAP7_75t_L g207 ( .A(n_73), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_74), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_75), .B(n_485), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_76), .A2(n_480), .B(n_488), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_77), .B(n_147), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_78), .Y(n_497) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_80), .B(n_484), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_82), .B(n_198), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_83), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_84), .B(n_147), .Y(n_211) );
INVx1_ASAP7_75t_L g458 ( .A(n_85), .Y(n_458) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_87), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_88), .B(n_159), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_89), .B(n_147), .Y(n_173) );
INVx2_ASAP7_75t_L g114 ( .A(n_90), .Y(n_114) );
OR2x2_ASAP7_75t_L g434 ( .A(n_90), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g462 ( .A(n_90), .B(n_436), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_92), .A2(n_103), .B1(n_147), .B2(n_148), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_93), .B(n_475), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_94), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_95), .A2(n_105), .B1(n_118), .B2(n_771), .Y(n_104) );
INVxp67_ASAP7_75t_L g500 ( .A(n_96), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_97), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_98), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g541 ( .A(n_99), .Y(n_541) );
INVx1_ASAP7_75t_L g562 ( .A(n_100), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_101), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_101), .Y(n_454) );
AND2x2_ASAP7_75t_L g490 ( .A(n_102), .B(n_164), .Y(n_490) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g772 ( .A(n_106), .Y(n_772) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g436 ( .A(n_113), .B(n_437), .Y(n_436) );
NOR2x2_ASAP7_75t_L g450 ( .A(n_114), .B(n_435), .Y(n_450) );
OR2x2_ASAP7_75t_L g467 ( .A(n_114), .B(n_436), .Y(n_467) );
OA211x2_ASAP7_75t_L g118 ( .A1(n_115), .A2(n_119), .B(n_121), .C(n_445), .Y(n_118) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g446 ( .A(n_120), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_122), .B(n_440), .Y(n_439) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx1_ASAP7_75t_SL g464 ( .A(n_127), .Y(n_464) );
OR3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_359), .C(n_408), .Y(n_127) );
NAND5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_274), .C(n_302), .D(n_332), .E(n_346), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_192), .B1(n_224), .B2(n_229), .C(n_240), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_131), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g254 ( .A(n_132), .Y(n_254) );
AND2x2_ASAP7_75t_L g262 ( .A(n_132), .B(n_168), .Y(n_262) );
AND2x2_ASAP7_75t_L g285 ( .A(n_132), .B(n_167), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_132), .B(n_179), .Y(n_300) );
OR2x2_ASAP7_75t_L g309 ( .A(n_132), .B(n_247), .Y(n_309) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_132), .Y(n_312) );
AND2x2_ASAP7_75t_L g420 ( .A(n_132), .B(n_247), .Y(n_420) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_163), .Y(n_132) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_133), .A2(n_180), .B(n_191), .Y(n_179) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_134), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_136), .B(n_137), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_160), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
INVx3_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_143), .Y(n_543) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
BUFx3_ASAP7_75t_L g236 ( .A(n_144), .Y(n_236) );
AND2x6_ASAP7_75t_L g480 ( .A(n_144), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_149), .A2(n_172), .B(n_173), .Y(n_171) );
INVx2_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_SL g205 ( .A1(n_149), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_149), .B(n_500), .Y(n_499) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_150), .A2(n_159), .B1(n_235), .B2(n_237), .Y(n_234) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
AND2x2_ASAP7_75t_L g476 ( .A(n_151), .B(n_156), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_151), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .C(n_158), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_154), .A2(n_177), .B(n_189), .C(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_154), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_177), .B1(n_197), .B2(n_199), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_177), .B1(n_250), .B2(n_251), .Y(n_249) );
INVx4_ASAP7_75t_L g554 ( .A(n_159), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g273 ( .A(n_160), .B(n_248), .C(n_249), .Y(n_273) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_161), .A2(n_171), .B(n_174), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_181), .B(n_188), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_205), .B(n_209), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_161), .A2(n_215), .B(n_220), .Y(n_214) );
AND2x4_ASAP7_75t_L g475 ( .A(n_161), .B(n_476), .Y(n_475) );
INVx4_ASAP7_75t_SL g489 ( .A(n_161), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_161), .B(n_476), .Y(n_563) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_164), .A2(n_204), .B(n_212), .Y(n_203) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_164), .A2(n_214), .B(n_223), .Y(n_213) );
INVx2_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_164), .A2(n_474), .B(n_477), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_164), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g535 ( .A(n_164), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_165), .B(n_312), .Y(n_368) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
OAI311xp33_ASAP7_75t_L g310 ( .A1(n_166), .A2(n_311), .A3(n_312), .B1(n_313), .C1(n_328), .Y(n_310) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
AND2x2_ASAP7_75t_L g271 ( .A(n_167), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g278 ( .A(n_167), .Y(n_278) );
AND2x2_ASAP7_75t_L g399 ( .A(n_167), .B(n_228), .Y(n_399) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_168), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g255 ( .A(n_168), .B(n_179), .Y(n_255) );
AND2x2_ASAP7_75t_L g307 ( .A(n_168), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_168), .B(n_254), .Y(n_321) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_178), .Y(n_168) );
INVx4_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_169), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_169), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
INVx2_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
AND2x2_ASAP7_75t_L g270 ( .A(n_179), .B(n_254), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_185), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_183), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_183), .A2(n_566), .B(n_567), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_185), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_210), .B(n_211), .Y(n_209) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g485 ( .A(n_187), .Y(n_485) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_200), .Y(n_192) );
OR2x2_ASAP7_75t_L g365 ( .A(n_193), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_193), .B(n_371), .Y(n_382) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_194), .B(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g239 ( .A(n_195), .Y(n_239) );
AND2x2_ASAP7_75t_L g306 ( .A(n_195), .B(n_233), .Y(n_306) );
AND2x2_ASAP7_75t_L g317 ( .A(n_195), .B(n_213), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_195), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_200), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_200), .B(n_267), .Y(n_311) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g298 ( .A(n_201), .B(n_257), .Y(n_298) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_213), .Y(n_201) );
INVx2_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
AND2x2_ASAP7_75t_L g325 ( .A(n_202), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
OR2x2_ASAP7_75t_L g342 ( .A(n_203), .B(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_203), .Y(n_405) );
AND2x2_ASAP7_75t_L g244 ( .A(n_213), .B(n_239), .Y(n_244) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g327 ( .A(n_213), .Y(n_327) );
INVx1_ASAP7_75t_L g343 ( .A(n_213), .Y(n_343) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_213), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_226), .B(n_331), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_226), .A2(n_316), .B1(n_365), .B2(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_227), .A2(n_409), .B(n_411), .C(n_429), .Y(n_408) );
INVx2_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
AND2x2_ASAP7_75t_L g319 ( .A(n_228), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_229), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g303 ( .A(n_230), .B(n_267), .Y(n_303) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g335 ( .A(n_231), .B(n_326), .Y(n_335) );
AND2x2_ASAP7_75t_L g354 ( .A(n_231), .B(n_268), .Y(n_354) );
AND2x4_ASAP7_75t_L g290 ( .A(n_232), .B(n_264), .Y(n_290) );
AND2x2_ASAP7_75t_L g428 ( .A(n_232), .B(n_404), .Y(n_428) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
INVx1_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
INVx1_ASAP7_75t_L g367 ( .A(n_233), .Y(n_367) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_236), .Y(n_487) );
INVx2_ASAP7_75t_L g555 ( .A(n_236), .Y(n_555) );
INVx1_ASAP7_75t_L g532 ( .A(n_238), .Y(n_532) );
OR2x2_ASAP7_75t_L g258 ( .A(n_239), .B(n_243), .Y(n_258) );
AND2x2_ASAP7_75t_L g267 ( .A(n_239), .B(n_268), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_239), .B(n_288), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .B1(n_256), .B2(n_259), .C(n_263), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_242), .A2(n_264), .B(n_266), .C(n_269), .Y(n_263) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_243), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_243), .B(n_265), .Y(n_371) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_243), .Y(n_378) );
AND2x2_ASAP7_75t_L g296 ( .A(n_244), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g333 ( .A(n_244), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
INVx2_ASAP7_75t_L g324 ( .A(n_246), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_246), .A2(n_257), .B1(n_374), .B2(n_376), .C1(n_377), .C2(n_379), .Y(n_373) );
AND2x2_ASAP7_75t_L g430 ( .A(n_246), .B(n_399), .Y(n_430) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
INVx1_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
AO21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_252), .Y(n_247) );
INVx3_ASAP7_75t_L g502 ( .A(n_248), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_248), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_248), .A2(n_538), .B(n_545), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_248), .B(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_248), .A2(n_561), .B(n_568), .Y(n_560) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g358 ( .A(n_255), .B(n_292), .Y(n_358) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_256), .A2(n_370), .B(n_372), .Y(n_369) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_257), .B(n_264), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_257), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx3_ASAP7_75t_L g323 ( .A(n_261), .Y(n_323) );
OR2x2_ASAP7_75t_L g375 ( .A(n_261), .B(n_297), .Y(n_375) );
AND2x2_ASAP7_75t_L g291 ( .A(n_262), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_262), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_262), .B(n_323), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_262), .B(n_319), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_262), .B(n_331), .Y(n_349) );
INVxp67_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_266), .A2(n_339), .B1(n_344), .B2(n_345), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_266), .B(n_371), .Y(n_401) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g387 ( .A(n_267), .B(n_378), .Y(n_387) );
AND2x2_ASAP7_75t_L g416 ( .A(n_267), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_267), .B(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g334 ( .A(n_268), .Y(n_334) );
BUFx2_ASAP7_75t_L g340 ( .A(n_268), .Y(n_340) );
INVx1_ASAP7_75t_L g425 ( .A(n_269), .Y(n_425) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_270), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g301 ( .A(n_271), .Y(n_301) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_272), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g284 ( .A(n_272), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g293 ( .A(n_272), .Y(n_293) );
INVx3_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
OR2x2_ASAP7_75t_L g397 ( .A(n_272), .B(n_398), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_282), .C(n_294), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_275), .A2(n_412), .B1(n_419), .B2(n_421), .C(n_422), .Y(n_411) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_289), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_285), .B(n_323), .Y(n_337) );
AND2x2_ASAP7_75t_L g379 ( .A(n_285), .B(n_319), .Y(n_379) );
INVx1_ASAP7_75t_SL g392 ( .A(n_286), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_286), .B(n_340), .Y(n_395) );
INVx1_ASAP7_75t_L g413 ( .A(n_287), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_291), .A2(n_381), .B1(n_383), .B2(n_387), .C(n_388), .Y(n_380) );
AND2x2_ASAP7_75t_L g407 ( .A(n_292), .B(n_399), .Y(n_407) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g391 ( .A(n_293), .Y(n_391) );
AOI21xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_298), .B(n_299), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g362 ( .A(n_297), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
INVx1_ASAP7_75t_L g376 ( .A(n_299), .Y(n_376) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_310), .Y(n_302) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_303), .A2(n_341), .A3(n_428), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g403 ( .A(n_306), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g424 ( .A(n_306), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_308), .B(n_323), .Y(n_351) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g426 ( .A(n_309), .B(n_323), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B1(n_322), .B2(n_325), .Y(n_313) );
NAND2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_317), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g356 ( .A(n_317), .B(n_340), .Y(n_356) );
AND2x2_ASAP7_75t_L g410 ( .A(n_317), .B(n_405), .Y(n_410) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_323), .A2(n_357), .A3(n_389), .B1(n_391), .B2(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_326), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_336), .C(n_338), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_334), .B(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_335), .A2(n_347), .B1(n_348), .B2(n_349), .C(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_345), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_355), .B2(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND4xp25_ASAP7_75t_SL g412 ( .A(n_355), .B(n_413), .C(n_414), .D(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_373), .C(n_380), .D(n_393), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_368), .C(n_369), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g390 ( .A(n_366), .Y(n_390) );
INVx2_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
OR2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_400), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_399), .B(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B(n_406), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g440 ( .A(n_433), .Y(n_440) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g444 ( .A(n_434), .Y(n_444) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_441), .B(n_446), .C(n_447), .D(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_459), .B2(n_766), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_465), .B2(n_468), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g767 ( .A(n_461), .Y(n_767) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g768 ( .A(n_463), .Y(n_768) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g769 ( .A(n_466), .Y(n_769) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g770 ( .A(n_468), .Y(n_770) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR5x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_639), .C(n_717), .D(n_741), .E(n_758), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_511), .B(n_557), .C(n_616), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_491), .Y(n_471) );
AND2x2_ASAP7_75t_L g570 ( .A(n_472), .B(n_493), .Y(n_570) );
INVx5_ASAP7_75t_SL g598 ( .A(n_472), .Y(n_598) );
AND2x2_ASAP7_75t_L g634 ( .A(n_472), .B(n_619), .Y(n_634) );
OR2x2_ASAP7_75t_L g673 ( .A(n_472), .B(n_492), .Y(n_673) );
OR2x2_ASAP7_75t_L g704 ( .A(n_472), .B(n_595), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_472), .B(n_608), .Y(n_740) );
AND2x2_ASAP7_75t_L g752 ( .A(n_472), .B(n_595), .Y(n_752) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_490), .Y(n_472) );
BUFx2_ASAP7_75t_L g527 ( .A(n_475), .Y(n_527) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_479), .A2(n_489), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_479), .A2(n_489), .B(n_550), .C(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .C(n_487), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_484), .A2(n_487), .B(n_519), .C(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g751 ( .A(n_491), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g614 ( .A(n_492), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_503), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_493), .B(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_493), .Y(n_607) );
INVx3_ASAP7_75t_L g622 ( .A(n_493), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_493), .B(n_503), .Y(n_646) );
OR2x2_ASAP7_75t_L g655 ( .A(n_493), .B(n_598), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_493), .B(n_619), .Y(n_659) );
AND2x2_ASAP7_75t_L g665 ( .A(n_493), .B(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g702 ( .A(n_493), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_493), .B(n_560), .Y(n_716) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_493) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_502), .A2(n_548), .B(n_556), .Y(n_547) );
OR2x2_ASAP7_75t_L g608 ( .A(n_503), .B(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_L g619 ( .A(n_503), .B(n_595), .Y(n_619) );
AND2x2_ASAP7_75t_L g631 ( .A(n_503), .B(n_622), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_503), .B(n_560), .Y(n_654) );
INVx1_ASAP7_75t_SL g666 ( .A(n_503), .Y(n_666) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g559 ( .A(n_504), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_504), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
AND2x2_ASAP7_75t_L g579 ( .A(n_513), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_513), .B(n_536), .Y(n_583) );
AND2x2_ASAP7_75t_L g586 ( .A(n_513), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_513), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g611 ( .A(n_513), .B(n_602), .Y(n_611) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_513), .Y(n_630) );
AND2x2_ASAP7_75t_L g651 ( .A(n_513), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g661 ( .A(n_513), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g707 ( .A(n_513), .B(n_590), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_513), .B(n_613), .Y(n_734) );
INVx5_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g604 ( .A(n_514), .Y(n_604) );
AND2x2_ASAP7_75t_L g670 ( .A(n_514), .B(n_602), .Y(n_670) );
AND2x2_ASAP7_75t_L g754 ( .A(n_514), .B(n_622), .Y(n_754) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_521), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_523), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_523), .Y(n_743) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
AND2x2_ASAP7_75t_L g573 ( .A(n_524), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g582 ( .A(n_524), .B(n_580), .Y(n_582) );
INVx5_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g613 ( .A(n_524), .B(n_547), .Y(n_613) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_526), .A2(n_528), .B(n_532), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g691 ( .A(n_536), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_536), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g724 ( .A(n_536), .B(n_590), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_536), .A2(n_647), .B(n_754), .C(n_755), .Y(n_753) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
BUFx2_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
INVx2_ASAP7_75t_L g578 ( .A(n_537), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .Y(n_538) );
INVx2_ASAP7_75t_L g580 ( .A(n_547), .Y(n_580) );
AND2x2_ASAP7_75t_L g587 ( .A(n_547), .B(n_578), .Y(n_587) );
AND2x2_ASAP7_75t_L g678 ( .A(n_547), .B(n_590), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI211x1_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_571), .B(n_584), .C(n_609), .Y(n_557) );
INVx1_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_570), .Y(n_558) );
INVx5_ASAP7_75t_SL g595 ( .A(n_560), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_560), .B(n_665), .Y(n_664) );
AOI311xp33_ASAP7_75t_L g683 ( .A1(n_560), .A2(n_684), .A3(n_686), .B(n_687), .C(n_693), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_560), .A2(n_631), .B(n_719), .C(n_722), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_564), .Y(n_561) );
INVxp67_ASAP7_75t_L g638 ( .A(n_570), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g571 ( .A(n_572), .B(n_575), .C(n_581), .D(n_583), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_572), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g629 ( .A(n_573), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_576), .B(n_582), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_576), .B(n_589), .Y(n_709) );
BUFx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_577), .B(n_590), .Y(n_727) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g602 ( .A(n_578), .Y(n_602) );
INVxp67_ASAP7_75t_L g637 ( .A(n_579), .Y(n_637) );
AND2x4_ASAP7_75t_L g589 ( .A(n_580), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g663 ( .A(n_580), .B(n_602), .Y(n_663) );
INVx1_ASAP7_75t_L g690 ( .A(n_580), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_580), .B(n_677), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_581), .B(n_651), .Y(n_671) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_582), .B(n_604), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_582), .B(n_651), .Y(n_750) );
INVx1_ASAP7_75t_L g761 ( .A(n_583), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_588), .B(n_591), .C(n_599), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
AND2x2_ASAP7_75t_L g600 ( .A(n_589), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_589), .B(n_651), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_589), .B(n_670), .Y(n_694) );
OR2x2_ASAP7_75t_L g610 ( .A(n_590), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g642 ( .A(n_590), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_590), .B(n_602), .Y(n_657) );
AND2x2_ASAP7_75t_L g714 ( .A(n_590), .B(n_670), .Y(n_714) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_590), .Y(n_721) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_592), .A2(n_604), .B1(n_726), .B2(n_728), .C(n_731), .Y(n_725) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g615 ( .A(n_595), .B(n_598), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_595), .B(n_665), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_595), .B(n_622), .Y(n_730) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g715 ( .A(n_597), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g729 ( .A(n_597), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_598), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g626 ( .A(n_598), .B(n_619), .Y(n_626) );
AND2x2_ASAP7_75t_L g696 ( .A(n_598), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_598), .B(n_645), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_598), .B(n_746), .Y(n_745) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_605), .Y(n_599) );
INVx2_ASAP7_75t_L g632 ( .A(n_600), .Y(n_632) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g652 ( .A(n_602), .Y(n_652) );
OR2x2_ASAP7_75t_L g656 ( .A(n_604), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g759 ( .A(n_604), .B(n_727), .Y(n_759) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_612), .B(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g763 ( .A(n_610), .Y(n_763) );
INVx2_ASAP7_75t_SL g677 ( .A(n_611), .Y(n_677) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_614), .A2(n_695), .B(n_759), .C(n_760), .Y(n_758) );
OAI322xp33_ASAP7_75t_SL g627 ( .A1(n_615), .A2(n_628), .A3(n_631), .B1(n_632), .B2(n_633), .C1(n_635), .C2(n_638), .Y(n_627) );
INVx2_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .B1(n_624), .B2(n_626), .C(n_627), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_SL g693 ( .A1(n_618), .A2(n_694), .B1(n_695), .B2(n_698), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_619), .B(n_622), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_619), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g692 ( .A(n_621), .B(n_654), .Y(n_692) );
INVx1_ASAP7_75t_L g682 ( .A(n_622), .Y(n_682) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_626), .A2(n_736), .B(n_738), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_628), .A2(n_661), .B(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g689 ( .A(n_630), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_630), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g746 ( .A(n_631), .Y(n_746) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_667), .C(n_683), .D(n_699), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_648), .C(n_660), .Y(n_640) );
INVx1_ASAP7_75t_L g732 ( .A(n_641), .Y(n_732) );
AND2x2_ASAP7_75t_L g680 ( .A(n_642), .B(n_663), .Y(n_680) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_647), .B(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B1(n_656), .B2(n_658), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_650), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g698 ( .A(n_651), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_651), .A2(n_690), .B(n_713), .C(n_715), .Y(n_712) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g697 ( .A(n_654), .Y(n_697) );
INVx1_ASAP7_75t_L g757 ( .A(n_655), .Y(n_757) );
NAND2xp33_ASAP7_75t_SL g747 ( .A(n_656), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g686 ( .A(n_665), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B(n_672), .C(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_679), .B2(n_681), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_677), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_682), .B(n_703), .Y(n_765) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_691), .B(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_705), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_715), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
NAND3xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_725), .C(n_735), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B(n_744), .C(n_753), .Y(n_741) );
INVx1_ASAP7_75t_L g762 ( .A(n_742), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_747), .B1(n_749), .B2(n_751), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI22x1_ASAP7_75t_SL g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
endmodule