module fake_jpeg_4533_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_47),
.B1(n_69),
.B2(n_26),
.Y(n_72)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_24),
.B1(n_31),
.B2(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_17),
.B1(n_25),
.B2(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_43),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_87),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_43),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_43),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_18),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_68),
.B1(n_62),
.B2(n_65),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_17),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_54),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_102),
.B1(n_110),
.B2(n_117),
.Y(n_130)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_43),
.B(n_25),
.C(n_66),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_107),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_20),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_111),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_56),
.B(n_30),
.Y(n_107)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_29),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_29),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_29),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_83),
.B1(n_82),
.B2(n_76),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_51),
.B1(n_89),
.B2(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_128),
.B1(n_131),
.B2(n_120),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_77),
.C(n_35),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_33),
.C(n_23),
.Y(n_168)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_133),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_89),
.B1(n_84),
.B2(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_93),
.B1(n_84),
.B2(n_30),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_93),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_139),
.B(n_23),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_114),
.Y(n_156)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_63),
.B(n_64),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_73),
.B1(n_45),
.B2(n_48),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_73),
.B1(n_32),
.B2(n_36),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_147),
.B1(n_88),
.B2(n_86),
.Y(n_153)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_110),
.B1(n_102),
.B2(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_109),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_165),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_110),
.B1(n_105),
.B2(n_96),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_166),
.B(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_103),
.B1(n_119),
.B2(n_97),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_174),
.B1(n_130),
.B2(n_121),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_109),
.B1(n_111),
.B2(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_116),
.B1(n_114),
.B2(n_86),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_104),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_98),
.B(n_32),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_33),
.B(n_23),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_49),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_164),
.C(n_168),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_36),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_88),
.CI(n_29),
.CON(n_165),
.SN(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_23),
.B(n_33),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_23),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_126),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_125),
.B1(n_137),
.B2(n_145),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_33),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_63),
.B1(n_33),
.B2(n_23),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_144),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_193),
.C(n_168),
.Y(n_204)
);

XOR2x2_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_142),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_150),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_138),
.A3(n_137),
.B1(n_125),
.B2(n_126),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_186),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_147),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_187),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_133),
.C(n_124),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_194),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_33),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_22),
.B(n_1),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_155),
.B(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_172),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_209),
.C(n_182),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_159),
.C(n_158),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_191),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_216),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_154),
.B1(n_173),
.B2(n_150),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_162),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_219),
.B(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_165),
.B(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_199),
.B1(n_194),
.B2(n_195),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_22),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVxp33_ASAP7_75t_SL g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_206),
.B(n_177),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_232),
.C(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_236),
.B1(n_202),
.B2(n_208),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_193),
.C(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_187),
.C(n_184),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_184),
.C(n_181),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_186),
.C(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_242),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_178),
.B(n_183),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_253),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_212),
.B1(n_211),
.B2(n_205),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_256),
.B1(n_235),
.B2(n_1),
.Y(n_269)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_219),
.B1(n_220),
.B2(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_221),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_201),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_22),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_232),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_229),
.B1(n_234),
.B2(n_9),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_233),
.C(n_228),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_264),
.A2(n_270),
.B(n_260),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_235),
.B1(n_8),
.B2(n_9),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_278),
.B1(n_11),
.B2(n_13),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_273),
.B(n_12),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_0),
.C(n_3),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_8),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_7),
.B(n_13),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_10),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_261),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_290),
.C(n_275),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_247),
.B(n_259),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_250),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_10),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_288),
.B(n_12),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_0),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.C(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_266),
.C(n_268),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_274),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_280),
.CI(n_283),
.CON(n_303),
.SN(n_303)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_299),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_10),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_297),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_303),
.B(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_13),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_293),
.B1(n_15),
.B2(n_298),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_15),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_302),
.C(n_308),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_312),
.C(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_310),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_5),
.B(n_6),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_5),
.C(n_6),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_5),
.Y(n_320)
);


endmodule