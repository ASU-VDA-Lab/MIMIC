module fake_jpeg_12696_n_46 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_27),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_2),
.A3(n_10),
.B1(n_19),
.B2(n_17),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_15),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.C(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_23),
.C(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_11),
.B(n_18),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.C(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_11),
.B1(n_12),
.B2(n_28),
.Y(n_35)
);

OA21x2_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_30),
.B(n_26),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.C(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OA21x2_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_32),
.B(n_37),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_40),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);


endmodule