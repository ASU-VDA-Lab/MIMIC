module fake_netlist_1_6767_n_33 (n_1, n_2, n_4, n_3, n_5, n_0, n_33);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_6;
wire n_7;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_0), .Y(n_9) );
INVx1_ASAP7_75t_SL g10 ( .A(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
NOR2xp33_ASAP7_75t_SL g13 ( .A(n_7), .B(n_1), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_1), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_6), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_1), .B(n_2), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_11), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_12), .B(n_7), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_8), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_17), .B(n_13), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_17), .B(n_13), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NOR4xp25_ASAP7_75t_SL g25 ( .A(n_23), .B(n_10), .C(n_3), .D(n_5), .Y(n_25) );
A2O1A1Ixp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_22), .B(n_21), .C(n_16), .Y(n_26) );
NAND4xp25_ASAP7_75t_L g27 ( .A(n_24), .B(n_10), .C(n_20), .D(n_22), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
NOR2x1_ASAP7_75t_SL g30 ( .A(n_26), .B(n_19), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_19), .B1(n_27), .B2(n_2), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI22xp33_ASAP7_75t_R g33 ( .A1(n_32), .A2(n_5), .B1(n_30), .B2(n_31), .Y(n_33) );
endmodule