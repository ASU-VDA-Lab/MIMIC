module fake_netlist_6_2907_n_1284 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1284);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1284;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_367;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx2_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_72),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_278),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_123),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_171),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_67),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_15),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_64),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_121),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_223),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_173),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_111),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_96),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_112),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_79),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_251),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_22),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_219),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_57),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_213),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_22),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_151),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_133),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_163),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_8),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_147),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_44),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_156),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_184),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_204),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_143),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_104),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_99),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_228),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_217),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_277),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_8),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_158),
.B(n_29),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_92),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_80),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_18),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_134),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_66),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_164),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_264),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_280),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_76),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_128),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_167),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_12),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_196),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_235),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_47),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_140),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_247),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_138),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_129),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_135),
.B(n_5),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_153),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_110),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_95),
.B(n_154),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_214),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_194),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_159),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_137),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_28),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_255),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_90),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_125),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_180),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_209),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_1),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_177),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_19),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_36),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_40),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_275),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_240),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_242),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_263),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_181),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_203),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_51),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_226),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_152),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_172),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_24),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_106),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_141),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_34),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_83),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_165),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_116),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_232),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_274),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_179),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_117),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_197),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_169),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_145),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_86),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_14),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_55),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_239),
.Y(n_411)
);

BUFx5_ASAP7_75t_L g412 ( 
.A(n_109),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_160),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_208),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_119),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_15),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_227),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_75),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_144),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_98),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_70),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_245),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_187),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_19),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_12),
.Y(n_426)
);

INVx4_ASAP7_75t_R g427 ( 
.A(n_53),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_284),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_220),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_63),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_101),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_256),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_11),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_265),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_189),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_105),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_270),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_102),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_150),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_161),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_200),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_146),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_89),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_11),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_14),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_41),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_192),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_259),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_246),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_221),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_233),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_257),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_269),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_45),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_237),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_50),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_85),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_2),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_132),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_193),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_46),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_71),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_126),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_94),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_215),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_78),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_122),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_21),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_139),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_178),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_231),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_28),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_18),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_176),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_234),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_59),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_93),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_229),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_50),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_207),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_199),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_29),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_224),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_253),
.Y(n_484)
);

BUFx5_ASAP7_75t_L g485 ( 
.A(n_16),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_107),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_4),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_60),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_43),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_250),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_73),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_16),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_91),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_485),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_287),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_485),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_287),
.B(n_58),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_290),
.A2(n_0),
.B(n_1),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_287),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_287),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_378),
.B(n_2),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_3),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

OAI22x1_ASAP7_75t_R g506 ( 
.A1(n_368),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

BUFx8_ASAP7_75t_SL g508 ( 
.A(n_379),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_308),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_305),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_6),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_305),
.Y(n_513)
);

BUFx8_ASAP7_75t_SL g514 ( 
.A(n_474),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_7),
.Y(n_515)
);

BUFx8_ASAP7_75t_SL g516 ( 
.A(n_483),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_378),
.B(n_7),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_294),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_310),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_305),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_305),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_322),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_307),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_292),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_319),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_335),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_308),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_308),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_376),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_308),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_393),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_381),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_366),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_366),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_419),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_359),
.B(n_61),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_313),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_444),
.B(n_9),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_366),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_366),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_297),
.B(n_10),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_374),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_374),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_351),
.A2(n_13),
.B1(n_17),
.B2(n_20),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_317),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_340),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_350),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_286),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_374),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_353),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_345),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_288),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_295),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_299),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_382),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_412),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_466),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_334),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_312),
.B(n_23),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_289),
.B(n_25),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_424),
.B(n_26),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_301),
.Y(n_570)
);

OAI22x1_ASAP7_75t_SL g571 ( 
.A1(n_389),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_285),
.B(n_62),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_326),
.A2(n_68),
.B(n_65),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_375),
.B(n_27),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_412),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_412),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_380),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_412),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_343),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_392),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_291),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_293),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_405),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_296),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_358),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_437),
.A2(n_460),
.B(n_303),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_312),
.B(n_31),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_298),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_302),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_304),
.Y(n_590)
);

OAI22x1_ASAP7_75t_L g591 ( 
.A1(n_396),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_591)
);

BUFx8_ASAP7_75t_SL g592 ( 
.A(n_372),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_309),
.A2(n_74),
.B(n_69),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_331),
.B(n_32),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

CKINVDCx6p67_ASAP7_75t_R g596 ( 
.A(n_467),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_321),
.B(n_325),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_327),
.B(n_33),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_478),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_328),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_306),
.Y(n_601)
);

OAI22x1_ASAP7_75t_SL g602 ( 
.A1(n_410),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_329),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_426),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_362),
.B(n_77),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_333),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_433),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_478),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_336),
.B(n_38),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_341),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_348),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_356),
.Y(n_613)
);

BUFx8_ASAP7_75t_SL g614 ( 
.A(n_390),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_397),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_357),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_360),
.B(n_39),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_363),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_311),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_314),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_364),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_377),
.A2(n_82),
.B(n_81),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_445),
.Y(n_623)
);

OA21x2_ASAP7_75t_L g624 ( 
.A1(n_385),
.A2(n_40),
.B(n_41),
.Y(n_624)
);

INVx6_ASAP7_75t_L g625 ( 
.A(n_427),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_454),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_394),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_316),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_487),
.B(n_42),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_395),
.B(n_398),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_399),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_401),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_458),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_413),
.B(n_43),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_468),
.Y(n_635)
);

CKINVDCx6p67_ASAP7_75t_R g636 ( 
.A(n_418),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_582),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_551),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_563),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_584),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_585),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_R g642 ( 
.A(n_523),
.B(n_472),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_R g643 ( 
.A(n_524),
.B(n_455),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_600),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_610),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_581),
.B(n_300),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_612),
.B(n_413),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_592),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_555),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_635),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_542),
.A2(n_337),
.B1(n_469),
.B2(n_462),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_R g652 ( 
.A(n_556),
.B(n_557),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_606),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_614),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_611),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_570),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_550),
.A2(n_473),
.B1(n_489),
.B2(n_480),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_496),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_589),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_601),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_613),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_616),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_621),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_500),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_619),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_503),
.B(n_538),
.C(n_566),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_522),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_579),
.B(n_477),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_500),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_631),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_615),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_508),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_500),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_636),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_514),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_574),
.B(n_300),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_R g678 ( 
.A(n_635),
.B(n_599),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_516),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_620),
.B(n_512),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_577),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_625),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_502),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_502),
.Y(n_684)
);

NOR2x1p5_ASAP7_75t_L g685 ( 
.A(n_596),
.B(n_315),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_502),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_R g687 ( 
.A(n_623),
.B(n_318),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_574),
.B(n_493),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_633),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_577),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_547),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_511),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_577),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_511),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_558),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_511),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_604),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_625),
.B(n_320),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_513),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_576),
.B(n_323),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_562),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_595),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_608),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_513),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_537),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_612),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_580),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_549),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_626),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_513),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_504),
.B(n_403),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_576),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_583),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_554),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_583),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_564),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_583),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_628),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_507),
.B(n_344),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_R g721 ( 
.A(n_517),
.B(n_324),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_509),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_597),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_597),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_658),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_605),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_650),
.B(n_586),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_657),
.B(n_546),
.C(n_587),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_678),
.B(n_517),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_642),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_677),
.B(n_495),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_680),
.B(n_677),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_674),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_653),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_652),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_704),
.Y(n_737)
);

AO221x1_ASAP7_75t_L g738 ( 
.A1(n_722),
.A2(n_591),
.B1(n_411),
.B2(n_422),
.C(n_421),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_680),
.B(n_521),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_704),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_655),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_664),
.B(n_521),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_670),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_720),
.B(n_512),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_661),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_662),
.B(n_494),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_683),
.B(n_521),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_715),
.B(n_629),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_684),
.B(n_540),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_686),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_692),
.B(n_540),
.Y(n_751)
);

AO221x1_ASAP7_75t_L g752 ( 
.A1(n_668),
.A2(n_431),
.B1(n_432),
.B2(n_423),
.C(n_408),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_709),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_699),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_651),
.A2(n_634),
.B1(n_594),
.B2(n_571),
.C(n_602),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_670),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_670),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_663),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_688),
.B(n_540),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_710),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_643),
.B(n_568),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_656),
.B(n_545),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_723),
.B(n_724),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_688),
.B(n_545),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_646),
.B(n_691),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_659),
.B(n_545),
.Y(n_766)
);

INVxp33_ASAP7_75t_L g767 ( 
.A(n_669),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_701),
.B(n_630),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_666),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_694),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_695),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_672),
.B(n_567),
.C(n_535),
.Y(n_772)
);

BUFx6f_ASAP7_75t_SL g773 ( 
.A(n_671),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_609),
.C(n_598),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_660),
.B(n_568),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_697),
.B(n_607),
.C(n_553),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_681),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_690),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_694),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_712),
.B(n_497),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_693),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_609),
.C(n_598),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_665),
.B(n_630),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_687),
.B(n_515),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_705),
.A2(n_622),
.B(n_593),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_702),
.B(n_515),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_703),
.B(n_617),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_696),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_711),
.Y(n_790)
);

BUFx5_ASAP7_75t_L g791 ( 
.A(n_712),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_708),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_637),
.B(n_617),
.C(n_499),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_700),
.B(n_698),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_714),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_712),
.B(n_501),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_711),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_685),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_712),
.B(n_505),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_707),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_716),
.B(n_510),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_718),
.B(n_527),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_640),
.B(n_532),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_735),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_794),
.B(n_761),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_741),
.B(n_518),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_727),
.A2(n_645),
.B(n_644),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_744),
.B(n_499),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_745),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_727),
.A2(n_530),
.B(n_528),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_758),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

BUFx5_ASAP7_75t_L g813 ( 
.A(n_769),
.Y(n_813)
);

BUFx4f_ASAP7_75t_L g814 ( 
.A(n_798),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_775),
.A2(n_573),
.B(n_536),
.C(n_439),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_730),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_733),
.B(n_436),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_803),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_765),
.B(n_706),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_728),
.A2(n_605),
.B1(n_417),
.B2(n_442),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_776),
.B(n_682),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_801),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_731),
.B(n_605),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_726),
.A2(n_605),
.B1(n_624),
.B2(n_572),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_801),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_731),
.B(n_647),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_753),
.B(n_675),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_775),
.A2(n_441),
.B(n_449),
.C(n_447),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_783),
.A2(n_355),
.B1(n_332),
.B2(n_338),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_760),
.B(n_719),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_759),
.B(n_764),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_768),
.Y(n_832)
);

BUFx8_ASAP7_75t_SL g833 ( 
.A(n_736),
.Y(n_833)
);

OAI21xp33_ASAP7_75t_L g834 ( 
.A1(n_787),
.A2(n_525),
.B(n_519),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_783),
.B(n_689),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_750),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_802),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_772),
.A2(n_339),
.B1(n_342),
.B2(n_330),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_802),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_754),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_785),
.B(n_572),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_791),
.B(n_498),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_729),
.B(n_624),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_746),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_771),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_756),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_762),
.B(n_572),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_743),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_777),
.A2(n_347),
.B1(n_349),
.B2(n_346),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_766),
.B(n_572),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_SL g852 ( 
.A1(n_738),
.A2(n_713),
.B1(n_639),
.B2(n_641),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_800),
.B(n_711),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_784),
.B(n_452),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_793),
.A2(n_748),
.B1(n_796),
.B2(n_781),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_780),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_788),
.B(n_780),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_757),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_778),
.B(n_526),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_796),
.A2(n_531),
.B(n_539),
.C(n_529),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_725),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_780),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_763),
.B(n_638),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_767),
.B(n_649),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_779),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_782),
.B(n_548),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_739),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_789),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_793),
.B(n_453),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_770),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_774),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_SL g872 ( 
.A(n_755),
.B(n_679),
.C(n_676),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_732),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_SL g874 ( 
.A1(n_792),
.A2(n_673),
.B1(n_648),
.B2(n_654),
.Y(n_874)
);

AND2x6_ASAP7_75t_SL g875 ( 
.A(n_795),
.B(n_506),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_734),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_737),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_740),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_790),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_797),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_773),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_773),
.A2(n_717),
.B1(n_565),
.B2(n_569),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_799),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_841),
.B(n_791),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_833),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_883),
.A2(n_855),
.B1(n_845),
.B2(n_820),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_823),
.A2(n_752),
.B(n_476),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_822),
.B(n_825),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_883),
.A2(n_481),
.B(n_484),
.C(n_457),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_817),
.A2(n_498),
.B1(n_486),
.B2(n_791),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_837),
.B(n_791),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_816),
.B(n_789),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_839),
.B(n_786),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_832),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_826),
.B(n_786),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_869),
.A2(n_843),
.B(n_831),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_809),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_819),
.B(n_352),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_824),
.A2(n_747),
.B(n_742),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_846),
.B(n_560),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_864),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_804),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_811),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_847),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_807),
.A2(n_749),
.B(n_751),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_862),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_805),
.B(n_354),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_842),
.A2(n_533),
.B(n_520),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_818),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_862),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_813),
.B(n_361),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_810),
.A2(n_534),
.B(n_533),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_865),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_870),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_813),
.B(n_365),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_828),
.A2(n_561),
.B(n_575),
.C(n_578),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_821),
.B(n_367),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_813),
.B(n_369),
.Y(n_918)
);

OAI21xp33_ASAP7_75t_SL g919 ( 
.A1(n_854),
.A2(n_552),
.B(n_543),
.Y(n_919)
);

AOI22x1_ASAP7_75t_L g920 ( 
.A1(n_844),
.A2(n_434),
.B1(n_370),
.B2(n_371),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_808),
.A2(n_541),
.B(n_534),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_860),
.A2(n_532),
.B(n_544),
.C(n_559),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_SL g924 ( 
.A1(n_835),
.A2(n_552),
.B(n_543),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_817),
.A2(n_498),
.B1(n_618),
.B2(n_603),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_874),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_867),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_830),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_861),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_850),
.A2(n_435),
.B(n_383),
.C(n_384),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_813),
.B(n_373),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_817),
.B(n_386),
.Y(n_932)
);

AO21x2_ASAP7_75t_L g933 ( 
.A1(n_815),
.A2(n_498),
.B(n_388),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_817),
.B(n_387),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_806),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_827),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_868),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_806),
.B(n_391),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_859),
.B(n_544),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_R g940 ( 
.A(n_872),
.B(n_400),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_848),
.A2(n_559),
.B(n_402),
.C(n_450),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_873),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_866),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_882),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_829),
.B(n_404),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_849),
.A2(n_856),
.B(n_812),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_881),
.B(n_857),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_836),
.B(n_406),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_838),
.B(n_407),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_840),
.B(n_414),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_944),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_897),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_895),
.A2(n_851),
.B(n_879),
.Y(n_953)
);

AOI22x1_ASAP7_75t_L g954 ( 
.A1(n_896),
.A2(n_880),
.B1(n_876),
.B2(n_877),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_905),
.A2(n_847),
.B(n_853),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_893),
.A2(n_834),
.B(n_812),
.Y(n_956)
);

BUFx2_ASAP7_75t_SL g957 ( 
.A(n_885),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_937),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_913),
.Y(n_960)
);

AOI22x1_ASAP7_75t_L g961 ( 
.A1(n_899),
.A2(n_878),
.B1(n_866),
.B2(n_856),
.Y(n_961)
);

CKINVDCx16_ASAP7_75t_R g962 ( 
.A(n_927),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_901),
.Y(n_963)
);

INVx5_ASAP7_75t_SL g964 ( 
.A(n_947),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_903),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_888),
.B(n_868),
.Y(n_966)
);

INVx6_ASAP7_75t_SL g967 ( 
.A(n_900),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_936),
.B(n_863),
.Y(n_968)
);

INVx6_ASAP7_75t_L g969 ( 
.A(n_937),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_914),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_922),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_926),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_886),
.A2(n_849),
.B(n_868),
.Y(n_973)
);

XOR2xp5_ASAP7_75t_L g974 ( 
.A(n_935),
.B(n_852),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_917),
.B(n_858),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_884),
.A2(n_814),
.B(n_871),
.Y(n_976)
);

CKINVDCx16_ASAP7_75t_R g977 ( 
.A(n_940),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_891),
.A2(n_849),
.B(n_814),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_941),
.A2(n_889),
.B(n_930),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_904),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_922),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_946),
.A2(n_88),
.B(n_84),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_928),
.B(n_898),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_906),
.B(n_588),
.Y(n_984)
);

AO21x2_ASAP7_75t_L g985 ( 
.A1(n_911),
.A2(n_603),
.B(n_590),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_904),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_909),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_908),
.A2(n_100),
.B(n_97),
.Y(n_988)
);

AO21x2_ASAP7_75t_L g989 ( 
.A1(n_915),
.A2(n_603),
.B(n_590),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_921),
.A2(n_108),
.B(n_103),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_947),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_939),
.Y(n_992)
);

AO21x2_ASAP7_75t_L g993 ( 
.A1(n_933),
.A2(n_618),
.B(n_590),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_920),
.A2(n_114),
.B(n_113),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_916),
.A2(n_428),
.B(n_415),
.Y(n_995)
);

AO21x2_ASAP7_75t_L g996 ( 
.A1(n_933),
.A2(n_632),
.B(n_618),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_922),
.Y(n_997)
);

BUFx2_ASAP7_75t_R g998 ( 
.A(n_887),
.Y(n_998)
);

AO21x2_ASAP7_75t_L g999 ( 
.A1(n_918),
.A2(n_632),
.B(n_430),
.Y(n_999)
);

BUFx4f_ASAP7_75t_L g1000 ( 
.A(n_943),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_906),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_910),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_912),
.A2(n_118),
.B(n_115),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_902),
.B(n_429),
.Y(n_1004)
);

AO21x2_ASAP7_75t_L g1005 ( 
.A1(n_931),
.A2(n_632),
.B(n_440),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_949),
.A2(n_465),
.B1(n_491),
.B2(n_475),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_910),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_945),
.A2(n_459),
.B1(n_471),
.B2(n_470),
.Y(n_1008)
);

BUFx8_ASAP7_75t_SL g1009 ( 
.A(n_929),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_892),
.Y(n_1010)
);

AND2x2_ASAP7_75t_SL g1011 ( 
.A(n_907),
.B(n_925),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_970),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_952),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_958),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_960),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_987),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_965),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_959),
.B(n_942),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_980),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_SL g1021 ( 
.A1(n_1011),
.A2(n_887),
.B1(n_938),
.B2(n_875),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_958),
.Y(n_1022)
);

OAI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_1010),
.A2(n_934),
.B1(n_932),
.B2(n_948),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_983),
.B(n_950),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_980),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_975),
.A2(n_890),
.B1(n_919),
.B2(n_924),
.Y(n_1026)
);

BUFx8_ASAP7_75t_SL g1027 ( 
.A(n_972),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_SL g1028 ( 
.A1(n_977),
.A2(n_438),
.B1(n_448),
.B2(n_451),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_955),
.A2(n_923),
.B(n_191),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_963),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_1007),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_SL g1032 ( 
.A1(n_974),
.A2(n_1006),
.B(n_1008),
.Y(n_1032)
);

OAI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_975),
.A2(n_464),
.B1(n_45),
.B2(n_46),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_SL g1034 ( 
.A1(n_972),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1008),
.A2(n_1006),
.B1(n_968),
.B2(n_979),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_986),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_986),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_991),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_966),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_966),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_969),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_954),
.A2(n_198),
.B(n_279),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_992),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_961),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_971),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_968),
.B(n_1004),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1004),
.B(n_48),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_971),
.Y(n_1048)
);

BUFx2_ASAP7_75t_R g1049 ( 
.A(n_957),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_971),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_969),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_971),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_981),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_981),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_981),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_981),
.Y(n_1056)
);

OA21x2_ASAP7_75t_L g1057 ( 
.A1(n_956),
.A2(n_49),
.B(n_52),
.Y(n_1057)
);

BUFx2_ASAP7_75t_R g1058 ( 
.A(n_1009),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_995),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_995),
.A2(n_976),
.B1(n_1000),
.B2(n_1005),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_973),
.A2(n_54),
.B(n_56),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_953),
.A2(n_205),
.B(n_120),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_997),
.Y(n_1063)
);

BUFx4f_ASAP7_75t_SL g1064 ( 
.A(n_967),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1009),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1013),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1012),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_1024),
.B(n_1000),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_1014),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1059),
.A2(n_998),
.B1(n_964),
.B2(n_1007),
.Y(n_1070)
);

NAND2xp33_ASAP7_75t_SL g1071 ( 
.A(n_1030),
.B(n_951),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1016),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_R g1073 ( 
.A(n_1064),
.B(n_962),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1018),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1021),
.B(n_964),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1032),
.B(n_951),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1021),
.B(n_964),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1046),
.B(n_1002),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_SL g1079 ( 
.A(n_1023),
.B(n_976),
.C(n_998),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1039),
.B(n_999),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1035),
.A2(n_999),
.B1(n_1005),
.B2(n_989),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1015),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_1014),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_1041),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1022),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1040),
.B(n_1001),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1012),
.B(n_997),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1022),
.B(n_997),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1023),
.B(n_978),
.C(n_994),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1017),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_1017),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1035),
.B(n_985),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1051),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1028),
.B(n_984),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_1041),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_1038),
.B(n_982),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_1065),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1028),
.B(n_993),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1033),
.A2(n_996),
.B(n_993),
.C(n_989),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_1043),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1037),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1047),
.B(n_1020),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1059),
.A2(n_996),
.B1(n_985),
.B2(n_57),
.C(n_1003),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1061),
.A2(n_988),
.B(n_990),
.C(n_130),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1048),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1019),
.B(n_124),
.Y(n_1106)
);

AND2x2_ASAP7_75t_SL g1107 ( 
.A(n_1060),
.B(n_127),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1020),
.B(n_131),
.Y(n_1108)
);

INVxp33_ASAP7_75t_L g1109 ( 
.A(n_1027),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1027),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1025),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1025),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_1045),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1036),
.B(n_281),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1036),
.B(n_136),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1049),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1031),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1019),
.B(n_142),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1053),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1034),
.B(n_148),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_1067),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_1091),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1066),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1085),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1112),
.Y(n_1125)
);

AND2x4_ASAP7_75t_SL g1126 ( 
.A(n_1088),
.B(n_1048),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1080),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1111),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1101),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1090),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1072),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1074),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1102),
.B(n_1057),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1075),
.B(n_1077),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1119),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1098),
.B(n_1057),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1087),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1068),
.B(n_1058),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1078),
.B(n_1057),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1107),
.B(n_1054),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1105),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1096),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1096),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1092),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1092),
.B(n_1055),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1090),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1081),
.A2(n_1044),
.B(n_1062),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1117),
.B(n_1069),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1113),
.Y(n_1149)
);

BUFx4f_ASAP7_75t_L g1150 ( 
.A(n_1069),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1086),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1108),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1079),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1105),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1089),
.A2(n_1062),
.B(n_1029),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1093),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1117),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1108),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1120),
.B(n_1056),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1094),
.B(n_1063),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1114),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1070),
.B(n_1050),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1114),
.B(n_1026),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1104),
.B(n_1042),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1076),
.B(n_1048),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1115),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1106),
.B(n_1052),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1118),
.B(n_149),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1084),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1099),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1099),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1082),
.B(n_155),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1129),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1129),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1156),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1136),
.B(n_1103),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1135),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1135),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1136),
.B(n_1104),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1122),
.B(n_1100),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_SL g1181 ( 
.A(n_1150),
.B(n_1110),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1145),
.B(n_1083),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1137),
.B(n_1097),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1145),
.B(n_1109),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1137),
.B(n_1071),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1121),
.B(n_1116),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_1127),
.B(n_1095),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1149),
.B(n_1146),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1161),
.B(n_1073),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1144),
.B(n_157),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1130),
.B(n_1151),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1123),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1164),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1132),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1134),
.B(n_1139),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1139),
.B(n_162),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1125),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1125),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1160),
.B(n_166),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1131),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1131),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1152),
.B(n_174),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1143),
.B(n_175),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1174),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1173),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1175),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1195),
.B(n_1170),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1188),
.B(n_1171),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1177),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1184),
.B(n_1142),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1193),
.B(n_1124),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1192),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1179),
.B(n_1165),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1193),
.B(n_1157),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1179),
.B(n_1165),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1178),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1189),
.B(n_1138),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1191),
.B(n_1133),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1182),
.B(n_1194),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1176),
.B(n_1158),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1176),
.B(n_1166),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1193),
.B(n_1157),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1187),
.B(n_1153),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1197),
.B(n_1147),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1205),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1218),
.B(n_1197),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_R g1227 ( 
.A1(n_1220),
.A2(n_1185),
.B(n_1180),
.C(n_1183),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1217),
.A2(n_1140),
.B1(n_1181),
.B2(n_1159),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1206),
.B(n_1186),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1204),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1208),
.B(n_1200),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1212),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1223),
.A2(n_1168),
.B(n_1190),
.C(n_1172),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1221),
.B(n_1201),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1211),
.B(n_1198),
.Y(n_1235)
);

OAI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_1227),
.A2(n_1213),
.B(n_1215),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1229),
.A2(n_1213),
.B1(n_1215),
.B2(n_1210),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1228),
.A2(n_1207),
.B1(n_1206),
.B2(n_1222),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1230),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1235),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1231),
.B(n_1219),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1233),
.A2(n_1214),
.B(n_1164),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_SL g1243 ( 
.A(n_1234),
.B(n_1196),
.C(n_1199),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1225),
.Y(n_1244)
);

NOR3xp33_ASAP7_75t_L g1245 ( 
.A(n_1232),
.B(n_1203),
.C(n_1202),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1226),
.A2(n_1206),
.B1(n_1163),
.B2(n_1162),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1242),
.A2(n_1164),
.B(n_1203),
.Y(n_1247)
);

AOI322xp5_ASAP7_75t_L g1248 ( 
.A1(n_1236),
.A2(n_1238),
.A3(n_1243),
.B1(n_1237),
.B2(n_1245),
.C1(n_1241),
.C2(n_1244),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1239),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1240),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1246),
.A2(n_1224),
.B(n_1148),
.C(n_1167),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1244),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1236),
.B(n_1209),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1248),
.B(n_1216),
.Y(n_1254)
);

NOR3x1_ASAP7_75t_L g1255 ( 
.A(n_1250),
.B(n_1253),
.C(n_1252),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1247),
.A2(n_1169),
.B(n_1155),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1254),
.B(n_1249),
.C(n_1251),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1255),
.Y(n_1258)
);

AOI211x1_ASAP7_75t_L g1259 ( 
.A1(n_1256),
.A2(n_1154),
.B(n_1141),
.C(n_1155),
.Y(n_1259)
);

NAND4xp25_ASAP7_75t_L g1260 ( 
.A(n_1258),
.B(n_1128),
.C(n_1126),
.D(n_182),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1259),
.A2(n_1154),
.B1(n_1141),
.B2(n_1126),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1257),
.A2(n_183),
.B(n_185),
.C(n_186),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1262),
.B(n_188),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1261),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1260),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1263),
.B(n_195),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1264),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_1265),
.B(n_201),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1267),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1266),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1268),
.Y(n_1271)
);

XNOR2xp5_ASAP7_75t_L g1272 ( 
.A(n_1271),
.B(n_1270),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1269),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1273),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1272),
.B(n_210),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1274),
.B(n_216),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1275),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1276),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1278),
.B(n_1277),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1278),
.B(n_236),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1279),
.A2(n_243),
.B1(n_248),
.B2(n_252),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1280),
.A2(n_254),
.B1(n_258),
.B2(n_260),
.Y(n_1282)
);

OR2x6_ASAP7_75t_L g1283 ( 
.A(n_1282),
.B(n_261),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1283),
.A2(n_1281),
.B1(n_268),
.B2(n_271),
.Y(n_1284)
);


endmodule