module fake_ariane_2827_n_611 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_611);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_611;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_261;
wire n_220;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_152;
wire n_405;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_115;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_108;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_588;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_102;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_606;
wire n_213;
wire n_110;
wire n_304;
wire n_583;
wire n_509;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_585;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_131;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_121;
wire n_118;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_116;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_127;
wire n_531;

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_0),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVxp33_ASAP7_75t_SL g110 ( 
.A(n_37),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_53),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_10),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_9),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_2),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_47),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_1),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_45),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_42),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_1),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_80),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_85),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_73),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_38),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_19),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_62),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_21),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_12),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_20),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_64),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_12),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_25),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_31),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_44),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_89),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_36),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_26),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_90),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_43),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_17),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_99),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_39),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_28),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_63),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_3),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_4),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_169),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_4),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_5),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_102),
.B(n_6),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_11),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_102),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_112),
.Y(n_234)
);

CKINVDCx6p67_ASAP7_75t_R g235 ( 
.A(n_192),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_143),
.B(n_22),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_103),
.A2(n_23),
.B(n_29),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

CKINVDCx8_ASAP7_75t_R g240 ( 
.A(n_104),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_116),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_105),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_108),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_32),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_109),
.B(n_35),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_109),
.B(n_123),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_120),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_149),
.B(n_46),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_106),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_172),
.B(n_83),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_120),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_133),
.A2(n_70),
.B1(n_82),
.B2(n_168),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_150),
.B(n_157),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_107),
.Y(n_264)
);

BUFx8_ASAP7_75t_L g265 ( 
.A(n_123),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_156),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_153),
.B(n_176),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_115),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_118),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_236),
.B(n_110),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_185),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_154),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_146),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_158),
.Y(n_279)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_159),
.B(n_187),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_211),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_239),
.B(n_179),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_193),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_239),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_195),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_206),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_101),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_224),
.B(n_122),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_219),
.B(n_194),
.Y(n_294)
);

BUFx6f_ASAP7_75t_SL g295 ( 
.A(n_237),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_219),
.A2(n_194),
.B1(n_168),
.B2(n_133),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_145),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_229),
.B(n_152),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_196),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_231),
.A2(n_130),
.B1(n_160),
.B2(n_179),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_208),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_138),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_196),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_235),
.B(n_136),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_210),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_200),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_190),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_222),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_221),
.B(n_132),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_228),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_200),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

NOR2x1p5_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_160),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_231),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_237),
.B1(n_207),
.B2(n_205),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_255),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_265),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_218),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_295),
.A2(n_225),
.B1(n_268),
.B2(n_207),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_262),
.B1(n_225),
.B2(n_254),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_309),
.B(n_240),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_255),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_285),
.B(n_240),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_301),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_234),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_271),
.Y(n_346)
);

OAI221xp5_ASAP7_75t_L g347 ( 
.A1(n_303),
.A2(n_267),
.B1(n_266),
.B2(n_269),
.C(n_233),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_225),
.B1(n_268),
.B2(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_295),
.A2(n_220),
.B1(n_218),
.B2(n_241),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_241),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_313),
.B(n_264),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_297),
.A2(n_242),
.B(n_245),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_313),
.B(n_234),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_220),
.B1(n_209),
.B2(n_201),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_199),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_199),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_198),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_288),
.B(n_198),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_197),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_292),
.B(n_201),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_197),
.Y(n_363)
);

NOR2x1_ASAP7_75t_R g364 ( 
.A(n_274),
.B(n_203),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_292),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_298),
.B(n_321),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_270),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_243),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_272),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_300),
.B(n_243),
.Y(n_371)
);

OR2x6_ASAP7_75t_L g372 ( 
.A(n_275),
.B(n_216),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_280),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_327),
.A2(n_294),
.B(n_324),
.C(n_318),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_280),
.B(n_305),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_280),
.B(n_305),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_296),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_326),
.A2(n_358),
.B(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_366),
.B(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_291),
.Y(n_382)
);

NOR2x1_ASAP7_75t_R g383 ( 
.A(n_354),
.B(n_291),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_341),
.B(n_324),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_324),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_319),
.B1(n_276),
.B2(n_284),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_347),
.A2(n_253),
.B1(n_223),
.B2(n_244),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_287),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_283),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_304),
.B(n_310),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_287),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_335),
.A2(n_314),
.B1(n_310),
.B2(n_141),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_348),
.A2(n_139),
.B1(n_166),
.B2(n_177),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_273),
.B(n_277),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_246),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_369),
.A2(n_281),
.B(n_289),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_371),
.A2(n_249),
.B(n_252),
.C(n_256),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_259),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_348),
.A2(n_140),
.B1(n_162),
.B2(n_173),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_337),
.A2(n_323),
.B(n_315),
.Y(n_407)
);

AND2x4_ASAP7_75t_SL g408 ( 
.A(n_368),
.B(n_217),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_367),
.B(n_257),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_250),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_329),
.B(n_250),
.Y(n_411)
);

O2A1O1Ixp5_ASAP7_75t_L g412 ( 
.A1(n_342),
.A2(n_322),
.B(n_249),
.C(n_184),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_364),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_331),
.B(n_263),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g417 ( 
.A1(n_346),
.A2(n_238),
.B(n_308),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_167),
.B1(n_128),
.B2(n_131),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_212),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_362),
.A2(n_113),
.B1(n_124),
.B2(n_127),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_332),
.B(n_250),
.Y(n_421)
);

AOI21xp33_ASAP7_75t_L g422 ( 
.A1(n_350),
.A2(n_355),
.B(n_373),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_368),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_352),
.B(n_129),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_345),
.A2(n_142),
.B1(n_151),
.B2(n_165),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_327),
.B(n_171),
.Y(n_427)
);

NOR3xp33_ASAP7_75t_L g428 ( 
.A(n_327),
.B(n_204),
.C(n_212),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_333),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_327),
.B(n_175),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_333),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_341),
.B(n_182),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_341),
.B(n_320),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_341),
.B(n_286),
.Y(n_435)
);

AOI221x1_ASAP7_75t_L g436 ( 
.A1(n_375),
.A2(n_374),
.B1(n_428),
.B2(n_376),
.C(n_407),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_312),
.B(n_202),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_230),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_230),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_230),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

AO31x2_ASAP7_75t_L g443 ( 
.A1(n_377),
.A2(n_202),
.A3(n_213),
.B(n_214),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_429),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_377),
.A2(n_202),
.A3(n_213),
.B(n_214),
.Y(n_445)
);

AO32x2_ASAP7_75t_L g446 ( 
.A1(n_398),
.A2(n_230),
.A3(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g447 ( 
.A1(n_382),
.A2(n_202),
.B1(n_213),
.B2(n_214),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_215),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_312),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_403),
.A2(n_392),
.B(n_400),
.Y(n_451)
);

AO21x1_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_435),
.B(n_403),
.Y(n_452)
);

O2A1O1Ixp33_ASAP7_75t_SL g453 ( 
.A1(n_416),
.A2(n_411),
.B(n_410),
.C(n_389),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_414),
.A2(n_434),
.B(n_404),
.C(n_406),
.Y(n_454)
);

BUFx12f_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_385),
.A2(n_388),
.B1(n_395),
.B2(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_409),
.B(n_423),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_R g460 ( 
.A(n_425),
.B(n_399),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_396),
.A2(n_424),
.B1(n_420),
.B2(n_386),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_422),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_412),
.A2(n_391),
.B(n_426),
.Y(n_466)
);

AO21x2_ASAP7_75t_L g467 ( 
.A1(n_418),
.A2(n_390),
.B(n_383),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_432),
.A2(n_327),
.B1(n_295),
.B2(n_301),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_432),
.A2(n_327),
.B1(n_295),
.B2(n_301),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_376),
.A2(n_379),
.B(n_374),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_333),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

AO31x2_ASAP7_75t_L g475 ( 
.A1(n_374),
.A2(n_376),
.A3(n_377),
.B(n_375),
.Y(n_475)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_378),
.A2(n_316),
.B1(n_296),
.B2(n_327),
.C(n_209),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_423),
.Y(n_477)
);

CKINVDCx11_ASAP7_75t_R g478 ( 
.A(n_431),
.Y(n_478)
);

BUFx2_ASAP7_75t_SL g479 ( 
.A(n_423),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_L g480 ( 
.A1(n_415),
.A2(n_327),
.B(n_339),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_376),
.A2(n_379),
.B(n_374),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_376),
.A2(n_379),
.B(n_374),
.Y(n_482)
);

O2A1O1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_415),
.A2(n_366),
.B(n_331),
.C(n_378),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_427),
.A2(n_295),
.B1(n_327),
.B2(n_378),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_376),
.A2(n_379),
.B(n_374),
.Y(n_485)
);

NOR3xp33_ASAP7_75t_L g486 ( 
.A(n_427),
.B(n_221),
.C(n_251),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_415),
.B(n_366),
.Y(n_487)
);

AO31x2_ASAP7_75t_L g488 ( 
.A1(n_374),
.A2(n_376),
.A3(n_377),
.B(n_375),
.Y(n_488)
);

AO21x2_ASAP7_75t_L g489 ( 
.A1(n_374),
.A2(n_376),
.B(n_417),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_384),
.A2(n_435),
.B(n_433),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_366),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

AO31x2_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_452),
.A3(n_490),
.B(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_472),
.A2(n_481),
.B(n_485),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_491),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_483),
.B(n_461),
.C(n_484),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_476),
.B(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_473),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_482),
.A2(n_489),
.B(n_451),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_442),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_469),
.B(n_470),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_478),
.Y(n_507)
);

AO31x2_ASAP7_75t_L g508 ( 
.A1(n_448),
.A2(n_454),
.A3(n_488),
.B(n_475),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_458),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_453),
.A2(n_449),
.B(n_466),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_467),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_439),
.A2(n_440),
.B(n_437),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_463),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_450),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_457),
.B(n_464),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_465),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_443),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_475),
.A2(n_488),
.B(n_460),
.C(n_446),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_446),
.A2(n_447),
.B(n_455),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_503),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_500),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_503),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_516),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g532 ( 
.A(n_506),
.B(n_495),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_501),
.Y(n_533)
);

BUFx8_ASAP7_75t_SL g534 ( 
.A(n_505),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_495),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_515),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_497),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_518),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_516),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_521),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_516),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_535),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_541),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_502),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_493),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_493),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_541),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_543),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_543),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_540),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_527),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_540),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_493),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_529),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_527),
.B(n_493),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_530),
.B(n_493),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_508),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_530),
.B(n_508),
.Y(n_564)
);

AND2x4_ASAP7_75t_SL g565 ( 
.A(n_554),
.B(n_531),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_555),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_538),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_545),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_538),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_560),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_533),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_534),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_539),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_547),
.Y(n_574)
);

NAND4xp25_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_520),
.C(n_507),
.D(n_533),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_571),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_570),
.B(n_562),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_566),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_558),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_565),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_568),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_572),
.B(n_548),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_573),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_576),
.Y(n_584)
);

AOI211xp5_ASAP7_75t_L g585 ( 
.A1(n_582),
.A2(n_575),
.B(n_572),
.C(n_573),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_548),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_580),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_581),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_577),
.Y(n_589)
);

AOI21xp33_ASAP7_75t_L g590 ( 
.A1(n_580),
.A2(n_551),
.B(n_552),
.Y(n_590)
);

NOR2x1_ASAP7_75t_L g591 ( 
.A(n_583),
.B(n_574),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_586),
.B(n_579),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_588),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_591),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_585),
.A2(n_558),
.B1(n_564),
.B2(n_565),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_594),
.A2(n_584),
.B(n_587),
.C(n_506),
.Y(n_596)
);

AOI222xp33_ASAP7_75t_L g597 ( 
.A1(n_596),
.A2(n_589),
.B1(n_593),
.B2(n_564),
.C1(n_578),
.C2(n_542),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_519),
.C(n_595),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_598),
.B(n_592),
.Y(n_599)
);

NAND4xp75_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_514),
.C(n_587),
.D(n_590),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_599),
.A2(n_562),
.B1(n_561),
.B2(n_547),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_601),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_600),
.B(n_588),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_603),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_604),
.A2(n_602),
.B1(n_563),
.B2(n_559),
.Y(n_605)
);

OAI211xp5_ASAP7_75t_SL g606 ( 
.A1(n_604),
.A2(n_556),
.B(n_510),
.C(n_522),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_605),
.A2(n_552),
.B1(n_553),
.B2(n_551),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_607),
.A2(n_606),
.B(n_524),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_513),
.B(n_524),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_609),
.A2(n_515),
.B(n_536),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_509),
.B1(n_532),
.B2(n_553),
.Y(n_611)
);


endmodule