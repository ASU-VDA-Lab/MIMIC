module fake_jpeg_29938_n_461 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_461);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_461;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_47),
.B(n_50),
.Y(n_138)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_51),
.B(n_59),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_29),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_58),
.B(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_0),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_65),
.B(n_67),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_18),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_33),
.A2(n_19),
.B1(n_40),
.B2(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_128)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_77),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_58),
.A2(n_27),
.B1(n_36),
.B2(n_38),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_27),
.B1(n_45),
.B2(n_43),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_112),
.A2(n_118),
.B1(n_119),
.B2(n_141),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_27),
.B1(n_45),
.B2(n_43),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_36),
.B1(n_38),
.B2(n_46),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_128),
.A2(n_134),
.B1(n_143),
.B2(n_149),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_36),
.B1(n_38),
.B2(n_26),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_36),
.B1(n_28),
.B2(n_39),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_42),
.B1(n_35),
.B2(n_25),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_68),
.A2(n_35),
.B1(n_25),
.B2(n_24),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_150),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_49),
.A2(n_24),
.B1(n_23),
.B2(n_36),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_71),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_72),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_55),
.B1(n_62),
.B2(n_70),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_52),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_53),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_61),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_155),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_130),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_69),
.C(n_47),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_173),
.C(n_112),
.Y(n_204)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_63),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_163),
.A2(n_183),
.B1(n_189),
.B2(n_192),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_103),
.B(n_75),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_165),
.B(n_168),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_80),
.B1(n_79),
.B2(n_56),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_103),
.B(n_57),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_170),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_48),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_89),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_171),
.B(n_174),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_111),
.B(n_76),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_87),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_142),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_178),
.B(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_185),
.Y(n_217)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_88),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_123),
.A2(n_84),
.B1(n_77),
.B2(n_85),
.Y(n_183)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_107),
.B(n_90),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_84),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_73),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_191),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_64),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_101),
.Y(n_192)
);

AND2x4_ASAP7_75t_SL g193 ( 
.A(n_107),
.B(n_1),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_194),
.Y(n_233)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_201),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_96),
.B(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_200),
.Y(n_246)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_5),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_96),
.B(n_5),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_150),
.A2(n_86),
.B1(n_83),
.B2(n_54),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_117),
.B1(n_133),
.B2(n_102),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_173),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_206),
.B1(n_213),
.B2(n_238),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_139),
.B1(n_116),
.B2(n_122),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_139),
.B1(n_116),
.B2(n_122),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_109),
.B(n_110),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_214),
.A2(n_152),
.B(n_177),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_113),
.B1(n_106),
.B2(n_97),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_216),
.A2(n_218),
.B1(n_227),
.B2(n_230),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_113),
.B1(n_125),
.B2(n_99),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_102),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_172),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_125),
.B1(n_99),
.B2(n_121),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_184),
.A2(n_121),
.B1(n_136),
.B2(n_117),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_188),
.A2(n_124),
.B1(n_6),
.B2(n_8),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_184),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_242),
.A2(n_243),
.B1(n_247),
.B2(n_156),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_200),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_238),
.B1(n_246),
.B2(n_241),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_10),
.B1(n_13),
.B2(n_155),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_174),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_248),
.B(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_151),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_250),
.B(n_256),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_153),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_259),
.C(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_221),
.B(n_160),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_257),
.B(n_262),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_261),
.B1(n_230),
.B2(n_218),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_185),
.C(n_173),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_158),
.B1(n_193),
.B2(n_198),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_210),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_191),
.B1(n_161),
.B2(n_197),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_277),
.B1(n_246),
.B2(n_208),
.Y(n_290)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_162),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_221),
.B(n_187),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_271),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_210),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_269),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_206),
.A2(n_179),
.B1(n_180),
.B2(n_157),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_270),
.A2(n_216),
.B1(n_227),
.B2(n_237),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_208),
.B(n_194),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_280),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_178),
.B(n_152),
.Y(n_276)
);

AOI22x1_ASAP7_75t_L g319 ( 
.A1(n_276),
.A2(n_283),
.B1(n_222),
.B2(n_215),
.Y(n_319)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_217),
.A2(n_159),
.B(n_172),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_176),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_154),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

OAI21x1_ASAP7_75t_SL g283 ( 
.A1(n_226),
.A2(n_189),
.B(n_195),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_175),
.C(n_189),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_231),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_225),
.B1(n_232),
.B2(n_223),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_289),
.A2(n_318),
.B1(n_235),
.B2(n_272),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_304),
.B1(n_270),
.B2(n_278),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_233),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_321),
.C(n_284),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_253),
.B(n_233),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_296),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_233),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_300),
.A2(n_306),
.B1(n_310),
.B2(n_275),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_213),
.B1(n_246),
.B2(n_225),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_254),
.A2(n_243),
.B1(n_245),
.B2(n_214),
.Y(n_310)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_205),
.A3(n_244),
.B1(n_236),
.B2(n_222),
.Y(n_316)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_276),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_317),
.B(n_319),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_257),
.A2(n_224),
.B1(n_215),
.B2(n_234),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_235),
.C(n_234),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_308),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_276),
.Y(n_324)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_291),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_291),
.C(n_296),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_326),
.B(n_327),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_299),
.A2(n_307),
.B(n_273),
.Y(n_327)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_224),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_335),
.Y(n_363)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_338),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_337),
.A2(n_344),
.B1(n_345),
.B2(n_307),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_298),
.Y(n_338)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_279),
.B(n_265),
.C(n_255),
.D(n_249),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_224),
.Y(n_375)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_341),
.A2(n_346),
.B1(n_348),
.B2(n_350),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_290),
.B(n_321),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_343),
.C(n_347),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_301),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_277),
.B1(n_254),
.B2(n_260),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_312),
.B(n_252),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_304),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_361),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_325),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_359),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_367),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_295),
.C(n_293),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_369),
.C(n_322),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_348),
.A2(n_306),
.B1(n_316),
.B2(n_320),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_358),
.A2(n_366),
.B1(n_324),
.B2(n_365),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_315),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_344),
.A2(n_320),
.B1(n_312),
.B2(n_313),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_345),
.A2(n_313),
.B1(n_315),
.B2(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_368),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_309),
.B1(n_308),
.B2(n_274),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_332),
.A2(n_264),
.B1(n_268),
.B2(n_269),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_282),
.C(n_285),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_262),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_375),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_379),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_328),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_328),
.C(n_349),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_389),
.C(n_394),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_381),
.A2(n_387),
.B1(n_396),
.B2(n_364),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_376),
.A2(n_349),
.B(n_337),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_393),
.B(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_330),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_386),
.B(n_392),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_358),
.A2(n_330),
.B1(n_339),
.B2(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_336),
.C(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_370),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_340),
.B(n_341),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_329),
.C(n_228),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g396 ( 
.A1(n_360),
.A2(n_329),
.B1(n_228),
.B2(n_13),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_397),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_373),
.B(n_382),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_408),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_359),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_410),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_397),
.A2(n_366),
.B1(n_351),
.B2(n_369),
.Y(n_406)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_409),
.A2(n_411),
.B1(n_401),
.B2(n_408),
.Y(n_428)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_375),
.B(n_351),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_384),
.B(n_383),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_391),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_395),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_353),
.C(n_352),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_389),
.C(n_384),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_414),
.C(n_403),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_409),
.A2(n_354),
.B1(n_391),
.B2(n_387),
.Y(n_417)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_398),
.B(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_424),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_385),
.C(n_377),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_404),
.C(n_403),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_402),
.B(n_416),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_413),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_428),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_415),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_407),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_431),
.B(n_399),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_438),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_433),
.A2(n_439),
.B(n_422),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_385),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_436),
.B(n_377),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_399),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_405),
.C(n_406),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_440),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_441),
.A2(n_447),
.B(n_439),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_428),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_445),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_435),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_446),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_419),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_442),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_450),
.C(n_437),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_440),
.C(n_416),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_454),
.A2(n_455),
.B(n_431),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_456),
.A2(n_457),
.B(n_429),
.Y(n_458)
);

OAI311xp33_ASAP7_75t_L g459 ( 
.A1(n_458),
.A2(n_451),
.A3(n_427),
.B1(n_436),
.C1(n_407),
.Y(n_459)
);

NAND5xp2_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_427),
.C(n_410),
.D(n_379),
.E(n_13),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_13),
.Y(n_461)
);


endmodule