module fake_ariane_1900_n_1184 (n_295, n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_289, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_294, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_299, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_291, n_20, n_292, n_174, n_275, n_100, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_297, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_290, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_293, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_14, n_163, n_88, n_186, n_141, n_296, n_298, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1184);

input n_295;
input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_289;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_294;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_299;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_291;
input n_20;
input n_292;
input n_174;
input n_275;
input n_100;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_297;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_290;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_293;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_296;
input n_298;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1184;

wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_479;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_1167;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_1154;
wire n_1166;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_1181;
wire n_445;
wire n_515;
wire n_379;
wire n_807;
wire n_765;
wire n_1131;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_336;
wire n_665;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_402;
wire n_1068;
wire n_1052;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_433;
wire n_600;
wire n_721;
wire n_795;
wire n_481;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_1153;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_1172;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_1160;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1085;
wire n_467;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_538;
wire n_352;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_654;
wire n_429;
wire n_455;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_459;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_617;
wire n_658;
wire n_705;
wire n_630;
wire n_616;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_673;
wire n_452;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_680;
wire n_571;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_1164;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_746;
wire n_456;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_615;
wire n_1070;
wire n_1027;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_739;
wire n_496;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_782;
wire n_650;
wire n_364;
wire n_856;
wire n_477;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1071;
wire n_484;
wire n_712;
wire n_411;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_797;
wire n_382;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_187),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_221),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_284),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_253),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_66),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_238),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_214),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_165),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_139),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_76),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_228),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_145),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_55),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_182),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_83),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_279),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_213),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_120),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_46),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_36),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_217),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_74),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_51),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_63),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_201),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_71),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_33),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_9),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_108),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_4),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_170),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_38),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_193),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_70),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_195),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_242),
.Y(n_350)
);

BUFx2_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_116),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_152),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_202),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_207),
.Y(n_355)
);

BUFx2_ASAP7_75t_R g356 ( 
.A(n_282),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_235),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_59),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_97),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_209),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_173),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_289),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_192),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_237),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_131),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_273),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_122),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_197),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_162),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_295),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_250),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_138),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_107),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_64),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_218),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_43),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_24),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_49),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_277),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_147),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_81),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_115),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_130),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_151),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_291),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_168),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_75),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_9),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_296),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_290),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_16),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_41),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_257),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_136),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_144),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_21),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_18),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_247),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_88),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_100),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_278),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_98),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_203),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_243),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_18),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_175),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_206),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_45),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_188),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_32),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_263),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_31),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_177),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_93),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_181),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_223),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_0),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_106),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_15),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_244),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_270),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_25),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_4),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_231),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_77),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_174),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_2),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_184),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_68),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_272),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_7),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_1),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_61),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_0),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_156),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_266),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_163),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_89),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_56),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_142),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_30),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_215),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_112),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_210),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_232),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_189),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_121),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_62),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_15),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_260),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_252),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_154),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_176),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_211),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_258),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_204),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_8),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_58),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_183),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_262),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_123),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_17),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_72),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_198),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_109),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_133),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_269),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_226),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_135),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_134),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_78),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_67),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_111),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_196),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_161),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_50),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_95),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_27),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_16),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_294),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_159),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_280),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_101),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_87),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_40),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_82),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_286),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_239),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_212),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_42),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_153),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_219),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_172),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_149),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_180),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g500 ( 
.A(n_65),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_234),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_370),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_328),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_337),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_370),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_346),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_409),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_395),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_340),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_362),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_433),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_444),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_344),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_460),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_484),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_436),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_345),
.B(n_1),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_392),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_483),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_385),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_472),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_373),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_431),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_438),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_397),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_453),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_461),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_500),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_402),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_347),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_466),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_442),
.B(n_2),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_300),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_302),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_301),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_306),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_426),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_442),
.B(n_3),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_309),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_312),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_351),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_313),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_315),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_319),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_338),
.B(n_3),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_339),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_341),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_354),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_303),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_358),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_359),
.B(n_5),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_361),
.B(n_5),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_304),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_356),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_368),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_305),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_308),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_307),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_375),
.B(n_6),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_376),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_320),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_329),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_499),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_377),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_398),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_428),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_355),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_311),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_388),
.B(n_6),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_314),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_390),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_391),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_412),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_318),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_414),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_322),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_323),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_325),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_326),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_500),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_432),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_327),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_330),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_501),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_437),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_441),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_331),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_443),
.B(n_7),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_445),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_R g600 ( 
.A(n_332),
.B(n_22),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_355),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_333),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_334),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_446),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_447),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_448),
.Y(n_606)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_335),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_449),
.B(n_8),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_336),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_342),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_348),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_450),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_349),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_350),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_534),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_534),
.B(n_355),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_576),
.B(n_451),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_589),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_589),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_546),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_544),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_510),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_513),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_545),
.B(n_316),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_540),
.B(n_400),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_541),
.B(n_439),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_521),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_519),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_601),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_566),
.B(n_457),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_458),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_548),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_570),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_550),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_310),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_557),
.B(n_324),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_561),
.B(n_360),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_554),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_555),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_556),
.Y(n_647)
);

OA21x2_ASAP7_75t_L g648 ( 
.A1(n_553),
.A2(n_578),
.B(n_560),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_558),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_563),
.B(n_355),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_568),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_564),
.B(n_465),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_573),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_542),
.B(n_317),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_590),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_591),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_595),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_503),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_596),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_604),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_605),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

NOR2x1_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_321),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_531),
.B(n_343),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_606),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_516),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_599),
.A2(n_468),
.B(n_467),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_565),
.B(n_469),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_538),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_559),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_502),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_567),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_369),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_504),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_522),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_506),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_505),
.A2(n_476),
.B(n_473),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_526),
.A2(n_489),
.B(n_480),
.Y(n_689)
);

BUFx12f_ASAP7_75t_L g690 ( 
.A(n_512),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_543),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_577),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_562),
.B(n_365),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_579),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_583),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_532),
.B(n_393),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_585),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_600),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_600),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_545),
.B(n_417),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_586),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_587),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_632),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_615),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_632),
.B(n_574),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_641),
.B(n_655),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_677),
.B(n_575),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g708 ( 
.A(n_690),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_698),
.B(n_588),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_698),
.B(n_699),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_668),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_699),
.B(n_607),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_676),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_624),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_676),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_669),
.B(n_592),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_625),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_622),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_696),
.B(n_593),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_669),
.B(n_597),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_619),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_694),
.B(n_509),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_683),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_686),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_615),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_623),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_676),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_661),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_638),
.B(n_533),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_623),
.Y(n_732)
);

INVx6_ASAP7_75t_L g733 ( 
.A(n_668),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_680),
.B(n_594),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_618),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_692),
.B(n_417),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_668),
.Y(n_737)
);

INVx4_ASAP7_75t_SL g738 ( 
.A(n_650),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_691),
.B(n_602),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_651),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_651),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_657),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

INVx4_ASAP7_75t_SL g745 ( 
.A(n_650),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_618),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_657),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_688),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_640),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_672),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_633),
.B(n_549),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_689),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_682),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_626),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_537),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_671),
.B(n_508),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_669),
.B(n_609),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_636),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_640),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_685),
.A2(n_613),
.B1(n_614),
.B2(n_603),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_673),
.B(n_536),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_637),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_670),
.B(n_518),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_645),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_656),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_654),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_695),
.B(n_610),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_675),
.B(n_611),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_656),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_617),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_675),
.B(n_571),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_639),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_662),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_697),
.B(n_701),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_675),
.B(n_527),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_664),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_642),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_702),
.B(n_511),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_621),
.B(n_507),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_653),
.B(n_535),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_646),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_647),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_674),
.B(n_515),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_649),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_652),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_725),
.B(n_520),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_708),
.B(n_693),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_726),
.B(n_685),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_704),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_730),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_705),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_755),
.B(n_753),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_707),
.Y(n_794)
);

AO22x2_ASAP7_75t_L g795 ( 
.A1(n_760),
.A2(n_687),
.B1(n_681),
.B2(n_684),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_743),
.B(n_621),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_705),
.B(n_703),
.Y(n_797)
);

AO22x2_ASAP7_75t_L g798 ( 
.A1(n_707),
.A2(n_523),
.B1(n_687),
.B2(n_681),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_731),
.B(n_621),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_734),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_710),
.B(n_648),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_704),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_737),
.B(n_630),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_775),
.A2(n_648),
.B1(n_629),
.B2(n_628),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_733),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_735),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_735),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_709),
.A2(n_700),
.B1(n_627),
.B2(n_644),
.Y(n_808)
);

AO22x2_ASAP7_75t_L g809 ( 
.A1(n_734),
.A2(n_684),
.B1(n_679),
.B2(n_678),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_728),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_770),
.B(n_634),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_712),
.B(n_635),
.Y(n_813)
);

AO22x2_ASAP7_75t_L g814 ( 
.A1(n_739),
.A2(n_679),
.B1(n_643),
.B2(n_659),
.Y(n_814)
);

AO22x2_ASAP7_75t_L g815 ( 
.A1(n_761),
.A2(n_658),
.B1(n_660),
.B2(n_665),
.Y(n_815)
);

OAI221xp5_ASAP7_75t_L g816 ( 
.A1(n_706),
.A2(n_663),
.B1(n_666),
.B2(n_667),
.C(n_498),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_778),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_778),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_780),
.B(n_650),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_716),
.B(n_616),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_763),
.B(n_384),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_727),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_739),
.A2(n_422),
.B1(n_482),
.B2(n_493),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_713),
.B(n_417),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_780),
.B(n_10),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_784),
.B(n_10),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_746),
.Y(n_827)
);

OAI221xp5_ASAP7_75t_L g828 ( 
.A1(n_754),
.A2(n_786),
.B1(n_785),
.B2(n_783),
.C(n_782),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_758),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_763),
.B(n_417),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_773),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_711),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_764),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_781),
.B(n_11),
.Y(n_835)
);

AOI22x1_ASAP7_75t_L g836 ( 
.A1(n_765),
.A2(n_420),
.B1(n_353),
.B2(n_357),
.Y(n_836)
);

AO22x2_ASAP7_75t_L g837 ( 
.A1(n_776),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_756),
.Y(n_838)
);

AO22x2_ASAP7_75t_L g839 ( 
.A1(n_771),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_721),
.A2(n_425),
.B1(n_363),
.B2(n_364),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_779),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_767),
.A2(n_429),
.B1(n_366),
.B2(n_367),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_766),
.Y(n_843)
);

OR2x2_ASAP7_75t_SL g844 ( 
.A(n_733),
.B(n_495),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_774),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_715),
.B(n_495),
.Y(n_846)
);

NAND2x1p5_ASAP7_75t_L g847 ( 
.A(n_729),
.B(n_495),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_769),
.B(n_650),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_717),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_779),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_768),
.Y(n_851)
);

AO22x2_ASAP7_75t_L g852 ( 
.A1(n_720),
.A2(n_751),
.B1(n_718),
.B2(n_714),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_719),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_724),
.B(n_772),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_749),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_722),
.B(n_495),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_759),
.A2(n_440),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_751),
.B(n_616),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_757),
.B(n_352),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_723),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_742),
.A2(n_747),
.B1(n_740),
.B2(n_741),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_777),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_744),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_744),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_736),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_736),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_791),
.B(n_752),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_854),
.B(n_752),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_SL g869 ( 
.A(n_835),
.B(n_748),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_813),
.B(n_811),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_789),
.B(n_799),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_851),
.B(n_748),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_826),
.B(n_750),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_793),
.B(n_750),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_804),
.B(n_738),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_SL g876 ( 
.A(n_796),
.B(n_378),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_808),
.B(n_738),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_817),
.B(n_736),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_SL g879 ( 
.A(n_818),
.B(n_379),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_797),
.B(n_745),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_859),
.B(n_745),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_855),
.B(n_380),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_825),
.B(n_381),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_819),
.B(n_382),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_SL g885 ( 
.A(n_829),
.B(n_383),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_842),
.B(n_387),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_831),
.B(n_389),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_SL g888 ( 
.A(n_810),
.B(n_394),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_790),
.B(n_802),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_806),
.B(n_396),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_807),
.B(n_399),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_812),
.B(n_403),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_840),
.B(n_404),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_787),
.B(n_19),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_861),
.B(n_864),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_863),
.B(n_405),
.Y(n_896)
);

NAND2xp33_ASAP7_75t_SL g897 ( 
.A(n_848),
.B(n_833),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_858),
.B(n_406),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_788),
.B(n_407),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_SL g900 ( 
.A(n_805),
.B(n_408),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_792),
.B(n_410),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_803),
.B(n_411),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_SL g903 ( 
.A(n_801),
.B(n_413),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_SL g904 ( 
.A(n_822),
.B(n_415),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_794),
.B(n_616),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_827),
.B(n_616),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_836),
.B(n_416),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_800),
.B(n_418),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_832),
.B(n_419),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_865),
.B(n_424),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_830),
.B(n_20),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_866),
.B(n_434),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_838),
.B(n_452),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_841),
.B(n_454),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_834),
.B(n_455),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_843),
.B(n_456),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_830),
.B(n_20),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_845),
.B(n_459),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_850),
.B(n_462),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_849),
.B(n_463),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_853),
.B(n_464),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_815),
.B(n_470),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_860),
.B(n_824),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_846),
.B(n_471),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_847),
.B(n_474),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_870),
.B(n_795),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_875),
.A2(n_856),
.B(n_820),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_889),
.A2(n_828),
.B(n_857),
.Y(n_928)
);

OAI21x1_ASAP7_75t_SL g929 ( 
.A1(n_878),
.A2(n_862),
.B(n_837),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_873),
.A2(n_862),
.B(n_816),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_871),
.B(n_795),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_906),
.A2(n_814),
.B(n_809),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_895),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_SL g934 ( 
.A1(n_911),
.A2(n_837),
.B(n_839),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_899),
.B(n_821),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_L g936 ( 
.A(n_869),
.B(n_814),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_903),
.A2(n_809),
.B(n_852),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_874),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_868),
.A2(n_923),
.B(n_881),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_872),
.A2(n_500),
.B(n_844),
.Y(n_940)
);

AO31x2_ASAP7_75t_L g941 ( 
.A1(n_909),
.A2(n_823),
.A3(n_798),
.B(n_500),
.Y(n_941)
);

NAND2x1_ASAP7_75t_L g942 ( 
.A(n_905),
.B(n_821),
.Y(n_942)
);

AOI221x1_ASAP7_75t_L g943 ( 
.A1(n_897),
.A2(n_823),
.B1(n_500),
.B2(n_496),
.C(n_494),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_907),
.A2(n_486),
.B(n_492),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_905),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_880),
.B(n_911),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_902),
.B(n_475),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_917),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_917),
.B(n_477),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_920),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_894),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_922),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_879),
.A2(n_487),
.B(n_491),
.C(n_490),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_877),
.A2(n_500),
.B(n_26),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_884),
.Y(n_955)
);

BUFx4_ASAP7_75t_SL g956 ( 
.A(n_913),
.Y(n_956)
);

AO31x2_ASAP7_75t_L g957 ( 
.A1(n_890),
.A2(n_23),
.A3(n_29),
.B(n_35),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_867),
.A2(n_37),
.B(n_39),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_901),
.B(n_478),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_891),
.A2(n_488),
.B(n_485),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_892),
.A2(n_481),
.B(n_479),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_883),
.B(n_44),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_SL g963 ( 
.A1(n_893),
.A2(n_47),
.B(n_48),
.C(n_52),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_919),
.B(n_53),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_915),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_885),
.B(n_54),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_888),
.B(n_908),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_887),
.A2(n_57),
.B(n_60),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_900),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_886),
.A2(n_69),
.B(n_73),
.Y(n_970)
);

CKINVDCx8_ASAP7_75t_R g971 ( 
.A(n_946),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_956),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_948),
.B(n_914),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_927),
.A2(n_925),
.B(n_924),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_951),
.B(n_898),
.Y(n_975)
);

AOI21x1_ASAP7_75t_L g976 ( 
.A1(n_930),
.A2(n_921),
.B(n_918),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_938),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_926),
.A2(n_916),
.B(n_896),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_928),
.A2(n_876),
.B(n_904),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_946),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_933),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_939),
.A2(n_882),
.B(n_910),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_952),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_936),
.A2(n_912),
.B1(n_80),
.B2(n_84),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_931),
.B(n_79),
.Y(n_985)
);

AO32x2_ASAP7_75t_L g986 ( 
.A1(n_934),
.A2(n_85),
.A3(n_86),
.B1(n_90),
.B2(n_92),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_963),
.A2(n_94),
.B(n_96),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_958),
.A2(n_99),
.B(n_102),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_937),
.A2(n_103),
.B(n_104),
.Y(n_989)
);

OAI21x1_ASAP7_75t_SL g990 ( 
.A1(n_929),
.A2(n_105),
.B(n_110),
.Y(n_990)
);

AO31x2_ASAP7_75t_L g991 ( 
.A1(n_943),
.A2(n_113),
.A3(n_114),
.B(n_117),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_932),
.A2(n_118),
.B(n_119),
.Y(n_992)
);

OA21x2_ASAP7_75t_L g993 ( 
.A1(n_970),
.A2(n_124),
.B(n_125),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_968),
.A2(n_126),
.B(n_127),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_940),
.A2(n_128),
.B(n_129),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_950),
.A2(n_132),
.B(n_137),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_935),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_997)
);

OAI221xp5_ASAP7_75t_L g998 ( 
.A1(n_955),
.A2(n_299),
.B1(n_148),
.B2(n_150),
.C(n_155),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_942),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_969),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_945),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_945),
.Y(n_1002)
);

AO31x2_ASAP7_75t_L g1003 ( 
.A1(n_962),
.A2(n_146),
.A3(n_157),
.B(n_158),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_965),
.A2(n_164),
.B1(n_169),
.B2(n_178),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_945),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_967),
.B(n_297),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_949),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_947),
.A2(n_179),
.B1(n_185),
.B2(n_186),
.Y(n_1008)
);

OA21x2_ASAP7_75t_L g1009 ( 
.A1(n_987),
.A2(n_944),
.B(n_966),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_972),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_977),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_981),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_975),
.B(n_941),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_992),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1005),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_992),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_990),
.B(n_964),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_983),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_980),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_985),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1007),
.B(n_941),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1007),
.B(n_941),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_978),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_1002),
.B(n_954),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_995),
.A2(n_988),
.B(n_974),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1003),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1003),
.Y(n_1027)
);

AO21x2_ASAP7_75t_L g1028 ( 
.A1(n_990),
.A2(n_953),
.B(n_960),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_978),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_1001),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_982),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_976),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_976),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_986),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_986),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_979),
.B(n_957),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_999),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_989),
.B(n_959),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_1000),
.B(n_973),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_996),
.A2(n_961),
.B1(n_957),
.B2(n_194),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_986),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1006),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_971),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_997),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1006),
.B(n_957),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1003),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1011),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1012),
.Y(n_1049)
);

XNOR2xp5_ASAP7_75t_L g1050 ( 
.A(n_1018),
.B(n_984),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1020),
.B(n_991),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_R g1052 ( 
.A(n_1017),
.B(n_994),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_1010),
.Y(n_1053)
);

OR2x4_ASAP7_75t_L g1054 ( 
.A(n_1043),
.B(n_991),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_1037),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_1018),
.B(n_1008),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1030),
.B(n_998),
.Y(n_1057)
);

XOR2xp5_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_1004),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_R g1059 ( 
.A(n_1017),
.B(n_994),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_1043),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1013),
.B(n_991),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1042),
.B(n_993),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_1017),
.B(n_993),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1022),
.B(n_190),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_1019),
.Y(n_1065)
);

XOR2xp5_ASAP7_75t_L g1066 ( 
.A(n_1044),
.B(n_191),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_R g1067 ( 
.A(n_1030),
.B(n_199),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_1021),
.B(n_200),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1015),
.B(n_205),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1024),
.B(n_208),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1034),
.B(n_216),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_1044),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1035),
.B(n_220),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_1045),
.B(n_1041),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_1036),
.B(n_222),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1038),
.B(n_224),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_1036),
.B(n_227),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_1038),
.B(n_229),
.Y(n_1078)
);

CKINVDCx11_ASAP7_75t_R g1079 ( 
.A(n_1038),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_1040),
.B(n_1028),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1029),
.B(n_230),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_1024),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1053),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_1028),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1048),
.B(n_1023),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1049),
.B(n_1029),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1051),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1047),
.B(n_1033),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1065),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_1032),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_1031),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1070),
.B(n_1046),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1061),
.B(n_1027),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1055),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_L g1095 ( 
.A(n_1057),
.B(n_1027),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1079),
.B(n_1026),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1071),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1073),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1081),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1064),
.B(n_1026),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1078),
.A2(n_1040),
.B1(n_1009),
.B2(n_1016),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1054),
.Y(n_1102)
);

AND2x4_ASAP7_75t_SL g1103 ( 
.A(n_1072),
.B(n_1016),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1062),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1076),
.B(n_1014),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1068),
.Y(n_1106)
);

AND2x4_ASAP7_75t_SL g1107 ( 
.A(n_1070),
.B(n_1014),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1101),
.A2(n_1078),
.B1(n_1050),
.B2(n_1063),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1085),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1090),
.B(n_1103),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_1104),
.B(n_1087),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1091),
.B(n_1056),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1083),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1088),
.B(n_1063),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1088),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1086),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1085),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1096),
.B(n_1077),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1086),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1109),
.B(n_1102),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1116),
.Y(n_1121)
);

NAND3x1_ASAP7_75t_L g1122 ( 
.A(n_1112),
.B(n_1094),
.C(n_1089),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1119),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1111),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1110),
.B(n_1104),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1115),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1114),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1111),
.B(n_1087),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1122),
.A2(n_1108),
.B1(n_1067),
.B2(n_1052),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1126),
.B(n_1097),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1121),
.B(n_1098),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1128),
.Y(n_1133)
);

AO221x2_ASAP7_75t_L g1134 ( 
.A1(n_1123),
.A2(n_1108),
.B1(n_1113),
.B2(n_1066),
.C(n_1058),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_1120),
.B(n_1113),
.Y(n_1135)
);

NOR4xp25_ASAP7_75t_SL g1136 ( 
.A(n_1124),
.B(n_1059),
.C(n_1080),
.D(n_1106),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1131),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1132),
.B(n_1125),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_1133),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1134),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1135),
.B(n_1124),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1130),
.B(n_1127),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1136),
.B(n_1127),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1133),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1131),
.B(n_1129),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1133),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1138),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1140),
.A2(n_1118),
.B(n_1095),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1144),
.B(n_1084),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1140),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1139),
.B(n_1068),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1141),
.B(n_1107),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1147),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1151),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1149),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_SL g1156 ( 
.A1(n_1150),
.A2(n_1152),
.B(n_1146),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1148),
.B(n_1143),
.C(n_1142),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1149),
.B(n_1137),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1153),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1155),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1158),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_1145),
.Y(n_1162)
);

NAND4xp75_ASAP7_75t_L g1163 ( 
.A(n_1160),
.B(n_1156),
.C(n_1157),
.D(n_1069),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1161),
.B(n_1105),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1159),
.B(n_1105),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_1162),
.B(n_1092),
.C(n_1093),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_1075),
.B1(n_1093),
.B2(n_1092),
.C(n_1100),
.Y(n_1167)
);

AOI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1163),
.A2(n_1025),
.B(n_1009),
.C(n_241),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1166),
.B(n_233),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1168),
.B(n_240),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1170),
.B(n_1167),
.Y(n_1171)
);

XOR2xp5_ASAP7_75t_L g1172 ( 
.A(n_1171),
.B(n_1169),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1171),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1173),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1172),
.B(n_245),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1174),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1175),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1174),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1177),
.A2(n_251),
.B1(n_254),
.B2(n_256),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1179),
.A2(n_1178),
.B(n_1176),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1180),
.B(n_259),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1181),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1182),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.C(n_267),
.Y(n_1183)
);

AOI211xp5_ASAP7_75t_L g1184 ( 
.A1(n_1183),
.A2(n_268),
.B(n_271),
.C(n_274),
.Y(n_1184)
);


endmodule