module fake_jpeg_29697_n_478 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_478);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_478;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_51),
.B(n_67),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_53),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_12),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_64),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_12),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_12),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_76),
.Y(n_134)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_10),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_78),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_0),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_94),
.Y(n_122)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_1),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_1),
.C(n_2),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_90),
.Y(n_142)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_91),
.B(n_92),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_97),
.B1(n_26),
.B2(n_94),
.Y(n_100)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_19),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_100),
.A2(n_108),
.B(n_112),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_32),
.B1(n_46),
.B2(n_41),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_106),
.A2(n_110),
.B1(n_63),
.B2(n_89),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_21),
.B1(n_26),
.B2(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_46),
.B1(n_41),
.B2(n_32),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_79),
.B1(n_91),
.B2(n_84),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_46),
.B1(n_41),
.B2(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_41),
.B1(n_46),
.B2(n_44),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_48),
.B1(n_45),
.B2(n_38),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_138),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_121),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_27),
.B1(n_44),
.B2(n_31),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_52),
.B(n_23),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_128),
.B(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_31),
.B1(n_42),
.B2(n_40),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_50),
.A2(n_23),
.B1(n_42),
.B2(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_19),
.B1(n_45),
.B2(n_38),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_80),
.B(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_53),
.B(n_28),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_62),
.A2(n_28),
.B1(n_48),
.B2(n_18),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_22),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_59),
.B(n_35),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_71),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_190),
.C(n_119),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_156),
.B(n_186),
.Y(n_232)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_158),
.Y(n_230)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_71),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_162),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_86),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_35),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_167),
.Y(n_224)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_35),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_22),
.B1(n_82),
.B2(n_93),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_176),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

CKINVDCx6p67_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_173),
.B1(n_175),
.B2(n_198),
.Y(n_210)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_114),
.A2(n_65),
.B1(n_22),
.B2(n_7),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_4),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_105),
.B1(n_131),
.B2(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_116),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_182),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_4),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_124),
.A2(n_113),
.B1(n_115),
.B2(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_192),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_113),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_8),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_197),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_136),
.B1(n_137),
.B2(n_147),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_8),
.B(n_9),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_193),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_9),
.B1(n_150),
.B2(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_9),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_9),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_117),
.A2(n_128),
.B1(n_143),
.B2(n_127),
.Y(n_198)
);

OR2x4_ASAP7_75t_L g199 ( 
.A(n_120),
.B(n_138),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_201),
.B(n_102),
.Y(n_237)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_135),
.A2(n_150),
.B1(n_133),
.B2(n_105),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_142),
.B(n_138),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_154),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_231),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_146),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_214),
.A2(n_190),
.B(n_157),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_110),
.B1(n_101),
.B2(n_145),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_219),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_155),
.A2(n_145),
.B1(n_106),
.B2(n_149),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_105),
.B1(n_131),
.B2(n_125),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_227),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_119),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_161),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_244),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_182),
.B(n_168),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_196),
.B(n_105),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_155),
.B(n_189),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_155),
.A2(n_111),
.B1(n_131),
.B2(n_189),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_243),
.A2(n_174),
.B1(n_199),
.B2(n_203),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_162),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_167),
.B(n_111),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_161),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_111),
.C(n_131),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_247),
.Y(n_299)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_258),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_205),
.B(n_216),
.Y(n_286)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_256),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_189),
.B1(n_174),
.B2(n_157),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_262),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_221),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_259),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_270),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_197),
.B(n_177),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_273),
.B(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_187),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_264),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_157),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_174),
.B1(n_154),
.B2(n_170),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_269),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_176),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_204),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_274),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_182),
.B(n_193),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_176),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_160),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_246),
.C(n_232),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_206),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_283),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_186),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_156),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_216),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_153),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_242),
.B(n_153),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_158),
.B(n_111),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_285),
.B(n_170),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_288),
.B(n_295),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_287),
.B(n_309),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_214),
.B(n_222),
.C(n_210),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_289),
.B(n_250),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_211),
.C(n_207),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_307),
.C(n_311),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_215),
.B1(n_230),
.B2(n_170),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_300),
.B1(n_236),
.B2(n_247),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_219),
.B(n_218),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_213),
.B1(n_218),
.B2(n_228),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_236),
.B(n_208),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_251),
.B(n_274),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_207),
.C(n_178),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_230),
.C(n_213),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_254),
.B(n_200),
.C(n_206),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_164),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_314),
.C(n_317),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_159),
.C(n_234),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_170),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_317),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_320),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_319),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_321),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_296),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_322),
.A2(n_348),
.B1(n_313),
.B2(n_314),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_257),
.B1(n_303),
.B2(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_327),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_263),
.Y(n_325)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_331),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_330),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_271),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_271),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

NOR3xp33_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_283),
.C(n_267),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_334),
.B(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_251),
.Y(n_335)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_276),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_337),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_296),
.A2(n_273),
.B(n_267),
.C(n_276),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_338),
.A2(n_346),
.B1(n_297),
.B2(n_292),
.Y(n_372)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_344),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_284),
.C(n_279),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_307),
.C(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_303),
.A2(n_255),
.B1(n_250),
.B2(n_253),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_270),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_306),
.A2(n_286),
.B1(n_305),
.B2(n_315),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_229),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_229),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_350),
.Y(n_355)
);

INVx13_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_351),
.B(n_309),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_308),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_354),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_308),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_373),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_323),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_304),
.B1(n_289),
.B2(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_311),
.Y(n_363)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_367),
.C(n_342),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_312),
.C(n_302),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_343),
.B(n_302),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_370),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_297),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_346),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_266),
.Y(n_373)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_292),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_322),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_381),
.Y(n_412)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_382),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_362),
.Y(n_381)
);

BUFx12_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_390),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_SL g384 ( 
.A(n_366),
.B(n_330),
.C(n_337),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_384),
.B(n_399),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_389),
.C(n_365),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_324),
.C(n_329),
.Y(n_389)
);

FAx1_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_324),
.CI(n_337),
.CON(n_390),
.SN(n_390)
);

BUFx12_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_396),
.B(n_354),
.Y(n_406)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_331),
.Y(n_398)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_400),
.B(n_401),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_339),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_404),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_357),
.B(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_403),
.B(n_393),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_373),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_352),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_406),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_367),
.C(n_356),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_417),
.C(n_395),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_357),
.B(n_371),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_416),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_378),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_396),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_387),
.A2(n_377),
.B1(n_338),
.B2(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_369),
.C(n_345),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_434),
.C(n_405),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_425),
.A2(n_412),
.B(n_403),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_402),
.C(n_404),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_430),
.C(n_433),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_427),
.A2(n_397),
.B1(n_340),
.B2(n_333),
.Y(n_444)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_429),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_420),
.B(n_388),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_395),
.C(n_386),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_431),
.B(n_435),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_432),
.A2(n_414),
.B(n_422),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_390),
.C(n_394),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_413),
.A2(n_384),
.B1(n_359),
.B2(n_391),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_423),
.Y(n_453)
);

AOI21xp33_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_407),
.B(n_418),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_445),
.B(n_448),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_407),
.C(n_406),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_421),
.C(n_424),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_426),
.A2(n_409),
.B(n_380),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_444),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_432),
.A2(n_391),
.B(n_338),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_423),
.A2(n_338),
.B1(n_299),
.B2(n_336),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_SL g448 ( 
.A(n_424),
.B(n_382),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_445),
.A2(n_338),
.B(n_382),
.C(n_344),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_247),
.B(n_209),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_459),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_454),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_277),
.C(n_272),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_440),
.B(n_248),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_455),
.B(n_459),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_350),
.B(n_248),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_458),
.A2(n_172),
.B(n_169),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_235),
.C(n_194),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_446),
.A3(n_438),
.B1(n_228),
.B2(n_194),
.C1(n_209),
.C2(n_163),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_464),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_158),
.A3(n_163),
.B1(n_169),
.B2(n_172),
.C1(n_235),
.C2(n_451),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_466),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_450),
.A2(n_452),
.B(n_454),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_457),
.C(n_462),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_468),
.B(n_469),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_457),
.C(n_460),
.Y(n_469)
);

OA21x2_ASAP7_75t_SL g474 ( 
.A1(n_468),
.A2(n_471),
.B(n_470),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_474),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_472),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_475),
.B(n_473),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_R g478 ( 
.A(n_477),
.B(n_476),
.Y(n_478)
);


endmodule