module real_aes_2162_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_0), .B(n_131), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_1), .A2(n_31), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_1), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_2), .A2(n_140), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_3), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_4), .B(n_131), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_5), .B(n_147), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_6), .B(n_147), .Y(n_539) );
INVx1_ASAP7_75t_L g138 ( .A(n_7), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_8), .B(n_147), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_9), .Y(n_764) );
NAND2xp33_ASAP7_75t_L g516 ( .A(n_10), .B(n_149), .Y(n_516) );
AND2x2_ASAP7_75t_L g168 ( .A(n_11), .B(n_156), .Y(n_168) );
AND2x2_ASAP7_75t_L g177 ( .A(n_12), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g153 ( .A(n_13), .Y(n_153) );
AOI221x1_ASAP7_75t_L g469 ( .A1(n_14), .A2(n_25), .B1(n_131), .B2(n_140), .C(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_15), .B(n_147), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_16), .B(n_763), .C(n_765), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_17), .B(n_131), .Y(n_512) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_18), .A2(n_156), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_19), .B(n_151), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_147), .Y(n_523) );
AO21x1_ASAP7_75t_L g534 ( .A1(n_21), .A2(n_131), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_22), .B(n_131), .Y(n_211) );
INVx1_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
NOR2xp33_ASAP7_75t_SL g760 ( .A(n_23), .B(n_116), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_24), .A2(n_90), .B1(n_131), .B2(n_241), .Y(n_240) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_26), .B(n_147), .Y(n_479) );
NAND2x1_ASAP7_75t_L g505 ( .A(n_27), .B(n_149), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_28), .Y(n_452) );
OR2x2_ASAP7_75t_L g154 ( .A(n_29), .B(n_87), .Y(n_154) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_29), .A2(n_87), .B(n_153), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_30), .B(n_149), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_31), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_32), .B(n_147), .Y(n_515) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_33), .A2(n_178), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_34), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_35), .B(n_149), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_36), .A2(n_140), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_37), .B(n_147), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_38), .A2(n_140), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g137 ( .A(n_39), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g141 ( .A(n_39), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g249 ( .A(n_39), .Y(n_249) );
OR2x6_ASAP7_75t_L g113 ( .A(n_40), .B(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g765 ( .A(n_40), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_41), .B(n_131), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_42), .B(n_131), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_43), .B(n_147), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_44), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_45), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_46), .B(n_149), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_47), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_48), .A2(n_140), .B(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_49), .A2(n_140), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_50), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_51), .B(n_149), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_52), .B(n_131), .Y(n_183) );
INVx1_ASAP7_75t_L g134 ( .A(n_53), .Y(n_134) );
INVx1_ASAP7_75t_L g144 ( .A(n_53), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_54), .B(n_147), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_55), .A2(n_62), .B1(n_120), .B2(n_121), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_55), .Y(n_120) );
AND2x2_ASAP7_75t_L g202 ( .A(n_56), .B(n_151), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_57), .B(n_149), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_58), .B(n_147), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_59), .B(n_149), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_60), .A2(n_140), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_61), .B(n_131), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_62), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_63), .B(n_131), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_64), .A2(n_140), .B(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g217 ( .A(n_65), .B(n_152), .Y(n_217) );
AO21x1_ASAP7_75t_L g536 ( .A1(n_66), .A2(n_140), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_67), .B(n_131), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_68), .B(n_149), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_69), .B(n_131), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_70), .B(n_149), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_71), .A2(n_95), .B1(n_140), .B2(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_72), .B(n_147), .Y(n_214) );
AND2x2_ASAP7_75t_L g490 ( .A(n_73), .B(n_152), .Y(n_490) );
INVx1_ASAP7_75t_L g136 ( .A(n_74), .Y(n_136) );
INVx1_ASAP7_75t_L g142 ( .A(n_74), .Y(n_142) );
AND2x2_ASAP7_75t_L g508 ( .A(n_75), .B(n_178), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_76), .B(n_149), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_77), .A2(n_140), .B(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_78), .A2(n_140), .B(n_145), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_79), .A2(n_140), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g197 ( .A(n_80), .B(n_152), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_81), .B(n_151), .Y(n_238) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
AND2x2_ASAP7_75t_L g494 ( .A(n_83), .B(n_178), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_84), .B(n_131), .Y(n_525) );
AND2x2_ASAP7_75t_L g155 ( .A(n_85), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g535 ( .A(n_86), .B(n_188), .Y(n_535) );
AND2x2_ASAP7_75t_L g482 ( .A(n_88), .B(n_178), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_89), .B(n_149), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_91), .B(n_147), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_92), .B(n_149), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_93), .A2(n_140), .B(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_94), .A2(n_140), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_96), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_97), .B(n_147), .Y(n_499) );
BUFx2_ASAP7_75t_L g216 ( .A(n_98), .Y(n_216) );
BUFx2_ASAP7_75t_L g107 ( .A(n_99), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_100), .A2(n_140), .B(n_514), .Y(n_513) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_755), .B(n_766), .Y(n_101) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_453), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g754 ( .A(n_105), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_117), .B(n_451), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_109), .B(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x6_ASAP7_75t_SL g741 ( .A(n_111), .B(n_112), .Y(n_741) );
AND2x6_ASAP7_75t_SL g743 ( .A(n_111), .B(n_113), .Y(n_743) );
OR2x2_ASAP7_75t_L g752 ( .A(n_111), .B(n_113), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
NAND2x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_448), .Y(n_117) );
NAND2x1p5_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_119), .Y(n_450) );
INVx4_ASAP7_75t_L g449 ( .A(n_122), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_122), .A2(n_460), .B1(n_741), .B2(n_745), .Y(n_744) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_356), .Y(n_122) );
NOR3xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_279), .C(n_314), .Y(n_123) );
OAI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_179), .B(n_231), .C(n_269), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_158), .Y(n_126) );
AND2x2_ASAP7_75t_L g262 ( .A(n_127), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_127), .B(n_268), .Y(n_302) );
AND2x2_ASAP7_75t_L g327 ( .A(n_127), .B(n_282), .Y(n_327) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_L g234 ( .A(n_128), .Y(n_234) );
OR2x2_ASAP7_75t_L g265 ( .A(n_128), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_128), .B(n_169), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_128), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g308 ( .A(n_128), .B(n_309), .Y(n_308) );
NOR2x1_ASAP7_75t_L g319 ( .A(n_128), .B(n_311), .Y(n_319) );
AND2x4_ASAP7_75t_L g336 ( .A(n_128), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g374 ( .A(n_128), .Y(n_374) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_128), .B(n_159), .Y(n_379) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_155), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_139), .B(n_151), .Y(n_129) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
AND2x6_ASAP7_75t_L g149 ( .A(n_133), .B(n_142), .Y(n_149) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g147 ( .A(n_135), .B(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
AND2x2_ASAP7_75t_L g143 ( .A(n_138), .B(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_138), .Y(n_244) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx3_ASAP7_75t_L g245 ( .A(n_141), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_142), .Y(n_251) );
AND2x4_ASAP7_75t_L g247 ( .A(n_143), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g243 ( .A(n_144), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_150), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_149), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_150), .A2(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_150), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_150), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_150), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_150), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_150), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_150), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_150), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_150), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_150), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_150), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_150), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_150), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_150), .A2(n_538), .B(n_539), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_151), .Y(n_161) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_151), .A2(n_240), .B(n_246), .Y(n_239) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_151), .A2(n_469), .B(n_473), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_151), .A2(n_496), .B(n_497), .Y(n_495) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_151), .A2(n_469), .B(n_473), .Y(n_575) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x4_ASAP7_75t_L g188 ( .A(n_153), .B(n_154), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_156), .A2(n_211), .B(n_212), .Y(n_210) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g170 ( .A(n_157), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_158), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_158), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_169), .Y(n_158) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_159), .Y(n_274) );
INVx2_ASAP7_75t_L g310 ( .A(n_159), .Y(n_310) );
INVx1_ASAP7_75t_L g337 ( .A(n_159), .Y(n_337) );
AND2x2_ASAP7_75t_L g436 ( .A(n_159), .B(n_346), .Y(n_436) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_160), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_160), .B(n_169), .Y(n_282) );
AOI21x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_168), .Y(n_160) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_161), .A2(n_502), .B(n_508), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_167), .Y(n_162) );
INVx2_ASAP7_75t_L g311 ( .A(n_169), .Y(n_311) );
INVx2_ASAP7_75t_L g346 ( .A(n_169), .Y(n_346) );
OR2x2_ASAP7_75t_L g431 ( .A(n_169), .B(n_263), .Y(n_431) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_177), .Y(n_169) );
INVx4_ASAP7_75t_L g178 ( .A(n_170), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_176), .Y(n_171) );
INVx3_ASAP7_75t_L g190 ( .A(n_178), .Y(n_190) );
AOI211xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_198), .B(n_218), .C(n_225), .Y(n_179) );
INVx2_ASAP7_75t_SL g320 ( .A(n_180), .Y(n_320) );
AND2x2_ASAP7_75t_L g326 ( .A(n_180), .B(n_199), .Y(n_326) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_189), .Y(n_180) );
INVx1_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
INVx1_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
INVx2_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
AND2x2_ASAP7_75t_L g277 ( .A(n_181), .B(n_201), .Y(n_277) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_181), .Y(n_306) );
OR2x2_ASAP7_75t_L g386 ( .A(n_181), .B(n_209), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_188), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_188), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_188), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_SL g519 ( .A(n_188), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_188), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g252 ( .A(n_189), .B(n_253), .Y(n_252) );
NOR2x1_ASAP7_75t_SL g284 ( .A(n_189), .B(n_209), .Y(n_284) );
AO21x1_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_191), .B(n_197), .Y(n_189) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_190), .A2(n_191), .B(n_197), .Y(n_224) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_190), .A2(n_476), .B(n_482), .Y(n_475) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_190), .A2(n_484), .B(n_490), .Y(n_483) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_190), .A2(n_484), .B(n_490), .Y(n_542) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_190), .A2(n_476), .B(n_482), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_196), .Y(n_191) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_221), .Y(n_298) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
OR2x2_ASAP7_75t_L g230 ( .A(n_200), .B(n_209), .Y(n_230) );
BUFx2_ASAP7_75t_L g254 ( .A(n_200), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_200), .B(n_306), .Y(n_305) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
AND2x2_ASAP7_75t_L g283 ( .A(n_201), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g293 ( .A(n_201), .Y(n_293) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_201), .B(n_209), .Y(n_331) );
OR2x2_ASAP7_75t_L g406 ( .A(n_201), .B(n_223), .Y(n_406) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_SL g219 ( .A(n_209), .Y(n_219) );
AND2x2_ASAP7_75t_L g278 ( .A(n_209), .B(n_223), .Y(n_278) );
AND2x2_ASAP7_75t_L g349 ( .A(n_209), .B(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g370 ( .A(n_209), .Y(n_370) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_217), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g292 ( .A(n_221), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
BUFx2_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
AND2x2_ASAP7_75t_L g259 ( .A(n_223), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g350 ( .A(n_223), .Y(n_350) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
OR2x2_ASAP7_75t_L g296 ( .A(n_227), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_SL g338 ( .A(n_227), .B(n_339), .Y(n_338) );
AOI322xp5_ASAP7_75t_L g375 ( .A1(n_227), .A2(n_254), .A3(n_376), .B1(n_378), .B2(n_381), .C1(n_383), .C2(n_385), .Y(n_375) );
AND2x2_ASAP7_75t_L g440 ( .A(n_227), .B(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_228), .B(n_254), .Y(n_264) );
AOI322xp5_ASAP7_75t_L g315 ( .A1(n_229), .A2(n_316), .A3(n_320), .B1(n_321), .B2(n_324), .C1(n_326), .C2(n_327), .Y(n_315) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g367 ( .A(n_230), .B(n_320), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_230), .A2(n_427), .B1(n_429), .B2(n_432), .Y(n_426) );
OR2x2_ASAP7_75t_L g444 ( .A(n_230), .B(n_393), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_254), .B(n_255), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AOI221xp5_ASAP7_75t_SL g294 ( .A1(n_233), .A2(n_270), .B1(n_295), .B2(n_298), .C(n_299), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_233), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_234), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g363 ( .A(n_234), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g392 ( .A(n_235), .Y(n_392) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_252), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_236), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g334 ( .A(n_236), .Y(n_334) );
OR2x2_ASAP7_75t_L g341 ( .A(n_236), .B(n_342), .Y(n_341) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g384 ( .A(n_237), .B(n_346), .Y(n_384) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x4_ASAP7_75t_L g263 ( .A(n_238), .B(n_239), .Y(n_263) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NOR2x1p5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_252), .B(n_313), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_252), .B(n_293), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_252), .Y(n_393) );
INVx1_ASAP7_75t_L g260 ( .A(n_253), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_261), .B1(n_264), .B2(n_265), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_SL g371 ( .A(n_259), .Y(n_371) );
AND2x2_ASAP7_75t_L g428 ( .A(n_260), .B(n_284), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_262), .B(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g300 ( .A(n_262), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_262), .B(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
INVx2_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
AND2x2_ASAP7_75t_L g361 ( .A(n_263), .B(n_345), .Y(n_361) );
INVx1_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI21xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_275), .B(n_276), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g354 ( .A(n_273), .Y(n_354) );
INVx2_ASAP7_75t_L g342 ( .A(n_274), .Y(n_342) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g339 ( .A(n_278), .B(n_293), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g399 ( .A1(n_278), .A2(n_376), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_294), .Y(n_279) );
AOI32xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .A3(n_285), .B1(n_289), .B2(n_292), .Y(n_280) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_281), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_281), .A2(n_370), .B1(n_388), .B2(n_390), .C(n_396), .Y(n_387) );
AND2x2_ASAP7_75t_L g407 ( .A(n_281), .B(n_288), .Y(n_407) );
BUFx2_ASAP7_75t_L g291 ( .A(n_282), .Y(n_291) );
INVx1_ASAP7_75t_L g416 ( .A(n_282), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_282), .Y(n_421) );
INVx1_ASAP7_75t_SL g414 ( .A(n_283), .Y(n_414) );
INVx2_ASAP7_75t_L g297 ( .A(n_284), .Y(n_297) );
AND2x2_ASAP7_75t_L g409 ( .A(n_285), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g381 ( .A(n_287), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g353 ( .A(n_288), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_288), .B(n_379), .Y(n_401) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g303 ( .A(n_297), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_297), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g417 ( .A(n_298), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_307), .B2(n_312), .Y(n_299) );
INVx2_ASAP7_75t_SL g391 ( .A(n_301), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_301), .B(n_430), .Y(n_432) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_303), .A2(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g348 ( .A(n_305), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g376 ( .A(n_308), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
INVx1_ASAP7_75t_L g410 ( .A(n_312), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_328), .C(n_351), .Y(n_314) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx2_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_317), .B(n_336), .Y(n_395) );
OR2x2_ASAP7_75t_L g434 ( .A(n_317), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_318), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g330 ( .A(n_320), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g397 ( .A(n_323), .B(n_334), .Y(n_397) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_326), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g438 ( .A(n_326), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_336), .B2(n_338), .C(n_340), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_329), .A2(n_352), .B(n_355), .Y(n_351) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_331), .B(n_425), .Y(n_424) );
INVxp33_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g343 ( .A(n_339), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_344), .B2(n_347), .Y(n_340) );
INVx2_ASAP7_75t_L g446 ( .A(n_342), .Y(n_446) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g425 ( .A(n_350), .Y(n_425) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_402), .Y(n_356) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_375), .C(n_387), .D(n_399), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_366), .C(n_368), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_363), .A2(n_369), .B(n_372), .Y(n_368) );
INVx2_ASAP7_75t_L g447 ( .A(n_364), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_365), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OR2x2_ASAP7_75t_L g442 ( .A(n_370), .B(n_406), .Y(n_442) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_377), .Y(n_413) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_379), .B(n_384), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_379), .A2(n_409), .B(n_411), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_379), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g437 ( .A(n_379), .Y(n_437) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp33_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B1(n_393), .B2(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_408), .C(n_418), .D(n_439), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_415), .B2(n_417), .Y(n_411) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI211xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_422), .B(n_426), .C(n_433), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B(n_438), .Y(n_433) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_443), .B(n_445), .Y(n_439) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OAI22x1_ASAP7_75t_L g458 ( .A1(n_449), .A2(n_459), .B1(n_739), .B2(n_742), .Y(n_458) );
INVxp33_ASAP7_75t_L g753 ( .A(n_451), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_753), .B(n_754), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_744), .B2(n_747), .C(n_748), .Y(n_454) );
INVx1_ASAP7_75t_L g747 ( .A(n_455), .Y(n_747) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_651), .Y(n_460) );
AND4x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_563), .C(n_590), .D(n_625), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_491), .B1(n_528), .B2(n_543), .C(n_547), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_465), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g604 ( .A(n_466), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g659 ( .A(n_466), .B(n_614), .Y(n_659) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g562 ( .A(n_467), .B(n_483), .Y(n_562) );
AND2x4_ASAP7_75t_L g598 ( .A(n_467), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g612 ( .A(n_467), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_468), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_SL g556 ( .A1(n_474), .A2(n_529), .B(n_557), .C(n_561), .Y(n_556) );
AND2x2_ASAP7_75t_L g577 ( .A(n_474), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_474), .B(n_529), .Y(n_717) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .Y(n_474) );
INVx2_ASAP7_75t_L g597 ( .A(n_475), .Y(n_597) );
BUFx3_ASAP7_75t_L g613 ( .A(n_475), .Y(n_613) );
INVxp67_ASAP7_75t_L g617 ( .A(n_475), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g596 ( .A(n_483), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_483), .B(n_575), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_483), .B(n_597), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_485), .B(n_489), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_491), .A2(n_626), .B(n_629), .C(n_639), .Y(n_625) );
AND2x2_ASAP7_75t_SL g491 ( .A(n_492), .B(n_509), .Y(n_491) );
OAI321xp33_ASAP7_75t_L g600 ( .A1(n_492), .A2(n_548), .A3(n_601), .B1(n_603), .B2(n_604), .C(n_606), .Y(n_600) );
AND2x2_ASAP7_75t_L g721 ( .A(n_492), .B(n_696), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_492), .Y(n_724) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
INVx5_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_493), .B(n_560), .Y(n_559) );
NOR2x1_ASAP7_75t_SL g591 ( .A(n_493), .B(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g636 ( .A(n_493), .Y(n_636) );
AND2x2_ASAP7_75t_L g738 ( .A(n_493), .B(n_510), .Y(n_738) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x2_ASAP7_75t_L g545 ( .A(n_501), .B(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_501), .Y(n_555) );
INVx4_ASAP7_75t_L g560 ( .A(n_501), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .Y(n_502) );
INVx1_ASAP7_75t_L g603 ( .A(n_509), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_R g706 ( .A1(n_509), .A2(n_545), .B(n_577), .C(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g726 ( .A(n_509), .B(n_551), .Y(n_726) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .Y(n_509) );
INVx1_ASAP7_75t_L g544 ( .A(n_510), .Y(n_544) );
INVx2_ASAP7_75t_L g550 ( .A(n_510), .Y(n_550) );
OR2x2_ASAP7_75t_L g569 ( .A(n_510), .B(n_560), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_510), .B(n_592), .Y(n_638) );
BUFx3_ASAP7_75t_L g645 ( .A(n_510), .Y(n_645) );
INVx1_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_517), .Y(n_621) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
INVx1_ASAP7_75t_L g663 ( .A(n_518), .Y(n_663) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_526), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_519), .B(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g592 ( .A1(n_519), .A2(n_520), .B(n_526), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AND2x2_ASAP7_75t_L g564 ( .A(n_528), .B(n_565), .Y(n_564) );
OAI31xp33_ASAP7_75t_L g715 ( .A1(n_528), .A2(n_716), .A3(n_718), .B(n_721), .Y(n_715) );
INVx1_ASAP7_75t_SL g733 ( .A(n_528), .Y(n_733) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AOI21xp33_ASAP7_75t_L g547 ( .A1(n_529), .A2(n_548), .B(n_556), .Y(n_547) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_529), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g656 ( .A(n_529), .Y(n_656) );
INVx2_ASAP7_75t_L g605 ( .A(n_530), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_530), .B(n_588), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_530), .B(n_587), .Y(n_697) );
NOR2xp33_ASAP7_75t_SL g705 ( .A(n_530), .B(n_656), .Y(n_705) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_531), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g585 ( .A(n_531), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g614 ( .A(n_531), .B(n_596), .Y(n_614) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g599 ( .A(n_533), .Y(n_599) );
OAI21x1_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_536), .B(n_540), .Y(n_533) );
INVx1_ASAP7_75t_L g541 ( .A(n_535), .Y(n_541) );
INVx2_ASAP7_75t_L g586 ( .A(n_542), .Y(n_586) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_542), .Y(n_646) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
AND2x2_ASAP7_75t_L g661 ( .A(n_544), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g572 ( .A(n_545), .B(n_566), .Y(n_572) );
INVx2_ASAP7_75t_SL g620 ( .A(n_545), .Y(n_620) );
INVx4_ASAP7_75t_L g551 ( .A(n_546), .Y(n_551) );
AND2x2_ASAP7_75t_L g649 ( .A(n_546), .B(n_592), .Y(n_649) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_546), .B(n_662), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_546), .B(n_560), .Y(n_684) );
INVx1_ASAP7_75t_L g690 ( .A(n_548), .Y(n_690) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g609 ( .A(n_549), .Y(n_609) );
OR2x2_ASAP7_75t_L g622 ( .A(n_549), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OR2x2_ASAP7_75t_L g674 ( .A(n_550), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g704 ( .A(n_550), .B(n_592), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_551), .B(n_554), .Y(n_580) );
AND2x2_ASAP7_75t_L g672 ( .A(n_551), .B(n_662), .Y(n_672) );
AND2x4_ASAP7_75t_L g734 ( .A(n_551), .B(n_613), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx2_ASAP7_75t_L g558 ( .A(n_553), .Y(n_558) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp67_ASAP7_75t_SL g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI322xp33_ASAP7_75t_SL g570 ( .A1(n_558), .A2(n_571), .A3(n_573), .B1(n_576), .B2(n_579), .C1(n_581), .C2(n_583), .Y(n_570) );
INVx1_ASAP7_75t_L g728 ( .A(n_558), .Y(n_728) );
OR2x2_ASAP7_75t_L g581 ( .A(n_559), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g607 ( .A(n_560), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_560), .B(n_608), .Y(n_623) );
INVx2_ASAP7_75t_L g650 ( .A(n_560), .Y(n_650) );
AND2x4_ASAP7_75t_L g662 ( .A(n_560), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_562), .B(n_578), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_568), .B(n_570), .Y(n_563) );
AND2x2_ASAP7_75t_L g631 ( .A(n_565), .B(n_598), .Y(n_631) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_566), .B(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g589 ( .A(n_567), .Y(n_589) );
AND2x4_ASAP7_75t_SL g671 ( .A(n_567), .B(n_586), .Y(n_671) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g579 ( .A(n_569), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_572), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g707 ( .A(n_574), .B(n_671), .Y(n_707) );
NOR4xp25_ASAP7_75t_L g711 ( .A(n_574), .B(n_588), .C(n_628), .D(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g588 ( .A(n_575), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g624 ( .A(n_575), .B(n_599), .Y(n_624) );
AND2x4_ASAP7_75t_L g688 ( .A(n_575), .B(n_599), .Y(n_688) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_578), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
OR2x2_ASAP7_75t_L g677 ( .A(n_585), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g731 ( .A(n_585), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_586), .B(n_598), .Y(n_632) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AOI211xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_593), .B(n_600), .C(n_615), .Y(n_590) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_596), .B(n_599), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_597), .B(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g679 ( .A(n_597), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_598), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g694 ( .A(n_598), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_610), .Y(n_606) );
AND2x4_ASAP7_75t_L g643 ( .A(n_607), .B(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g737 ( .A(n_607), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_SL g641 ( .A(n_613), .Y(n_641) );
AND2x2_ASAP7_75t_L g700 ( .A(n_614), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g714 ( .A(n_614), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_618), .B(n_622), .C(n_624), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_616), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g692 ( .A(n_617), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g713 ( .A(n_617), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
OR2x2_ASAP7_75t_L g702 ( .A(n_620), .B(n_644), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_623), .A2(n_630), .B1(n_632), .B2(n_633), .Y(n_629) );
INVx1_ASAP7_75t_SL g720 ( .A(n_624), .Y(n_720) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_635), .B(n_644), .Y(n_686) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_638), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_646), .B2(n_647), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI21xp5_ASAP7_75t_SL g653 ( .A1(n_644), .A2(n_654), .B(n_657), .Y(n_653) );
AND2x2_ASAP7_75t_L g682 ( .A(n_644), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND3x2_ASAP7_75t_L g648 ( .A(n_645), .B(n_649), .C(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g710 ( .A(n_645), .B(n_667), .Y(n_710) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g695 ( .A(n_650), .B(n_696), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_652), .B(n_708), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_668), .C(n_689), .D(n_706), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_664), .B2(n_666), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_660), .A2(n_674), .B1(n_694), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g675 ( .A(n_662), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_664), .A2(n_687), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_673), .B2(n_676), .C(n_680), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_683), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_683), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_692), .B(n_694), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g723 ( .A1(n_704), .A2(n_724), .B(n_725), .C(n_727), .Y(n_723) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_715), .C(n_722), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_729), .B1(n_732), .B2(n_734), .C(n_735), .Y(n_722) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
CKINVDCx11_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g746 ( .A(n_742), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
CKINVDCx6p67_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_SL g769 ( .A(n_758), .Y(n_769) );
OR2x2_ASAP7_75t_SL g758 ( .A(n_759), .B(n_761), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
BUFx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
endmodule