module fake_jpeg_7731_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_40),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_25),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_56),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_43),
.B(n_25),
.C(n_31),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_57),
.B(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_18),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_23),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_27),
.B1(n_19),
.B2(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_78),
.B1(n_95),
.B2(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_83),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_34),
.B(n_35),
.C(n_30),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_79),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_17),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_101),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_R g121 ( 
.A(n_99),
.B(n_35),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_79),
.B(n_17),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_12),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_14),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_96),
.B1(n_112),
.B2(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_58),
.B1(n_46),
.B2(n_51),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_72),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_62),
.C(n_64),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_34),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_122),
.Y(n_140)
);

OAI22x1_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_97),
.B1(n_110),
.B2(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_128),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_81),
.B(n_73),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_77),
.B1(n_93),
.B2(n_92),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_92),
.B1(n_84),
.B2(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_94),
.B1(n_84),
.B2(n_23),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_143),
.B(n_150),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_144),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_102),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_108),
.B1(n_109),
.B2(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_153),
.B1(n_105),
.B2(n_124),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_105),
.B(n_98),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_101),
.C(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_132),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_151),
.C(n_143),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_125),
.B1(n_137),
.B2(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_162),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_13),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_14),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_138),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_170),
.C(n_176),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_164),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_179),
.C(n_183),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_161),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_160),
.B1(n_145),
.B2(n_158),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_182),
.B1(n_175),
.B2(n_139),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_155),
.B1(n_145),
.B2(n_147),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_155),
.B1(n_177),
.B2(n_147),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_179),
.C(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_174),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_0),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_151),
.B1(n_149),
.B2(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_186),
.A2(n_173),
.B(n_139),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_0),
.B(n_1),
.Y(n_196)
);

AOI21x1_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_7),
.B(n_3),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_194),
.A2(n_188),
.B1(n_185),
.B2(n_8),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_197),
.B(n_193),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_2),
.B(n_3),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.Y(n_201)
);


endmodule