module real_jpeg_9896_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_178;
wire n_67;
wire n_79;
wire n_76;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_62),
.B1(n_68),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_1),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_129),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_129),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_129),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_69),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_69),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_62),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_71),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_57),
.B1(n_62),
.B2(n_68),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_52),
.B(n_64),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_12),
.A2(n_62),
.B1(n_68),
.B2(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_12),
.B(n_156),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_12),
.A2(n_38),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_12),
.B(n_38),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_209),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_51),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_51),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_13),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_15),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_17),
.A2(n_62),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_17),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_17),
.A2(n_51),
.B1(n_52),
.B2(n_89),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_89),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_17),
.A2(n_38),
.B1(n_39),
.B2(n_89),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_21),
.B(n_93),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_79),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_23),
.B1(n_73),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_59),
.C(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_25),
.B(n_36),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_26),
.A2(n_33),
.B1(n_82),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_26),
.A2(n_33),
.B1(n_192),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_26),
.A2(n_33),
.B1(n_194),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_26),
.A2(n_33),
.B1(n_225),
.B2(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_27),
.A2(n_28),
.B1(n_137),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_27),
.A2(n_28),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_29),
.B(n_44),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_29),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_30),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_33),
.B(n_133),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_50),
.B2(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_38),
.B(n_55),
.Y(n_237)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_39),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_41),
.A2(n_43),
.B1(n_77),
.B2(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_41),
.A2(n_43),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_41),
.A2(n_43),
.B1(n_200),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_41),
.A2(n_43),
.B1(n_223),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_41),
.A2(n_43),
.B1(n_159),
.B2(n_230),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_43),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_43),
.B(n_133),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_54),
.B1(n_58),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_49),
.A2(n_54),
.B1(n_92),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_49),
.A2(n_54),
.B1(n_124),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_49),
.A2(n_54),
.B1(n_152),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_49),
.A2(n_54),
.B1(n_178),
.B2(n_232),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_66)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_54),
.B(n_133),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_66),
.B1(n_70),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_61),
.A2(n_66),
.B1(n_88),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_62),
.A2(n_63),
.B(n_133),
.C(n_134),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_73),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_75),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.C(n_90),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_81),
.B(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_110),
.B2(n_111),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_101),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_105),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_141),
.B(n_264),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_138),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_116),
.B(n_138),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_120),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_119),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_121),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_125),
.C(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_183),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_165),
.B(n_182),
.Y(n_143)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_144),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_162),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_162),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_157),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_151),
.B1(n_157),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_166),
.B(n_168),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_172),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_177),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_180),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_181),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_262),
.C(n_263),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_256),
.B(n_261),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_242),
.B(n_255),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_227),
.B(n_241),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_217),
.B(n_226),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_206),
.B(n_216),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_195),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_205),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_205),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_201),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_228),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.CI(n_224),
.CON(n_220),
.SN(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.CI(n_234),
.CON(n_228),
.SN(n_228)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_243),
.B(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_252),
.C(n_253),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_251),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);


endmodule