module fake_jpeg_7715_n_49 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_49);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_27),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_28),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_8),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.C(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_12),
.C(n_13),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_14),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_15),
.B(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_31),
.Y(n_45)
);

XNOR2x1_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.C(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_43),
.C(n_44),
.Y(n_49)
);


endmodule