module real_jpeg_2911_n_16 (n_5, n_4, n_8, n_0, n_12, n_408, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_407, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_408;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_407;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_0),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_0),
.B(n_97),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_99),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_0),
.B(n_62),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_0),
.B(n_54),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_0),
.B(n_29),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_0),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_26),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_4),
.B(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_4),
.B(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_4),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_54),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_29),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_4),
.B(n_23),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_4),
.B(n_26),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_6),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_6),
.B(n_97),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_6),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_6),
.B(n_34),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_9),
.B(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_9),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_23),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_9),
.B(n_26),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_9),
.B(n_34),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_34),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_13),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_13),
.B(n_97),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_62),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_13),
.B(n_54),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_13),
.B(n_29),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_14),
.B(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_14),
.B(n_54),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_29),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_23),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_29),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_15),
.B(n_99),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_15),
.B(n_54),
.Y(n_268)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_57),
.B(n_83),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_57),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_25),
.C(n_28),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_21),
.A2(n_22),
.B1(n_28),
.B2(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_21),
.A2(n_22),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_22),
.B(n_285),
.C(n_286),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_23),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_25),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_25),
.A2(n_49),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_25),
.B(n_268),
.C(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_28),
.A2(n_48),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_28),
.A2(n_48),
.B1(n_248),
.B2(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_28),
.B(n_170),
.C(n_249),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_29),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_53),
.C(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_31),
.A2(n_40),
.B1(n_61),
.B2(n_185),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_32),
.B(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_32),
.B(n_130),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_33),
.B(n_104),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_33),
.B(n_134),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_33),
.B(n_156),
.Y(n_331)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_38),
.A2(n_39),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_38),
.B(n_314),
.C(n_316),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_38),
.A2(n_39),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_38),
.B(n_354),
.C(n_357),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.C(n_52),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_45),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.C(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_53),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_53),
.B(n_227),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_53),
.A2(n_76),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_56),
.A2(n_77),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_78),
.C(n_79),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_58),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_68),
.C(n_73),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_59),
.B(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_64),
.C(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_61),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_61),
.B(n_182),
.C(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_61),
.A2(n_185),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_61),
.B(n_167),
.C(n_339),
.Y(n_382)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_65),
.B(n_137),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_66),
.B(n_134),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_68),
.B(n_73),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.C(n_72),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_389),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_69),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_70),
.A2(n_71),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_71),
.B(n_122),
.C(n_190),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_72),
.B(n_388),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_77),
.B(n_167),
.C(n_323),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_78),
.B(n_79),
.Y(n_403)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_401),
.B(n_405),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_374),
.A3(n_392),
.B1(n_399),
.B2(n_400),
.C(n_407),
.Y(n_85)
);

AOI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_304),
.A3(n_363),
.B1(n_368),
.B2(n_373),
.C(n_408),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_240),
.C(n_300),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_206),
.B(n_239),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_174),
.B(n_205),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_149),
.B(n_173),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_126),
.B(n_148),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_106),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_93),
.B(n_106),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.C(n_105),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_95),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_96),
.B(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_137),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_116),
.C(n_120),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_112),
.C(n_113),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_121),
.A2(n_122),
.B1(n_190),
.B2(n_192),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_121),
.A2(n_122),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_123),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_122),
.B(n_234),
.C(n_331),
.Y(n_354)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_139),
.B(n_147),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_132),
.B(n_138),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_184),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_163),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_162),
.C(n_163),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_159),
.C(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_172),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_166),
.C(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_167),
.A2(n_171),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_167),
.A2(n_171),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_169),
.A2(n_170),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_176),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_194),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_195),
.C(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_186),
.B2(n_187),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_188),
.C(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_184),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_204),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_224),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_222),
.B2(n_223),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_211),
.B(n_223),
.C(n_224),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_220),
.C(n_221),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_255),
.C(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_234),
.A2(n_235),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g369 ( 
.A1(n_241),
.A2(n_370),
.B(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_273),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_242),
.B(n_273),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_259),
.C(n_260),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_246),
.C(n_253),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_257),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_260),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_272),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_265),
.C(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_268),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_268),
.A2(n_269),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_299),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_288),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_275),
.B(n_288),
.C(n_299),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_280),
.C(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_284),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_297),
.C(n_298),
.Y(n_311)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_302),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_333),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_305),
.B(n_333),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_317),
.C(n_332),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_317),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_311),
.C(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_326),
.C(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_348),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_348),
.C(n_362),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_342),
.C(n_343),
.Y(n_390)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_346),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_359),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_352),
.C(n_353),
.Y(n_391)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_351),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_360),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_364),
.A2(n_369),
.B(n_372),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_365),
.B(n_366),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_375),
.B(n_376),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_393),
.Y(n_400)
);

FAx1_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_384),
.CI(n_391),
.CON(n_376),
.SN(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_382),
.C(n_383),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_387),
.C(n_390),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_396),
.C(n_398),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_404),
.Y(n_405)
);


endmodule