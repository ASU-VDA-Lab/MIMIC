module fake_jpeg_3729_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_60),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_59),
.B1(n_23),
.B2(n_17),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_30),
.B1(n_28),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_50),
.B1(n_14),
.B2(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_30),
.B1(n_28),
.B2(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_27),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_35),
.B1(n_42),
.B2(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_71),
.B1(n_79),
.B2(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_72),
.Y(n_97)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_74),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_35),
.B1(n_26),
.B2(n_14),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_29),
.B1(n_16),
.B2(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_44),
.B(n_47),
.C(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_42),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_72),
.C(n_64),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_97),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_68),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_54),
.C(n_66),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_102),
.B1(n_74),
.B2(n_51),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_54),
.B1(n_33),
.B2(n_34),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_54),
.B(n_76),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_118),
.B(n_95),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_91),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_54),
.B(n_70),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_109),
.B(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_69),
.B1(n_63),
.B2(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_112),
.B1(n_40),
.B2(n_39),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_40),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_69),
.B1(n_40),
.B2(n_51),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_87),
.B1(n_98),
.B2(n_96),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_82),
.B(n_101),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_34),
.B(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_124),
.C(n_125),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_110),
.B(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_128),
.B(n_116),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_117),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_88),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_102),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_112),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_93),
.CI(n_82),
.CON(n_127),
.SN(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_118),
.B1(n_108),
.B2(n_114),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_142),
.B1(n_127),
.B2(n_131),
.Y(n_143)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_103),
.B(n_107),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_129),
.C(n_130),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_108),
.B(n_109),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_136),
.B(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_140),
.C(n_123),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_125),
.C(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.C(n_151),
.Y(n_153)
);

AOI21x1_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_116),
.B(n_22),
.Y(n_146)
);

XOR2x1_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_22),
.C(n_21),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_134),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_1),
.C(n_4),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_140),
.C(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_147),
.C(n_148),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_136),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_136),
.B1(n_5),
.B2(n_7),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_151),
.C(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_150),
.C(n_144),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_152),
.B(n_154),
.C(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_163),
.B(n_10),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_11),
.B(n_72),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_11),
.Y(n_167)
);


endmodule