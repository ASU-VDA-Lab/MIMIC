module fake_jpeg_18293_n_299 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_265;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_13),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_21),
.B1(n_30),
.B2(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_62),
.B(n_64),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_65),
.B(n_70),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_27),
.B1(n_34),
.B2(n_42),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_33),
.B(n_15),
.C(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_76),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_80),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_36),
.B1(n_23),
.B2(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_72)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_40),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_75),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_83),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_41),
.B1(n_38),
.B2(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_44),
.C(n_40),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_28),
.C(n_29),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_19),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_67),
.B(n_88),
.Y(n_111)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_30),
.B1(n_21),
.B2(n_14),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_93),
.B1(n_28),
.B2(n_20),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_17),
.B(n_19),
.C(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_19),
.B1(n_43),
.B2(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_19),
.B1(n_17),
.B2(n_26),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_29),
.B1(n_26),
.B2(n_2),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_28),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_29),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_11),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_20),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_65),
.B1(n_74),
.B2(n_100),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_64),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_120),
.B1(n_126),
.B2(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_68),
.A2(n_29),
.B1(n_26),
.B2(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_133),
.B1(n_127),
.B2(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_73),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_150),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_152),
.B1(n_154),
.B2(n_118),
.Y(n_169)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_148),
.Y(n_179)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_153),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_75),
.B1(n_93),
.B2(n_94),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_109),
.A2(n_80),
.B1(n_97),
.B2(n_96),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_81),
.B1(n_89),
.B2(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_134),
.B1(n_117),
.B2(n_119),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_106),
.B(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_97),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_12),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_12),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_110),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_167),
.A2(n_185),
.B(n_187),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_180),
.B1(n_142),
.B2(n_84),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_136),
.Y(n_216)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_109),
.B1(n_115),
.B2(n_107),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_110),
.B1(n_134),
.B2(n_117),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_144),
.B1(n_155),
.B2(n_148),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_194),
.B1(n_138),
.B2(n_139),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_137),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_108),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_133),
.B(n_135),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_140),
.B(n_84),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_125),
.B1(n_129),
.B2(n_135),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_200),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_143),
.B(n_165),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_175),
.B(n_192),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_147),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_172),
.B1(n_183),
.B2(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_206),
.B1(n_215),
.B2(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_138),
.C(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_191),
.C(n_179),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_156),
.B1(n_151),
.B2(n_129),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_132),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_142),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_140),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_225),
.B1(n_228),
.B2(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_227),
.C(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_176),
.C(n_193),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_176),
.B(n_181),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_202),
.B1(n_206),
.B2(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_170),
.C(n_146),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_238),
.C(n_107),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_172),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_209),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_170),
.C(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_208),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_248),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_217),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_212),
.C(n_196),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_254),
.C(n_256),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_201),
.B1(n_214),
.B2(n_205),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_190),
.B1(n_235),
.B2(n_237),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_211),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_205),
.C(n_204),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_204),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_256),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_225),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_195),
.C(n_177),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_235),
.B(n_232),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_264),
.B(n_229),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_267),
.C(n_254),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_259),
.B1(n_263),
.B2(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_252),
.C(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_123),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_242),
.C(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_273),
.C(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_266),
.B1(n_269),
.B2(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_237),
.C(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_229),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_121),
.C(n_123),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_250),
.B1(n_105),
.B2(n_78),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_61),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_282),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_78),
.B1(n_105),
.B2(n_166),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_166),
.B1(n_101),
.B2(n_79),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_285),
.A3(n_276),
.B1(n_270),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_289),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_290),
.B(n_283),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_282),
.B(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_292),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.C(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_283),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_4),
.Y(n_299)
);


endmodule