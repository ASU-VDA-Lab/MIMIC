module fake_jpeg_23441_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_1),
.B(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_57),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_26),
.B1(n_25),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_25),
.B1(n_33),
.B2(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_26),
.B1(n_36),
.B2(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_26),
.B1(n_36),
.B2(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_37),
.B1(n_22),
.B2(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_29),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_27),
.B1(n_37),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_79),
.B1(n_84),
.B2(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_1),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_28),
.B1(n_24),
.B2(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_28),
.B1(n_32),
.B2(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_31),
.B1(n_32),
.B2(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_34),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_85),
.B1(n_40),
.B2(n_39),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_20),
.B1(n_31),
.B2(n_2),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_0),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_20),
.B(n_40),
.C(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_108),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_116),
.B1(n_100),
.B2(n_109),
.Y(n_154)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_102),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_71),
.B1(n_96),
.B2(n_98),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_111),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_80),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_114),
.Y(n_153)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_89),
.B1(n_67),
.B2(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_50),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_1),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_54),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_65),
.C(n_64),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_145),
.Y(n_167)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_89),
.B1(n_69),
.B2(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_149),
.B1(n_90),
.B2(n_108),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_140),
.B1(n_143),
.B2(n_154),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_55),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_71),
.B1(n_61),
.B2(n_63),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_87),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_71),
.B1(n_61),
.B2(n_63),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_74),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_97),
.A2(n_64),
.B1(n_72),
.B2(n_78),
.Y(n_149)
);

FAx1_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_43),
.CI(n_57),
.CON(n_150),
.SN(n_150)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_125),
.B(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_159),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_168),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_106),
.B(n_112),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_166),
.B(n_174),
.Y(n_200)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_95),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_106),
.B(n_122),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_10),
.B(n_12),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_95),
.B(n_122),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_123),
.B1(n_114),
.B2(n_124),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_178),
.B1(n_183),
.B2(n_130),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_73),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_182),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_107),
.B1(n_43),
.B2(n_8),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_6),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_186),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_188),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_126),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_6),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_7),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_9),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_139),
.C(n_136),
.Y(n_207)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_197),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_219),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_149),
.B1(n_150),
.B2(n_129),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_206),
.B1(n_214),
.B2(n_181),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_150),
.B(n_141),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_203),
.B(n_213),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_126),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_216),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_152),
.B1(n_136),
.B2(n_139),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_217),
.B(n_221),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_144),
.B1(n_11),
.B2(n_12),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_191),
.B1(n_171),
.B2(n_188),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_138),
.B(n_11),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_138),
.B1(n_11),
.B2(n_12),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_162),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_13),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_13),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_164),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_160),
.A2(n_13),
.B(n_14),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_224),
.Y(n_246)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_240),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_167),
.C(n_192),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_189),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_211),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_186),
.B1(n_182),
.B2(n_163),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_242),
.A2(n_197),
.B1(n_214),
.B2(n_213),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_163),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_199),
.C(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_253),
.C(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_207),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_198),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_263),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_194),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_251),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_234),
.B(n_226),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_249),
.C(n_230),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_276),
.C(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_261),
.B(n_236),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_234),
.B(n_228),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_274),
.B(n_277),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_233),
.B(n_241),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_231),
.C(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_204),
.B1(n_228),
.B2(n_210),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_217),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_287),
.C(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_265),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_288),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_247),
.C(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_159),
.C(n_212),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_252),
.C(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_271),
.C(n_227),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_14),
.Y(n_300)
);

XOR2x1_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_203),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_278),
.B1(n_271),
.B2(n_203),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_201),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_273),
.C(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_301),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_299),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_304),
.B(n_307),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_299),
.B(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

NAND2x1_ASAP7_75t_SL g306 ( 
.A(n_293),
.B(n_288),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_180),
.B(n_272),
.C(n_268),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_293),
.B(n_284),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_14),
.B(n_15),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_268),
.B(n_181),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_306),
.A3(n_303),
.B1(n_190),
.B2(n_188),
.C1(n_168),
.C2(n_17),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_15),
.B(n_313),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_309),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);


endmodule