module fake_netlist_6_845_n_1987 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1987);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1987;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_131),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_181),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_55),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_30),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_6),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_77),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_62),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_115),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_112),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_73),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_45),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_25),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_143),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_24),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_6),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_26),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_85),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_142),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_153),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_50),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_88),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_75),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_59),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_37),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_8),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_114),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_7),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_151),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_193),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_122),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_61),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_171),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_10),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_71),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_61),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_124),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_59),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_10),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_21),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_33),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_191),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_116),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_195),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_74),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_48),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_107),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_161),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_12),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_97),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_23),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_28),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_54),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_26),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_128),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_120),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_132),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_113),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_74),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_175),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_135),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_4),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_23),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_130),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_103),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_1),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_0),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_72),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_178),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_71),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_69),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_98),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_46),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_118),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_64),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_152),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_48),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_57),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_93),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_5),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_32),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_187),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_127),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_83),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_34),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_109),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_19),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_121),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_65),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_11),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_82),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_43),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_89),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_55),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_99),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_19),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_70),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_31),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_63),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_119),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_17),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_100),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_104),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_165),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_52),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_162),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_15),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_167),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_186),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_149),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_42),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_67),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_28),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_54),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_192),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_108),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_53),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_73),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_31),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_170),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_41),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_173),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_43),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_35),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_36),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_92),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_13),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_17),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_179),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_69),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_58),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_156),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_21),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_169),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_155),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_29),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_84),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_14),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_51),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_47),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_57),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_3),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_94),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_154),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_200),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_230),
.B(n_0),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_272),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_198),
.B(n_2),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_212),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_198),
.B(n_2),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_243),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_323),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_254),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_276),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_259),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_234),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_298),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_303),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_252),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_262),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_261),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_270),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_274),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_275),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_276),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_282),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_299),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_301),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_199),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_304),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_306),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_276),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_310),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_206),
.B(n_3),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_311),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_315),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_276),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_309),
.B(n_7),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_320),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_325),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_328),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_329),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_276),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_289),
.B(n_9),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_224),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_309),
.B(n_9),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_330),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_246),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_294),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_251),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_334),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_246),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_238),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_196),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_339),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_342),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_221),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_342),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_238),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_348),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_296),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_229),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_289),
.B(n_11),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_207),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_235),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_350),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_207),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_354),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_242),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_355),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_391),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_201),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_199),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_201),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_202),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_247),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_332),
.B(n_14),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_203),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_244),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_203),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_202),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_264),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_248),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_205),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_249),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_204),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_429),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_442),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_205),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_459),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_425),
.B(n_332),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_459),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_208),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_448),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_211),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_459),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_465),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_208),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_462),
.B(n_213),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_396),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_460),
.B(n_396),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_478),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_398),
.B(n_210),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_460),
.B(n_218),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_467),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_407),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_408),
.B(n_210),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_408),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_449),
.B(n_241),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_412),
.B(n_214),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_245),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_413),
.B(n_238),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_479),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_413),
.B(n_214),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_416),
.B(n_250),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_255),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_393),
.B(n_256),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_421),
.B(n_215),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_424),
.B(n_257),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_424),
.B(n_427),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_437),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_468),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_265),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_468),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_450),
.B(n_215),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_483),
.B(n_238),
.Y(n_560)
);

CKINVDCx8_ASAP7_75t_R g561 ( 
.A(n_455),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_471),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_475),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_480),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_482),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_544),
.A2(n_392),
.B1(n_428),
.B2(n_420),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_496),
.B(n_455),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_527),
.B(n_397),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_557),
.B(n_544),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_531),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_557),
.B(n_470),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_531),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_517),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_557),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_557),
.B(n_473),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_SL g584 ( 
.A1(n_507),
.A2(n_452),
.B(n_443),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_559),
.B(n_439),
.C(n_402),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_557),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_556),
.A2(n_557),
.B1(n_560),
.B2(n_508),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_513),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_557),
.B(n_473),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_526),
.B(n_400),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_514),
.B(n_405),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_526),
.B(n_417),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_531),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_549),
.B(n_443),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_515),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_493),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_515),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_559),
.A2(n_399),
.B1(n_347),
.B2(n_233),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_561),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_493),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_493),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_556),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_526),
.B(n_422),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_431),
.B1(n_456),
.B2(n_394),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_507),
.B(n_423),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_560),
.B(n_238),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_561),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_514),
.B(n_426),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_509),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_509),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_531),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_509),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_509),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_451),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_561),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_522),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_522),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_518),
.B(n_430),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_518),
.B(n_433),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_510),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_563),
.B(n_441),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_520),
.B(n_447),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_516),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_549),
.B(n_452),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_563),
.B(n_453),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_523),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_538),
.A2(n_438),
.B1(n_440),
.B2(n_435),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_520),
.B(n_457),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_525),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_549),
.B(n_463),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_516),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_496),
.B(n_492),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_556),
.B(n_263),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_R g651 ( 
.A(n_568),
.B(n_432),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_508),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_514),
.B(n_476),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_532),
.B(n_536),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_532),
.B(n_454),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_519),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_519),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_538),
.A2(n_456),
.B1(n_431),
.B2(n_267),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_528),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_548),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_551),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_503),
.B(n_263),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_501),
.B(n_477),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_535),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_517),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_454),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_536),
.B(n_458),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_508),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_510),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_528),
.Y(n_671)
);

AO22x2_ASAP7_75t_L g672 ( 
.A1(n_569),
.A2(n_364),
.B1(n_314),
.B2(n_292),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_568),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_530),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_548),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_498),
.B(n_529),
.Y(n_676)
);

INVxp33_ASAP7_75t_SL g677 ( 
.A(n_524),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_498),
.B(n_362),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_551),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_541),
.B(n_263),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_535),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_501),
.B(n_484),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_444),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_530),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_560),
.A2(n_324),
.B1(n_345),
.B2(n_335),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_529),
.B(n_445),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_549),
.B(n_463),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_524),
.B(n_458),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_533),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_541),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_533),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_498),
.B(n_271),
.Y(n_693)
);

AO21x2_ASAP7_75t_L g694 ( 
.A1(n_534),
.A2(n_288),
.B(n_283),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_534),
.B(n_446),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_540),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_539),
.B(n_464),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_549),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_539),
.B(n_461),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

NOR2x1p5_ASAP7_75t_L g702 ( 
.A(n_527),
.B(n_204),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_546),
.B(n_466),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_552),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_551),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_527),
.B(n_464),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_552),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_503),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_503),
.B(n_279),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_553),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_540),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_541),
.B(n_263),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_537),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_541),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_553),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_499),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_503),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_503),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_498),
.B(n_291),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_682),
.B(n_472),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_661),
.B(n_543),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_719),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_691),
.Y(n_725)
);

AND2x4_ASAP7_75t_SL g726 ( 
.A(n_626),
.B(n_406),
.Y(n_726)
);

INVx8_ASAP7_75t_L g727 ( 
.A(n_643),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_588),
.A2(n_474),
.B1(n_418),
.B2(n_415),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_587),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_587),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_691),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_675),
.B(n_543),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_576),
.B(n_543),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_543),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_652),
.B(n_481),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_589),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_603),
.B(n_613),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_652),
.B(n_487),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_598),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_598),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_600),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_600),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_607),
.B(n_611),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_669),
.A2(n_490),
.B1(n_411),
.B2(n_410),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_703),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_632),
.B(n_543),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_703),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_664),
.B(n_547),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_639),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_716),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_669),
.A2(n_547),
.B1(n_521),
.B2(n_560),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_582),
.B(n_547),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_716),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_710),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_710),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_720),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_642),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_628),
.B(n_547),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_628),
.B(n_547),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_582),
.B(n_560),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_689),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_647),
.B(n_521),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_718),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_578),
.A2(n_521),
.B1(n_560),
.B2(n_222),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_586),
.B(n_560),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_666),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_647),
.B(n_521),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_574),
.B(n_697),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_630),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_628),
.B(n_499),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_586),
.B(n_560),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_708),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_676),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_574),
.B(n_521),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_642),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_583),
.B(n_216),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_720),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_644),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_666),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_590),
.B(n_216),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_697),
.B(n_219),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_718),
.B(n_499),
.Y(n_782)
);

NAND2x1p5_ASAP7_75t_L g783 ( 
.A(n_698),
.B(n_499),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_718),
.Y(n_784)
);

AND2x2_ASAP7_75t_SL g785 ( 
.A(n_612),
.B(n_263),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_671),
.B(n_560),
.Y(n_787)
);

BUFx5_ASAP7_75t_L g788 ( 
.A(n_720),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_671),
.B(n_560),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_584),
.B(n_219),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_585),
.B(n_222),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_663),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_223),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_630),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_573),
.B(n_223),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_674),
.Y(n_796)
);

INVx8_ASAP7_75t_L g797 ( 
.A(n_643),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_596),
.A2(n_300),
.B1(n_305),
.B2(n_318),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_663),
.B(n_499),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_715),
.B(n_356),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_689),
.B(n_558),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_555),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_690),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_692),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_670),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_555),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_700),
.B(n_701),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_700),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_640),
.B(n_558),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_715),
.B(n_356),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_686),
.B(n_225),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_701),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_708),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_683),
.B(n_373),
.C(n_562),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_225),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_711),
.B(n_562),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_699),
.B(n_566),
.C(n_565),
.Y(n_818)
);

AND2x6_ASAP7_75t_SL g819 ( 
.A(n_643),
.B(n_280),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_670),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_705),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_616),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_694),
.A2(n_554),
.B1(n_550),
.B2(n_542),
.Y(n_823)
);

BUFx5_ASAP7_75t_L g824 ( 
.A(n_680),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_565),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_715),
.B(n_356),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_709),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_709),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_678),
.A2(n_566),
.B(n_571),
.C(n_570),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_577),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_603),
.B(n_567),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_643),
.B(n_287),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_717),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_694),
.A2(n_542),
.B1(n_550),
.B2(n_554),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_704),
.B(n_228),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_596),
.A2(n_352),
.B1(n_381),
.B2(n_375),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_624),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_651),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_616),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_626),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_625),
.B(n_555),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_649),
.B(n_356),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_633),
.B(n_555),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_659),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_684),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_610),
.B(n_268),
.C(n_258),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_592),
.B(n_228),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_622),
.B(n_567),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_596),
.A2(n_349),
.B1(n_346),
.B2(n_341),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_712),
.B(n_555),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_655),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_655),
.B(n_570),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_614),
.B(n_240),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_667),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_668),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_596),
.A2(n_322),
.B1(n_337),
.B2(n_240),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_656),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_693),
.A2(n_542),
.B(n_554),
.C(n_550),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_656),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_653),
.B(n_361),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_668),
.B(n_572),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_580),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_687),
.B(n_361),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_711),
.B(n_708),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_637),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_687),
.B(n_571),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_687),
.B(n_232),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_637),
.B(n_648),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_591),
.B(n_273),
.C(n_269),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_613),
.B(n_564),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_687),
.B(n_366),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_637),
.B(n_572),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_657),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_648),
.B(n_572),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_648),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_627),
.B(n_366),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_626),
.B(n_572),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_629),
.B(n_368),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_657),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_702),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_708),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_660),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_679),
.A2(n_612),
.B(n_602),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_766),
.B(n_623),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_863),
.B(n_623),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_733),
.A2(n_602),
.B(n_595),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_779),
.B(n_677),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_743),
.B(n_694),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_729),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_750),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_773),
.A2(n_601),
.B(n_593),
.C(n_609),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_768),
.B(n_806),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_768),
.B(n_677),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_792),
.B(n_619),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_781),
.A2(n_672),
.B(n_638),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_782),
.A2(n_602),
.B(n_595),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_729),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_750),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_763),
.B(n_635),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_782),
.A2(n_646),
.B(n_595),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_784),
.B(n_635),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_730),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_761),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_878),
.B(n_635),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_781),
.B(n_631),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_722),
.B(n_658),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_812),
.A2(n_672),
.B(n_220),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_820),
.B(n_575),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_799),
.A2(n_665),
.B(n_660),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_722),
.B(n_673),
.C(n_685),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_730),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_723),
.A2(n_688),
.B(n_646),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_762),
.B(n_707),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_865),
.Y(n_916)
);

CKINVDCx10_ASAP7_75t_R g917 ( 
.A(n_832),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_800),
.A2(n_696),
.B(n_681),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_SL g919 ( 
.A1(n_787),
.A2(n_340),
.B(n_319),
.C(n_321),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_838),
.B(n_735),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_799),
.A2(n_706),
.B(n_696),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_792),
.A2(n_672),
.B1(n_312),
.B2(n_371),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_738),
.B(n_673),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_377),
.B(n_338),
.C(n_333),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_812),
.A2(n_672),
.B(n_220),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_767),
.B(n_707),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_756),
.B(n_619),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_800),
.A2(n_713),
.B(n_706),
.Y(n_928)
);

OAI321xp33_ASAP7_75t_L g929 ( 
.A1(n_816),
.A2(n_835),
.A3(n_795),
.B1(n_793),
.B2(n_790),
.C(n_880),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_R g930 ( 
.A(n_737),
.B(n_236),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_767),
.B(n_707),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_774),
.B(n_253),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_724),
.B(n_564),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_756),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_774),
.A2(n_649),
.B1(n_714),
.B2(n_680),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_746),
.B(n_713),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_732),
.A2(n_688),
.B(n_646),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_758),
.A2(n_688),
.B(n_579),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_792),
.B(n_619),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_769),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_789),
.A2(n_599),
.B(n_597),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_825),
.B(n_232),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_794),
.B(n_285),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_736),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_728),
.B(n_802),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_851),
.A2(n_504),
.B(n_494),
.C(n_495),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_748),
.B(n_649),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_649),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_865),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_816),
.B(n_835),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_792),
.A2(n_343),
.B1(n_359),
.B2(n_380),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_739),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_847),
.B(n_861),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_877),
.A2(n_226),
.B(n_217),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_756),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_848),
.B(n_232),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_865),
.A2(n_649),
.B1(n_714),
.B2(n_680),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_853),
.A2(n_387),
.B(n_331),
.C(n_376),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_750),
.B(n_619),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_852),
.B(n_855),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_870),
.B(n_597),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_750),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_788),
.B(n_680),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_786),
.B(n_599),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_856),
.B(n_260),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_758),
.A2(n_579),
.B(n_577),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_759),
.A2(n_579),
.B(n_577),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_847),
.B(n_577),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_796),
.B(n_604),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_727),
.B(n_564),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_740),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_777),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_759),
.A2(n_579),
.B(n_577),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_770),
.A2(n_581),
.B(n_579),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_861),
.B(n_581),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_777),
.B(n_619),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_777),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_L g979 ( 
.A(n_788),
.B(n_680),
.Y(n_979)
);

AO21x1_ASAP7_75t_L g980 ( 
.A1(n_793),
.A2(n_605),
.B(n_604),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_770),
.A2(n_594),
.B(n_581),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_790),
.A2(n_295),
.B(n_239),
.C(n_237),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_741),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_882),
.B(n_606),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_734),
.A2(n_594),
.B(n_581),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_804),
.B(n_606),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_809),
.B(n_608),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_726),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_744),
.B(n_581),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_877),
.B(n_594),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_813),
.B(n_608),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_741),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_L g993 ( 
.A1(n_880),
.A2(n_226),
.B(n_217),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_760),
.A2(n_620),
.B(n_615),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_879),
.A2(n_617),
.B(n_594),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_879),
.A2(n_885),
.B(n_752),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_742),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_742),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_L g999 ( 
.A(n_846),
.B(n_372),
.C(n_368),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_765),
.A2(n_620),
.B(n_615),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_831),
.B(n_260),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_862),
.A2(n_617),
.B(n_594),
.Y(n_1002)
);

CKINVDCx11_ASAP7_75t_R g1003 ( 
.A(n_819),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_771),
.A2(n_650),
.B(n_645),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_811),
.A2(n_650),
.B(n_645),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_811),
.A2(n_634),
.B(n_621),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_869),
.A2(n_617),
.B(n_662),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_828),
.B(n_621),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_726),
.B(n_260),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_777),
.B(n_617),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_808),
.B(n_617),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_749),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_749),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_837),
.B(n_844),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_772),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_845),
.B(n_618),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_791),
.A2(n_829),
.B(n_857),
.C(n_854),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_817),
.B(n_618),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_868),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_840),
.A2(n_662),
.B(n_636),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_817),
.B(n_618),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_772),
.B(n_618),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_788),
.B(n_618),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_727),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_788),
.B(n_636),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_788),
.B(n_636),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_757),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_778),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_727),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_805),
.A2(n_495),
.B(n_494),
.C(n_502),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_817),
.B(n_805),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_821),
.B(n_636),
.Y(n_1033)
);

NAND2x1_ASAP7_75t_SL g1034 ( 
.A(n_864),
.B(n_207),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_821),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_815),
.B(n_369),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_814),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_840),
.A2(n_662),
.B(n_636),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_814),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_725),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_L g1041 ( 
.A(n_832),
.Y(n_1041)
);

O2A1O1Ixp5_ASAP7_75t_L g1042 ( 
.A1(n_826),
.A2(n_502),
.B(n_504),
.C(n_512),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_827),
.A2(n_512),
.B(n_511),
.C(n_506),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_731),
.A2(n_714),
.B1(n_680),
.B2(n_662),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_827),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_833),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_818),
.A2(n_385),
.B(n_295),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_826),
.A2(n_714),
.B(n_537),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_833),
.A2(n_511),
.B(n_506),
.C(n_505),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_864),
.B(n_662),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_871),
.B(n_572),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_872),
.A2(n_385),
.B(n_239),
.C(n_237),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_725),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_859),
.A2(n_714),
.B(n_537),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_751),
.A2(n_714),
.B(n_537),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_754),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_788),
.B(n_572),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_872),
.B(n_277),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_810),
.B(n_369),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_801),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_783),
.A2(n_511),
.B(n_506),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_745),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_755),
.A2(n_380),
.B1(n_372),
.B2(n_378),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_SL g1064 ( 
.A(n_950),
.B(n_780),
.C(n_776),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_936),
.A2(n_783),
.B(n_830),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_950),
.A2(n_785),
.B1(n_747),
.B2(n_753),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_953),
.B(n_801),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_918),
.A2(n_875),
.B(n_807),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_953),
.B(n_883),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_895),
.B(n_832),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_929),
.B(n_764),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_908),
.A2(n_797),
.B1(n_849),
.B2(n_836),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_908),
.A2(n_797),
.B(n_843),
.C(n_850),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1058),
.A2(n_797),
.B(n_841),
.C(n_876),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_930),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_890),
.A2(n_803),
.B(n_823),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_907),
.B(n_822),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_894),
.B(n_822),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_895),
.B(n_839),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_1039),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_SL g1082 ( 
.A1(n_923),
.A2(n_227),
.B1(n_231),
.B2(n_358),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1024),
.B(n_839),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_982),
.A2(n_798),
.B(n_873),
.C(n_866),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_891),
.Y(n_1085)
);

OA21x2_ASAP7_75t_L g1086 ( 
.A1(n_980),
.A2(n_834),
.B(n_881),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_905),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_934),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1024),
.B(n_858),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_913),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_889),
.B(n_785),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1029),
.B(n_858),
.Y(n_1092)
);

OAI22x1_ASAP7_75t_L g1093 ( 
.A1(n_923),
.A2(n_358),
.B1(n_360),
.B2(n_363),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_893),
.A2(n_884),
.B(n_881),
.C(n_874),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_945),
.A2(n_884),
.B(n_874),
.C(n_860),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_963),
.A2(n_979),
.B(n_996),
.Y(n_1096)
);

CKINVDCx8_ASAP7_75t_R g1097 ( 
.A(n_917),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_1052),
.B(n_360),
.C(n_390),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_901),
.A2(n_830),
.B(n_842),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_945),
.A2(n_873),
.B1(n_860),
.B2(n_389),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_932),
.B(n_942),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_903),
.A2(n_830),
.B(n_824),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_932),
.A2(n_378),
.B(n_383),
.C(n_389),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_990),
.A2(n_383),
.B1(n_293),
.B2(n_278),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_934),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_888),
.A2(n_824),
.B(n_572),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_897),
.A2(n_369),
.B1(n_284),
.B2(n_266),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_990),
.A2(n_351),
.B1(n_281),
.B2(n_286),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_956),
.B(n_290),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_914),
.A2(n_824),
.B(n_505),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_960),
.B(n_1014),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1015),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1017),
.A2(n_357),
.B(n_307),
.C(n_308),
.Y(n_1113)
);

CKINVDCx8_ASAP7_75t_R g1114 ( 
.A(n_988),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_937),
.A2(n_824),
.B(n_505),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1014),
.B(n_824),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_920),
.B(n_297),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_1052),
.B(n_363),
.C(n_388),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1023),
.A2(n_824),
.B(n_500),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1023),
.A2(n_500),
.B(n_497),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_SL g1121 ( 
.A(n_934),
.B(n_365),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_920),
.A2(n_266),
.B1(n_284),
.B2(n_537),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1029),
.B(n_78),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1056),
.B(n_302),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1025),
.A2(n_500),
.B(n_497),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1032),
.B(n_313),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_L g1127 ( 
.A1(n_912),
.A2(n_365),
.B1(n_388),
.B2(n_386),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_906),
.B(n_955),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1025),
.A2(n_497),
.B(n_537),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1015),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1026),
.A2(n_537),
.B(n_110),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1026),
.A2(n_537),
.B(n_111),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_982),
.A2(n_266),
.B(n_284),
.C(n_353),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_SL g1134 ( 
.A(n_1019),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1057),
.A2(n_91),
.B(n_79),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_954),
.A2(n_390),
.B1(n_386),
.B2(n_384),
.C(n_379),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_SL g1137 ( 
.A(n_886),
.B(n_384),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_997),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_969),
.B(n_344),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_969),
.B(n_327),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_930),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1031),
.A2(n_326),
.B1(n_317),
.B2(n_316),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_955),
.B(n_379),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_955),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_924),
.A2(n_18),
.B(n_20),
.C(n_22),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_905),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1050),
.A2(n_374),
.B1(n_370),
.B2(n_367),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_898),
.A2(n_902),
.B(n_947),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_976),
.A2(n_146),
.B(n_90),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_940),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_922),
.B(n_374),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_899),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_976),
.A2(n_140),
.B(n_96),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1031),
.B(n_370),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_955),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_951),
.B(n_367),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_910),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_964),
.B(n_190),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_916),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_999),
.A2(n_184),
.B1(n_183),
.B2(n_180),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_915),
.A2(n_176),
.B(n_163),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_926),
.A2(n_931),
.B(n_938),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1050),
.A2(n_159),
.B1(n_157),
.B2(n_147),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1059),
.B(n_20),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_SL g1166 ( 
.A1(n_943),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_904),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_909),
.A2(n_27),
.B(n_29),
.C(n_35),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1011),
.A2(n_139),
.B(n_138),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1037),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1011),
.A2(n_136),
.B(n_133),
.Y(n_1171)
);

XOR2x2_ASAP7_75t_SL g1172 ( 
.A(n_933),
.B(n_37),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_944),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1037),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_943),
.B(n_38),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_911),
.A2(n_126),
.B(n_125),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_975),
.A2(n_123),
.B(n_117),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_964),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_925),
.A2(n_989),
.B(n_993),
.C(n_1001),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_966),
.B(n_887),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_964),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_916),
.A2(n_80),
.B1(n_39),
.B2(n_40),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_981),
.A2(n_76),
.B(n_40),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1010),
.A2(n_38),
.B(n_41),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1062),
.B(n_44),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1010),
.A2(n_44),
.B(n_46),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1036),
.B(n_47),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_1003),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1062),
.B(n_49),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_989),
.A2(n_1016),
.B(n_1054),
.C(n_1055),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_952),
.B(n_49),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_978),
.B(n_51),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_972),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_978),
.B(n_52),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_983),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_992),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_949),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1047),
.B(n_60),
.C(n_66),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_949),
.B(n_67),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_933),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_978),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1016),
.A2(n_68),
.B(n_70),
.C(n_72),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1063),
.B(n_1012),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1013),
.B(n_1027),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1028),
.B(n_68),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1035),
.B(n_75),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1009),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1034),
.B(n_76),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1051),
.A2(n_1002),
.B(n_985),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1041),
.B(n_984),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_924),
.A2(n_961),
.B(n_1046),
.C(n_1041),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_958),
.B(n_1022),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1018),
.B(n_1021),
.Y(n_1214)
);

AOI221x1_ASAP7_75t_L g1215 ( 
.A1(n_1168),
.A2(n_967),
.B1(n_968),
.B2(n_974),
.C(n_1007),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1114),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1096),
.A2(n_928),
.B(n_1061),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1181),
.B(n_962),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1101),
.B(n_1060),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1151),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1085),
.Y(n_1221)
);

INVx5_ASAP7_75t_L g1222 ( 
.A(n_1105),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1163),
.A2(n_973),
.B(n_1053),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1210),
.A2(n_994),
.B(n_1004),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1083),
.Y(n_1225)
);

AOI221xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1168),
.A2(n_946),
.B1(n_1030),
.B2(n_987),
.C(n_970),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1097),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1088),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1149),
.A2(n_1053),
.B(n_1040),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1117),
.A2(n_948),
.B(n_1043),
.C(n_935),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1076),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_1175),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1065),
.A2(n_1040),
.B(n_1038),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1088),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1111),
.A2(n_978),
.B1(n_962),
.B2(n_1022),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1172),
.B(n_1060),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1072),
.A2(n_1179),
.B(n_1190),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1153),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1167),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1087),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1141),
.B(n_971),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1081),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1105),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1117),
.A2(n_1175),
.B(n_1064),
.C(n_1152),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1070),
.B(n_971),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1173),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1112),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1095),
.A2(n_995),
.A3(n_1033),
.B(n_1020),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1155),
.B(n_971),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1080),
.B(n_892),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1071),
.B(n_892),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1109),
.B(n_900),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1077),
.A2(n_921),
.B(n_1000),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1181),
.B(n_1068),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1113),
.A2(n_896),
.B(n_939),
.C(n_977),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1200),
.B(n_991),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1128),
.A2(n_986),
.B(n_1008),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1105),
.Y(n_1258)
);

NAND3x1_ASAP7_75t_L g1259 ( 
.A(n_1152),
.B(n_957),
.C(n_1044),
.Y(n_1259)
);

OAI22x1_ASAP7_75t_L g1260 ( 
.A1(n_1157),
.A2(n_959),
.B1(n_919),
.B2(n_965),
.Y(n_1260)
);

AOI221x1_ASAP7_75t_L g1261 ( 
.A1(n_1183),
.A2(n_941),
.B1(n_1006),
.B2(n_1005),
.C(n_1048),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1069),
.A2(n_1106),
.B(n_1110),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1207),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1130),
.B(n_959),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1157),
.A2(n_1049),
.B(n_927),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1074),
.A2(n_927),
.B(n_1042),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1126),
.B(n_1087),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1075),
.A2(n_1094),
.A3(n_1212),
.B(n_1099),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1193),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1116),
.A2(n_1067),
.B(n_1102),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_SL g1271 ( 
.A(n_1181),
.B(n_1188),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1204),
.A3(n_1080),
.B(n_1214),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1196),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1176),
.A2(n_1078),
.B(n_1214),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1123),
.B(n_1174),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1078),
.A2(n_1139),
.B(n_1140),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1120),
.A2(n_1125),
.B(n_1150),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1119),
.A2(n_1129),
.B(n_1177),
.Y(n_1278)
);

NAND3x1_ASAP7_75t_L g1279 ( 
.A(n_1187),
.B(n_1211),
.C(n_1185),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1121),
.A2(n_1071),
.B(n_1203),
.C(n_1206),
.Y(n_1280)
);

AOI21xp33_ASAP7_75t_L g1281 ( 
.A1(n_1133),
.A2(n_1104),
.B(n_1108),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1086),
.A2(n_1169),
.B(n_1171),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1079),
.B(n_1180),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1170),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1154),
.A2(n_1159),
.B(n_1203),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1084),
.A2(n_1204),
.B(n_1086),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1209),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1158),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1086),
.A2(n_1162),
.B(n_1186),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1068),
.B(n_1145),
.Y(n_1290)
);

AND2x6_ASAP7_75t_L g1291 ( 
.A(n_1213),
.B(n_1123),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1135),
.A2(n_1131),
.B(n_1132),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1090),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1205),
.A2(n_1206),
.A3(n_1127),
.B(n_1191),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1147),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1083),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1084),
.A2(n_1092),
.B(n_1089),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1202),
.A2(n_1103),
.B(n_1159),
.C(n_1194),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1205),
.A2(n_1184),
.A3(n_1164),
.B(n_1199),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1199),
.A2(n_1093),
.A3(n_1182),
.B(n_1189),
.Y(n_1300)
);

BUFx10_ASAP7_75t_L g1301 ( 
.A(n_1134),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1092),
.A2(n_1066),
.B(n_1091),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1073),
.A2(n_1066),
.B1(n_1100),
.B2(n_1107),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1134),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_SL g1305 ( 
.A(n_1105),
.B(n_1156),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1156),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1165),
.A2(n_1122),
.B(n_1107),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1192),
.A2(n_1194),
.B(n_1143),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1202),
.A2(n_1192),
.B(n_1144),
.C(n_1161),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1185),
.A2(n_1189),
.A3(n_1197),
.B(n_1138),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1147),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1156),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1160),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1160),
.B(n_1124),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1156),
.A2(n_1178),
.B(n_1145),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1201),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1146),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1178),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1208),
.A2(n_1146),
.B(n_1195),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1142),
.Y(n_1320)
);

OAI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1137),
.A2(n_1136),
.B(n_1198),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1148),
.A2(n_1098),
.A3(n_1118),
.B(n_1198),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1098),
.B(n_1118),
.C(n_1195),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1082),
.B(n_1166),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1096),
.A2(n_628),
.B(n_840),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1175),
.B(n_950),
.C(n_953),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1111),
.A2(n_950),
.B1(n_953),
.B2(n_945),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_L g1329 ( 
.A1(n_1117),
.A2(n_950),
.B(n_953),
.C(n_1058),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1085),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1151),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1095),
.A2(n_980),
.A3(n_1074),
.B(n_1075),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1101),
.B(n_950),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1117),
.A2(n_950),
.B(n_953),
.C(n_929),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1072),
.A2(n_950),
.B(n_953),
.Y(n_1337)
);

CKINVDCx8_ASAP7_75t_R g1338 ( 
.A(n_1151),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1085),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1151),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1163),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1096),
.A2(n_628),
.B(n_840),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1111),
.B(n_768),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1087),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1072),
.A2(n_950),
.B(n_953),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1095),
.A2(n_980),
.A3(n_1074),
.B(n_1075),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1096),
.A2(n_628),
.B(n_840),
.Y(n_1348)
);

AO32x2_ASAP7_75t_L g1349 ( 
.A1(n_1166),
.A2(n_1197),
.A3(n_1182),
.B1(n_1108),
.B2(n_1104),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1095),
.A2(n_980),
.A3(n_1074),
.B(n_1075),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1111),
.B(n_768),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1096),
.A2(n_628),
.B(n_840),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1095),
.A2(n_1163),
.B(n_980),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1072),
.A2(n_950),
.B(n_953),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1111),
.B(n_950),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_SL g1356 ( 
.A1(n_1179),
.A2(n_950),
.B(n_953),
.C(n_1168),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1168),
.A2(n_950),
.B1(n_982),
.B2(n_953),
.C(n_925),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1096),
.A2(n_628),
.B(n_840),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1072),
.A2(n_950),
.B(n_953),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1096),
.A2(n_1210),
.B(n_1149),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1085),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1111),
.A2(n_950),
.B1(n_953),
.B2(n_722),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1085),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1151),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1220),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1332),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1334),
.B(n_1232),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1363),
.A2(n_1327),
.B1(n_1244),
.B2(n_1320),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1324),
.A2(n_1327),
.B1(n_1303),
.B2(n_1323),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1221),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1340),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1355),
.B(n_1328),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1335),
.A2(n_1323),
.B(n_1321),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1228),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1238),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1328),
.A2(n_1343),
.B1(n_1351),
.B2(n_1354),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1232),
.B(n_1252),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1228),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1321),
.A2(n_1354),
.B1(n_1345),
.B2(n_1337),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1337),
.A2(n_1345),
.B1(n_1360),
.B2(n_1307),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1307),
.A2(n_1291),
.B1(n_1360),
.B2(n_1319),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1227),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1239),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1246),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1281),
.A2(n_1237),
.B1(n_1285),
.B2(n_1236),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1237),
.A2(n_1291),
.B1(n_1274),
.B2(n_1317),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1284),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1338),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1216),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1291),
.A2(n_1274),
.B1(n_1283),
.B2(n_1267),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1231),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1279),
.A2(n_1219),
.B1(n_1291),
.B2(n_1251),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1301),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1314),
.B(n_1256),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1253),
.A2(n_1348),
.B(n_1359),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1302),
.A2(n_1329),
.B1(n_1245),
.B2(n_1287),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1222),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1305),
.B(n_1222),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1263),
.Y(n_1401)
);

CKINVDCx6p67_ASAP7_75t_R g1402 ( 
.A(n_1242),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1275),
.A2(n_1249),
.B1(n_1259),
.B2(n_1241),
.Y(n_1403)
);

CKINVDCx8_ASAP7_75t_R g1404 ( 
.A(n_1304),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1365),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1222),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1275),
.A2(n_1240),
.B1(n_1295),
.B2(n_1362),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1275),
.A2(n_1240),
.B1(n_1295),
.B2(n_1339),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1276),
.A2(n_1356),
.B(n_1230),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1301),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1228),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1322),
.B(n_1294),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1269),
.A2(n_1273),
.B1(n_1364),
.B2(n_1331),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1311),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1293),
.A2(n_1313),
.B1(n_1344),
.B2(n_1308),
.Y(n_1415)
);

BUFx8_ASAP7_75t_L g1416 ( 
.A(n_1288),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1357),
.B(n_1280),
.Y(n_1417)
);

BUFx8_ASAP7_75t_L g1418 ( 
.A(n_1234),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1349),
.A2(n_1235),
.B1(n_1357),
.B2(n_1308),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1272),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1260),
.A2(n_1265),
.B1(n_1250),
.B2(n_1264),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1265),
.A2(n_1286),
.B1(n_1271),
.B2(n_1349),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1234),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1349),
.A2(n_1297),
.B1(n_1296),
.B2(n_1225),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1294),
.B(n_1300),
.Y(n_1425)
);

CKINVDCx6p67_ASAP7_75t_R g1426 ( 
.A(n_1234),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1243),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1225),
.A2(n_1296),
.B1(n_1322),
.B2(n_1292),
.Y(n_1428)
);

AND2x4_ASAP7_75t_SL g1429 ( 
.A(n_1243),
.B(n_1258),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1353),
.A2(n_1270),
.B1(n_1300),
.B2(n_1316),
.Y(n_1430)
);

INVx6_ASAP7_75t_L g1431 ( 
.A(n_1243),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1322),
.B(n_1294),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1353),
.A2(n_1300),
.B1(n_1282),
.B2(n_1277),
.Y(n_1433)
);

CKINVDCx6p67_ASAP7_75t_R g1434 ( 
.A(n_1312),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1277),
.A2(n_1266),
.B1(n_1223),
.B2(n_1224),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1272),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1258),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1318),
.A2(n_1218),
.B1(n_1290),
.B2(n_1254),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1258),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1306),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1309),
.A2(n_1298),
.B1(n_1299),
.B2(n_1342),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1299),
.A2(n_1352),
.B1(n_1325),
.B2(n_1289),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1261),
.A2(n_1215),
.B1(n_1257),
.B2(n_1299),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1272),
.B(n_1226),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1333),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1315),
.A2(n_1229),
.B1(n_1233),
.B2(n_1341),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1255),
.A2(n_1217),
.B1(n_1226),
.B2(n_1268),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1268),
.B(n_1350),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1333),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1278),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1326),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1333),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1347),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1347),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1248),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1248),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1330),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1336),
.A2(n_1346),
.B1(n_1358),
.B2(n_1361),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1347),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1262),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1350),
.A2(n_1248),
.B1(n_950),
.B2(n_1327),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1350),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1355),
.B(n_1334),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1221),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1324),
.A2(n_722),
.B1(n_908),
.B2(n_950),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1221),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1227),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_722),
.B2(n_908),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1216),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1227),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1327),
.A2(n_1363),
.B1(n_1324),
.B2(n_950),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1305),
.B(n_1181),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1327),
.A2(n_1363),
.B1(n_1324),
.B2(n_950),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1344),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1324),
.A2(n_722),
.B1(n_908),
.B2(n_950),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1324),
.A2(n_722),
.B1(n_908),
.B2(n_950),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1221),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1221),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1324),
.A2(n_722),
.B1(n_908),
.B2(n_950),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1305),
.B(n_1181),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1240),
.Y(n_1486)
);

CKINVDCx16_ASAP7_75t_R g1487 ( 
.A(n_1216),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1222),
.Y(n_1488)
);

BUFx8_ASAP7_75t_L g1489 ( 
.A(n_1332),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_722),
.B2(n_908),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1216),
.Y(n_1491)
);

INVx4_ASAP7_75t_SL g1492 ( 
.A(n_1291),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1327),
.A2(n_1363),
.B1(n_1324),
.B2(n_950),
.Y(n_1493)
);

AOI22x1_ASAP7_75t_L g1494 ( 
.A1(n_1337),
.A2(n_1354),
.B1(n_1360),
.B2(n_1345),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1222),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1222),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1324),
.A2(n_722),
.B1(n_908),
.B2(n_950),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_722),
.B2(n_908),
.Y(n_1499)
);

BUFx8_ASAP7_75t_L g1500 ( 
.A(n_1332),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1228),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1327),
.A2(n_950),
.B1(n_953),
.B2(n_908),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1227),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1221),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1492),
.B(n_1412),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1441),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1469),
.A2(n_1479),
.B1(n_1480),
.B2(n_1484),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1457),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1446),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1450),
.Y(n_1510)
);

INVxp33_ASAP7_75t_L g1511 ( 
.A(n_1388),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1472),
.A2(n_1490),
.B1(n_1499),
.B2(n_1494),
.Y(n_1512)
);

BUFx2_ASAP7_75t_SL g1513 ( 
.A(n_1399),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1486),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1455),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1425),
.B(n_1420),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1463),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1492),
.B(n_1432),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1405),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1420),
.B(n_1436),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1498),
.A2(n_1370),
.B1(n_1475),
.B2(n_1493),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1436),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1445),
.B(n_1462),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1449),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1367),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1464),
.B(n_1396),
.Y(n_1527)
);

AO21x2_ASAP7_75t_L g1528 ( 
.A1(n_1397),
.A2(n_1444),
.B(n_1447),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1371),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1451),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1376),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1462),
.B(n_1381),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1381),
.B(n_1454),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1475),
.A2(n_1477),
.B1(n_1493),
.B2(n_1466),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1456),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1459),
.A2(n_1443),
.B(n_1435),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1456),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1384),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1385),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1477),
.A2(n_1482),
.B1(n_1468),
.B2(n_1465),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1433),
.A2(n_1422),
.B(n_1409),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1444),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1417),
.B(n_1419),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1467),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1478),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1470),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1481),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1407),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1483),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1435),
.A2(n_1433),
.B(n_1461),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1458),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1380),
.B(n_1453),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1465),
.A2(n_1495),
.B(n_1466),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1460),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1399),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1415),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1407),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1372),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1468),
.B(n_1482),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1380),
.B(n_1369),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1415),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1399),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1495),
.A2(n_1502),
.B(n_1386),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1502),
.A2(n_1393),
.B1(n_1386),
.B2(n_1382),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1448),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1430),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1403),
.B(n_1400),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1378),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1430),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1428),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1391),
.A2(n_1368),
.B1(n_1377),
.B2(n_1398),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1489),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1424),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1391),
.A2(n_1377),
.B1(n_1398),
.B2(n_1408),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1422),
.A2(n_1387),
.B(n_1421),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1408),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1424),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1489),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1442),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1413),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1400),
.Y(n_1584)
);

CKINVDCx14_ASAP7_75t_R g1585 ( 
.A(n_1390),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1500),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1421),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1387),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1406),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1488),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1488),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1496),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1496),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1496),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1500),
.A2(n_1366),
.B1(n_1389),
.B2(n_1410),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1496),
.Y(n_1597)
);

INVx8_ASAP7_75t_L g1598 ( 
.A(n_1497),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1497),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1439),
.B(n_1437),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1476),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1402),
.A2(n_1487),
.B1(n_1395),
.B2(n_1491),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1366),
.A2(n_1416),
.B1(n_1394),
.B2(n_1401),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1476),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1485),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1485),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1438),
.B(n_1440),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1521),
.A2(n_1394),
.B1(n_1411),
.B2(n_1375),
.C(n_1473),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1560),
.B(n_1427),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1434),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1560),
.B(n_1375),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1508),
.B(n_1555),
.Y(n_1612)
);

AND2x4_ASAP7_75t_SL g1613 ( 
.A(n_1607),
.B(n_1392),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1514),
.B(n_1525),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_SL g1615 ( 
.A(n_1570),
.B(n_1411),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1526),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1527),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1534),
.A2(n_1503),
.B1(n_1474),
.B2(n_1429),
.C(n_1416),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1507),
.A2(n_1379),
.B1(n_1501),
.B2(n_1423),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1519),
.B(n_1471),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1536),
.A2(n_1431),
.B(n_1426),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1555),
.B(n_1431),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1585),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1511),
.B(n_1561),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1512),
.A2(n_1418),
.B(n_1379),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_R g1626 ( 
.A(n_1575),
.B(n_1383),
.Y(n_1626)
);

AND2x4_ASAP7_75t_SL g1627 ( 
.A(n_1607),
.B(n_1418),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1540),
.A2(n_1379),
.B1(n_1423),
.B2(n_1501),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1514),
.B(n_1404),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1553),
.B(n_1431),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1577),
.A2(n_1423),
.B1(n_1501),
.B2(n_1566),
.Y(n_1631)
);

NAND2xp33_ASAP7_75t_L g1632 ( 
.A(n_1563),
.B(n_1554),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_SL g1633 ( 
.A1(n_1567),
.A2(n_1574),
.B(n_1562),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1563),
.A2(n_1589),
.B1(n_1588),
.B2(n_1549),
.C(n_1579),
.Y(n_1634)
);

AO32x2_ASAP7_75t_L g1635 ( 
.A1(n_1565),
.A2(n_1523),
.A3(n_1516),
.B1(n_1568),
.B2(n_1542),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1586),
.A2(n_1582),
.B(n_1589),
.C(n_1588),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1549),
.A2(n_1579),
.B(n_1559),
.C(n_1582),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1551),
.A2(n_1542),
.B(n_1568),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1570),
.A2(n_1559),
.B1(n_1607),
.B2(n_1544),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1570),
.A2(n_1607),
.B1(n_1544),
.B2(n_1602),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1546),
.B(n_1557),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1551),
.A2(n_1569),
.B(n_1572),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1545),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1505),
.B(n_1518),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1583),
.A2(n_1607),
.B(n_1573),
.C(n_1570),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1545),
.Y(n_1648)
);

AO32x2_ASAP7_75t_L g1649 ( 
.A1(n_1565),
.A2(n_1516),
.A3(n_1520),
.B1(n_1580),
.B2(n_1576),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1599),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1528),
.A2(n_1537),
.B(n_1569),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1505),
.B(n_1518),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1578),
.A2(n_1532),
.B1(n_1603),
.B2(n_1596),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1532),
.A2(n_1578),
.B1(n_1573),
.B2(n_1576),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1524),
.B(n_1557),
.Y(n_1656)
);

AO32x2_ASAP7_75t_L g1657 ( 
.A1(n_1565),
.A2(n_1520),
.A3(n_1580),
.B1(n_1578),
.B2(n_1522),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1575),
.Y(n_1658)
);

INVxp67_ASAP7_75t_SL g1659 ( 
.A(n_1552),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1531),
.B(n_1538),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1661)
);

OAI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1558),
.A2(n_1564),
.B(n_1541),
.C(n_1572),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1587),
.A2(n_1581),
.B1(n_1575),
.B2(n_1505),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1547),
.B(n_1548),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1581),
.A2(n_1606),
.B(n_1605),
.C(n_1601),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1581),
.A2(n_1601),
.B(n_1606),
.C(n_1605),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1584),
.A2(n_1565),
.B1(n_1591),
.B2(n_1590),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1584),
.A2(n_1604),
.B(n_1595),
.C(n_1594),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1600),
.B(n_1550),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1543),
.B(n_1535),
.Y(n_1670)
);

INVx5_ASAP7_75t_L g1671 ( 
.A(n_1535),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_SL g1672 ( 
.A(n_1543),
.B(n_1513),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1509),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1635),
.B(n_1541),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1635),
.B(n_1541),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1649),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1673),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1639),
.A2(n_1604),
.B1(n_1556),
.B2(n_1590),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1644),
.B(n_1515),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1614),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1640),
.B(n_1515),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1664),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1632),
.B(n_1594),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1633),
.A2(n_1604),
.B1(n_1556),
.B2(n_1598),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1646),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1517),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1666),
.B(n_1537),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1640),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_R g1691 ( 
.A(n_1621),
.B(n_1530),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1657),
.B(n_1649),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1510),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1664),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1650),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1671),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1543),
.Y(n_1697)
);

INVxp33_ASAP7_75t_L g1698 ( 
.A(n_1638),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1643),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1627),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1654),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1651),
.B(n_1506),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1611),
.B(n_1593),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1668),
.B(n_1530),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1661),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1656),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1530),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1621),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1652),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1679),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1710),
.B(n_1612),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1682),
.B(n_1659),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1686),
.B(n_1653),
.C(n_1685),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1698),
.A2(n_1655),
.B(n_1641),
.Y(n_1715)
);

CKINVDCx12_ASAP7_75t_R g1716 ( 
.A(n_1697),
.Y(n_1716)
);

INVx5_ASAP7_75t_SL g1717 ( 
.A(n_1697),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1709),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1677),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1677),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1678),
.A2(n_1647),
.B(n_1615),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1656),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1683),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1636),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1703),
.B(n_1669),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1710),
.B(n_1672),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1680),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1699),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1617),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1699),
.B(n_1662),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1680),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1686),
.B(n_1637),
.C(n_1634),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1683),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1709),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1698),
.A2(n_1634),
.B1(n_1608),
.B2(n_1625),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1681),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1706),
.B(n_1662),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1681),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1695),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1685),
.A2(n_1642),
.B1(n_1631),
.B2(n_1608),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1681),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1707),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1700),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1695),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1688),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1687),
.Y(n_1747)
);

AND2x2_ASAP7_75t_SL g1748 ( 
.A(n_1676),
.B(n_1613),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1700),
.A2(n_1625),
.B1(n_1663),
.B2(n_1618),
.Y(n_1749)
);

AOI31xp33_ASAP7_75t_L g1750 ( 
.A1(n_1678),
.A2(n_1626),
.A3(n_1665),
.B(n_1618),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1688),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1688),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1676),
.A2(n_1631),
.B1(n_1609),
.B2(n_1611),
.C(n_1616),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1721),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1718),
.B(n_1676),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1743),
.B(n_1707),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1718),
.B(n_1692),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1719),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1684),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1697),
.Y(n_1761)
);

NAND2x1_ASAP7_75t_L g1762 ( 
.A(n_1722),
.B(n_1709),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1721),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1730),
.B(n_1623),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1720),
.Y(n_1765)
);

AND2x2_ASAP7_75t_SL g1766 ( 
.A(n_1748),
.B(n_1692),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1720),
.B(n_1684),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1728),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1728),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1735),
.B(n_1674),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1737),
.B(n_1674),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1732),
.B(n_1694),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1701),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1701),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1715),
.A2(n_1697),
.B1(n_1689),
.B2(n_1708),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1738),
.B(n_1701),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1737),
.B(n_1674),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1748),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1727),
.B(n_1697),
.Y(n_1780)
);

AND2x4_ASAP7_75t_SL g1781 ( 
.A(n_1744),
.B(n_1696),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1739),
.B(n_1742),
.Y(n_1782)
);

AND2x4_ASAP7_75t_SL g1783 ( 
.A(n_1744),
.B(n_1696),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1732),
.B(n_1694),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1739),
.B(n_1693),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1729),
.B(n_1704),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1693),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1725),
.B(n_1697),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1746),
.B(n_1751),
.Y(n_1790)
);

XNOR2xp5_ASAP7_75t_L g1791 ( 
.A(n_1749),
.B(n_1658),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1711),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1746),
.B(n_1675),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1751),
.B(n_1675),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1724),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1758),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1758),
.Y(n_1797)
);

NAND2xp67_ASAP7_75t_L g1798 ( 
.A(n_1781),
.B(n_1622),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1765),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1779),
.B(n_1727),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1765),
.Y(n_1801)
);

OR2x6_ASAP7_75t_L g1802 ( 
.A(n_1762),
.B(n_1722),
.Y(n_1802)
);

O2A1O1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1762),
.A2(n_1750),
.B(n_1733),
.C(n_1714),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1781),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1779),
.Y(n_1805)
);

NAND2x1_ASAP7_75t_L g1806 ( 
.A(n_1780),
.B(n_1727),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1766),
.B(n_1717),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1782),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1755),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1782),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1766),
.B(n_1717),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1768),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1782),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1773),
.B(n_1752),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1791),
.A2(n_1776),
.B(n_1736),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1768),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1773),
.B(n_1752),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1791),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1790),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1766),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1761),
.B(n_1717),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1744),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1790),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1769),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1781),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1759),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1764),
.A2(n_1741),
.B1(n_1753),
.B2(n_1665),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1775),
.B(n_1740),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1780),
.B(n_1620),
.Y(n_1831)
);

NOR2x1p5_ASAP7_75t_SL g1832 ( 
.A(n_1754),
.B(n_1702),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1759),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1775),
.B(n_1745),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1767),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1761),
.B(n_1717),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1767),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1756),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1777),
.A2(n_1700),
.B1(n_1624),
.B2(n_1723),
.C(n_1734),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1777),
.B(n_1713),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1772),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1805),
.B(n_1815),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1806),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1796),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1821),
.B(n_1780),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1846)
);

OAI32xp33_ASAP7_75t_L g1847 ( 
.A1(n_1829),
.A2(n_1755),
.A3(n_1757),
.B1(n_1760),
.B2(n_1770),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1821),
.B(n_1783),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1796),
.Y(n_1849)
);

INVx2_ASAP7_75t_SL g1850 ( 
.A(n_1806),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1801),
.Y(n_1851)
);

NAND3xp33_ASAP7_75t_L g1852 ( 
.A(n_1802),
.B(n_1609),
.C(n_1756),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1801),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1838),
.B(n_1774),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1809),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1818),
.B(n_1831),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1812),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1827),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1840),
.B(n_1755),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1807),
.B(n_1789),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1839),
.B(n_1789),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1807),
.B(n_1757),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1811),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1822),
.B(n_1629),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1830),
.B(n_1788),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1808),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1834),
.B(n_1788),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1812),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1816),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1840),
.B(n_1785),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1811),
.B(n_1757),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1816),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1808),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1810),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1800),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1835),
.B(n_1785),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1800),
.B(n_1726),
.Y(n_1877)
);

INVxp33_ASAP7_75t_L g1878 ( 
.A(n_1822),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1837),
.B(n_1787),
.Y(n_1879)
);

XOR2x2_ASAP7_75t_L g1880 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1855),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1846),
.A2(n_1836),
.B(n_1804),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1858),
.B(n_1804),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1875),
.B(n_1828),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1863),
.B(n_1828),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1878),
.A2(n_1802),
.B1(n_1852),
.B2(n_1848),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1844),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1877),
.B(n_1824),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1856),
.B(n_1802),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1843),
.A2(n_1802),
.B(n_1824),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1843),
.A2(n_1824),
.B1(n_1716),
.B2(n_1689),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1850),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1844),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1847),
.A2(n_1760),
.B1(n_1690),
.B2(n_1770),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1847),
.A2(n_1850),
.B(n_1861),
.C(n_1854),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1864),
.B(n_1833),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1862),
.B(n_1824),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1862),
.A2(n_1783),
.B1(n_1675),
.B2(n_1697),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1845),
.A2(n_1832),
.B(n_1760),
.C(n_1783),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1845),
.A2(n_1716),
.B1(n_1841),
.B2(n_1833),
.Y(n_1900)
);

AOI221x1_ASAP7_75t_L g1901 ( 
.A1(n_1849),
.A2(n_1826),
.B1(n_1797),
.B2(n_1823),
.C(n_1799),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1860),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1860),
.A2(n_1841),
.B1(n_1691),
.B2(n_1770),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1849),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1851),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1851),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1897),
.B(n_1871),
.Y(n_1907)
);

AOI21xp33_ASAP7_75t_L g1908 ( 
.A1(n_1889),
.A2(n_1871),
.B(n_1866),
.Y(n_1908)
);

OAI321xp33_ASAP7_75t_L g1909 ( 
.A1(n_1886),
.A2(n_1859),
.A3(n_1876),
.B1(n_1874),
.B2(n_1873),
.C(n_1866),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1902),
.B(n_1859),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1892),
.B(n_1873),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1881),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1881),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1883),
.B(n_1865),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1857),
.C(n_1853),
.Y(n_1915)
);

OAI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1895),
.A2(n_1867),
.B(n_1874),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1904),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_L g1918 ( 
.A(n_1894),
.B(n_1857),
.C(n_1853),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1901),
.B(n_1868),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1904),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1882),
.A2(n_1872),
.B(n_1869),
.C(n_1868),
.Y(n_1921)
);

OAI21xp33_ASAP7_75t_L g1922 ( 
.A1(n_1880),
.A2(n_1876),
.B(n_1798),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1870),
.Y(n_1923)
);

AOI211x1_ASAP7_75t_L g1924 ( 
.A1(n_1885),
.A2(n_1872),
.B(n_1869),
.C(n_1826),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_L g1925 ( 
.A(n_1890),
.B(n_1879),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1887),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1893),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1913),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1912),
.B(n_1896),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1907),
.B(n_1888),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1917),
.Y(n_1931)
);

OAI321xp33_ASAP7_75t_L g1932 ( 
.A1(n_1916),
.A2(n_1891),
.A3(n_1900),
.B1(n_1899),
.B2(n_1903),
.C(n_1884),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1919),
.Y(n_1933)
);

OAI21xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1925),
.A2(n_1898),
.B(n_1905),
.Y(n_1934)
);

XNOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1919),
.B(n_1906),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1920),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1919),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1910),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1907),
.B(n_1810),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1928),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1933),
.A2(n_1915),
.B1(n_1918),
.B2(n_1914),
.Y(n_1941)
);

NOR4xp25_ASAP7_75t_L g1942 ( 
.A(n_1933),
.B(n_1909),
.C(n_1921),
.D(n_1927),
.Y(n_1942)
);

AOI211xp5_ASAP7_75t_L g1943 ( 
.A1(n_1932),
.A2(n_1908),
.B(n_1922),
.C(n_1923),
.Y(n_1943)
);

NOR3xp33_ASAP7_75t_L g1944 ( 
.A(n_1929),
.B(n_1923),
.C(n_1926),
.Y(n_1944)
);

NAND4xp75_ASAP7_75t_L g1945 ( 
.A(n_1937),
.B(n_1924),
.C(n_1911),
.D(n_1910),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1939),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1937),
.B(n_1934),
.C(n_1936),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1930),
.B(n_1938),
.Y(n_1948)
);

AOI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1931),
.A2(n_1911),
.B1(n_1879),
.B2(n_1870),
.C(n_1825),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1935),
.A2(n_1813),
.B1(n_1825),
.B2(n_1820),
.Y(n_1950)
);

NAND4xp25_ASAP7_75t_L g1951 ( 
.A(n_1943),
.B(n_1930),
.C(n_1938),
.D(n_1939),
.Y(n_1951)
);

AOI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1942),
.A2(n_1941),
.B1(n_1947),
.B2(n_1944),
.C(n_1940),
.Y(n_1952)
);

AOI21xp33_ASAP7_75t_SL g1953 ( 
.A1(n_1946),
.A2(n_1935),
.B(n_1817),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1945),
.Y(n_1954)
);

XNOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1948),
.B(n_1610),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1950),
.A2(n_1819),
.B(n_1813),
.Y(n_1956)
);

O2A1O1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1949),
.A2(n_1820),
.B(n_1819),
.C(n_1814),
.Y(n_1957)
);

AOI211xp5_ASAP7_75t_L g1958 ( 
.A1(n_1952),
.A2(n_1619),
.B(n_1628),
.C(n_1814),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1954),
.A2(n_1619),
.B1(n_1691),
.B2(n_1628),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1953),
.A2(n_1817),
.B(n_1667),
.C(n_1630),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1951),
.A2(n_1787),
.B(n_1690),
.C(n_1795),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1955),
.A2(n_1772),
.B(n_1784),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1957),
.A2(n_1832),
.B(n_1690),
.C(n_1795),
.Y(n_1963)
);

AOI211xp5_ASAP7_75t_L g1964 ( 
.A1(n_1956),
.A2(n_1754),
.B(n_1795),
.C(n_1763),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1958),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1960),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1959),
.B(n_1754),
.Y(n_1967)
);

NAND4xp75_ASAP7_75t_L g1968 ( 
.A(n_1962),
.B(n_1705),
.C(n_1794),
.D(n_1793),
.Y(n_1968)
);

AO22x1_ASAP7_75t_L g1969 ( 
.A1(n_1961),
.A2(n_1705),
.B1(n_1763),
.B2(n_1747),
.Y(n_1969)
);

XOR2x2_ASAP7_75t_L g1970 ( 
.A(n_1964),
.B(n_1963),
.Y(n_1970)
);

OAI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1966),
.A2(n_1763),
.B1(n_1734),
.B2(n_1747),
.C(n_1696),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1965),
.B(n_1712),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1969),
.B(n_1724),
.C(n_1784),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1970),
.B(n_1967),
.Y(n_1974)
);

AO22x2_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1972),
.B1(n_1967),
.B2(n_1968),
.Y(n_1975)
);

OAI22x1_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1973),
.B1(n_1971),
.B2(n_1696),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1976),
.Y(n_1977)
);

XNOR2xp5_ASAP7_75t_L g1978 ( 
.A(n_1976),
.B(n_1798),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1977),
.B(n_1597),
.Y(n_1979)
);

AOI22x1_ASAP7_75t_L g1980 ( 
.A1(n_1978),
.A2(n_1696),
.B1(n_1792),
.B2(n_1556),
.Y(n_1980)
);

INVx4_ASAP7_75t_L g1981 ( 
.A(n_1979),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1980),
.A2(n_1792),
.B(n_1786),
.Y(n_1982)
);

NAND2x1p5_ASAP7_75t_L g1983 ( 
.A(n_1981),
.B(n_1597),
.Y(n_1983)
);

AOI21xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1983),
.A2(n_1982),
.B(n_1598),
.Y(n_1984)
);

OAI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1786),
.B1(n_1556),
.B2(n_1723),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1794),
.B1(n_1793),
.B2(n_1778),
.C(n_1771),
.Y(n_1986)
);

AOI211xp5_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1556),
.B(n_1597),
.C(n_1592),
.Y(n_1987)
);


endmodule