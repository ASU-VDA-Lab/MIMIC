module fake_ariane_1416_n_1237 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1237);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1237;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_209;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_174;
wire n_275;
wire n_204;
wire n_1232;
wire n_1211;
wire n_996;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_38),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_1),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_44),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_23),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_16),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_80),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_63),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_55),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_107),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_135),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_118),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_31),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

BUFx8_ASAP7_75t_SL g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_51),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_22),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_34),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_58),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_114),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_155),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_126),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_26),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_59),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_30),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_37),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_93),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_213),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_184),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_177),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_174),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_177),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

BUFx2_ASAP7_75t_R g255 ( 
.A(n_178),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_187),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_189),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_194),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_251),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_237),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_253),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_239),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_242),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_255),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_233),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_242),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_242),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_233),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_253),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_284),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_292),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_293),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_270),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_273),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_273),
.B(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_276),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_307),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_310),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_295),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_298),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_278),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_263),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_279),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_272),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_280),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_300),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_300),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_281),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_269),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_331),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_361),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_290),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_286),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_287),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_328),
.B(n_267),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_286),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_323),
.B(n_268),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

BUFx8_ASAP7_75t_SL g388 ( 
.A(n_322),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_286),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_302),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_308),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_229),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_317),
.B(n_182),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_318),
.B(n_178),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_317),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_319),
.B(n_180),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_225),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_355),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_340),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_388),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_340),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_373),
.A2(n_323),
.B1(n_350),
.B2(n_352),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_360),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_407),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_368),
.A2(n_357),
.B(n_356),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_388),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_335),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_387),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_360),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_395),
.A2(n_398),
.B1(n_368),
.B2(n_397),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_404),
.A2(n_344),
.B1(n_339),
.B2(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_349),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_321),
.B1(n_333),
.B2(n_362),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_301),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_351),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_365),
.B(n_354),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

NOR2x1_ASAP7_75t_L g445 ( 
.A(n_367),
.B(n_179),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_364),
.B(n_275),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_379),
.A2(n_176),
.B(n_183),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_180),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_371),
.A2(n_223),
.B1(n_188),
.B2(n_191),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_372),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_215),
.B(n_176),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_375),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_181),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_383),
.A2(n_181),
.B1(n_227),
.B2(n_231),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_374),
.B(n_275),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_374),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_399),
.A2(n_196),
.B(n_192),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_380),
.B(n_227),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_370),
.Y(n_475)
);

CKINVDCx11_ASAP7_75t_R g476 ( 
.A(n_370),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_390),
.A2(n_231),
.B1(n_223),
.B2(n_205),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_374),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_275),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_401),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_390),
.B(n_197),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_402),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_402),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_386),
.A2(n_214),
.B1(n_206),
.B2(n_207),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_403),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_411),
.B(n_377),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_476),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_426),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_423),
.B(n_377),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_426),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_403),
.C(n_396),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_476),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_415),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_403),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_422),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_415),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_422),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_R g521 ( 
.A(n_475),
.B(n_403),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_447),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_475),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_433),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_438),
.B(n_378),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_446),
.B(n_378),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_487),
.B(n_378),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_427),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_429),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_R g533 ( 
.A(n_417),
.B(n_378),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_418),
.A2(n_190),
.B1(n_199),
.B2(n_216),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_490),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_490),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_417),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_487),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_416),
.B(n_275),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_489),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_489),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_416),
.B(n_0),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_437),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_416),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_430),
.B(n_0),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_468),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_431),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_430),
.B(n_434),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_430),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_486),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_486),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_486),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_441),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_378),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_470),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_465),
.C(n_455),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_532),
.B(n_462),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_502),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_509),
.A2(n_436),
.B1(n_479),
.B2(n_451),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_556),
.B(n_445),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_515),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_533),
.B(n_483),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_516),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_533),
.B(n_470),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_517),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_520),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_525),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_555),
.B(n_410),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_523),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_507),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_524),
.B(n_454),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_534),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_534),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_535),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_443),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_539),
.B(n_443),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_512),
.B(n_518),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_535),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_521),
.B(n_425),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_521),
.B(n_428),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_541),
.B(n_428),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_563),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_511),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_567),
.A2(n_550),
.B1(n_526),
.B2(n_469),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_571),
.A2(n_526),
.B1(n_503),
.B2(n_550),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_568),
.B(n_504),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_522),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_585),
.B(n_527),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_584),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_569),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_595),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_578),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_505),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_569),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_548),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_588),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_593),
.B(n_500),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_584),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_596),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_600),
.B(n_553),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_572),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_598),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_589),
.B(n_506),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_596),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_586),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_577),
.B(n_513),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_603),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_569),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_603),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_583),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_605),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_589),
.B(n_497),
.C(n_477),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_601),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_605),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_574),
.B(n_552),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_601),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_573),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_576),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_601),
.B(n_513),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_565),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_583),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_576),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_583),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_604),
.B(n_513),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_557),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_581),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_590),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_582),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_572),
.A2(n_469),
.B1(n_554),
.B2(n_540),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_590),
.B(n_546),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_583),
.B(n_547),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_582),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_542),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_587),
.B(n_545),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_591),
.B(n_443),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_604),
.B(n_531),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_587),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_587),
.B(n_558),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_592),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_592),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_592),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_587),
.B(n_513),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_572),
.B(n_559),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_602),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_602),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_572),
.B(n_529),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_602),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_572),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_566),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_566),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_566),
.B(n_560),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_570),
.B(n_529),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_570),
.B(n_544),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_615),
.B(n_508),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_629),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_634),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_630),
.B(n_531),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_637),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_641),
.Y(n_695)
);

INVxp33_ASAP7_75t_L g696 ( 
.A(n_664),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_625),
.B(n_530),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_617),
.B(n_622),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_633),
.B(n_538),
.Y(n_699)
);

BUFx8_ASAP7_75t_L g700 ( 
.A(n_674),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_609),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_653),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_656),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_659),
.Y(n_707)
);

XOR2xp5_ASAP7_75t_L g708 ( 
.A(n_611),
.B(n_503),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_661),
.Y(n_709)
);

XOR2xp5_ASAP7_75t_L g710 ( 
.A(n_621),
.B(n_501),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_687),
.B(n_549),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_665),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_618),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_673),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_627),
.Y(n_715)
);

INVx4_ASAP7_75t_SL g716 ( 
.A(n_640),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_677),
.Y(n_717)
);

BUFx5_ASAP7_75t_L g718 ( 
.A(n_606),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_619),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_625),
.B(n_543),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_608),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_614),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_614),
.Y(n_723)
);

XOR2xp5_ASAP7_75t_L g724 ( 
.A(n_668),
.B(n_510),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_626),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_610),
.B(n_519),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_626),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_635),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_673),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_635),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_613),
.B(n_549),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_613),
.B(n_549),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_660),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_610),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_660),
.Y(n_737)
);

BUFx6f_ASAP7_75t_SL g738 ( 
.A(n_651),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_667),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_642),
.A2(n_463),
.B(n_564),
.Y(n_740)
);

BUFx6f_ASAP7_75t_SL g741 ( 
.A(n_671),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_667),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_613),
.B(n_679),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_672),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_672),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_675),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_682),
.A2(n_528),
.B(n_544),
.Y(n_747)
);

CKINVDCx14_ASAP7_75t_R g748 ( 
.A(n_640),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_669),
.B(n_549),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_675),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_676),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_680),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_654),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_680),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_681),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_683),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_685),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_646),
.Y(n_759)
);

INVxp33_ASAP7_75t_SL g760 ( 
.A(n_658),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_639),
.Y(n_761)
);

AOI21x1_ASAP7_75t_L g762 ( 
.A1(n_678),
.A2(n_461),
.B(n_469),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_645),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_624),
.B(n_570),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_638),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_639),
.Y(n_766)
);

XOR2x2_ASAP7_75t_L g767 ( 
.A(n_645),
.B(n_1),
.Y(n_767)
);

BUFx5_ASAP7_75t_L g768 ( 
.A(n_606),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_684),
.B(n_452),
.Y(n_769)
);

XNOR2x2_ASAP7_75t_L g770 ( 
.A(n_663),
.B(n_472),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_688),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_740),
.B(n_678),
.C(n_650),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_736),
.B(n_720),
.Y(n_773)
);

AND2x4_ASAP7_75t_SL g774 ( 
.A(n_714),
.B(n_658),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_719),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_713),
.B(n_606),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_726),
.B(n_607),
.C(n_662),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_738),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_715),
.B(n_606),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_708),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_697),
.B(n_640),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_696),
.B(n_682),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_698),
.B(n_606),
.Y(n_784)
);

BUFx8_ASAP7_75t_L g785 ( 
.A(n_738),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_691),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_695),
.B(n_612),
.Y(n_787)
);

BUFx8_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_694),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_2),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_731),
.B(n_623),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_765),
.B(n_616),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_702),
.B(n_631),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_703),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_705),
.B(n_631),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_770),
.A2(n_607),
.B(n_662),
.C(n_636),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_693),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_706),
.B(n_620),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_763),
.B(n_2),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_701),
.A2(n_684),
.B1(n_754),
.B2(n_710),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_707),
.B(n_620),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_712),
.B(n_643),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_704),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_709),
.B(n_643),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_747),
.B(n_684),
.Y(n_805)
);

INVx8_ASAP7_75t_L g806 ( 
.A(n_741),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_699),
.B(n_652),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_716),
.B(n_623),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_749),
.B(n_652),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_700),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_759),
.B(n_655),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_748),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_757),
.B(n_655),
.Y(n_813)
);

BUFx6f_ASAP7_75t_SL g814 ( 
.A(n_765),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_717),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_743),
.B(n_682),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_716),
.B(n_623),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_758),
.B(n_666),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_724),
.B(n_3),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_743),
.B(n_623),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_718),
.B(n_632),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_700),
.B(n_3),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_733),
.B(n_666),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_718),
.B(n_632),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_734),
.B(n_671),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_765),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_764),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_764),
.B(n_671),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_711),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_4),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_761),
.B(n_624),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_766),
.B(n_624),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_721),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_771),
.B(n_638),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_767),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_722),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_723),
.B(n_636),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_725),
.B(n_638),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_718),
.B(n_632),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_727),
.B(n_638),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_782),
.Y(n_842)
);

AO22x2_ASAP7_75t_L g843 ( 
.A1(n_777),
.A2(n_730),
.B1(n_729),
.B2(n_728),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_794),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_786),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_815),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_803),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_789),
.Y(n_848)
);

OAI221xp5_ASAP7_75t_L g849 ( 
.A1(n_777),
.A2(n_230),
.B1(n_226),
.B2(n_222),
.C(n_215),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_773),
.B(n_775),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_810),
.Y(n_851)
);

NAND2x1p5_ASAP7_75t_L g852 ( 
.A(n_808),
.B(n_616),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_828),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_787),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_834),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_778),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_812),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_837),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_793),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_772),
.B(n_718),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_795),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_817),
.B(n_616),
.Y(n_862)
);

OAI221xp5_ASAP7_75t_L g863 ( 
.A1(n_796),
.A2(n_215),
.B1(n_632),
.B2(n_670),
.C(n_737),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_791),
.B(n_616),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_800),
.A2(n_732),
.B1(n_739),
.B2(n_735),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_798),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_816),
.B(n_742),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_838),
.Y(n_868)
);

AO22x2_ASAP7_75t_L g869 ( 
.A1(n_783),
.A2(n_744),
.B1(n_746),
.B2(n_745),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_816),
.B(n_750),
.Y(n_870)
);

AO22x2_ASAP7_75t_L g871 ( 
.A1(n_776),
.A2(n_751),
.B1(n_753),
.B2(n_752),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_801),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_804),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_826),
.B(n_649),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_779),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_806),
.B(n_688),
.Y(n_878)
);

AO22x2_ASAP7_75t_L g879 ( 
.A1(n_784),
.A2(n_755),
.B1(n_756),
.B2(n_689),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_781),
.B(n_4),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_5),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_778),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_827),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_807),
.B(n_718),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_831),
.A2(n_768),
.B1(n_769),
.B2(n_688),
.Y(n_887)
);

AO22x2_ASAP7_75t_L g888 ( 
.A1(n_827),
.A2(n_689),
.B1(n_580),
.B2(n_575),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_811),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_799),
.A2(n_768),
.B1(n_657),
.B2(n_649),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_797),
.B(n_768),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_790),
.A2(n_657),
.B1(n_561),
.B2(n_544),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_841),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_816),
.B(n_835),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_809),
.B(n_823),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_836),
.A2(n_768),
.B1(n_410),
.B2(n_686),
.Y(n_896)
);

NAND2x1p5_ASAP7_75t_L g897 ( 
.A(n_826),
.B(n_686),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_825),
.B(n_768),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_805),
.A2(n_410),
.B1(n_686),
.B2(n_474),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_832),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_780),
.B(n_762),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_821),
.B(n_686),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_805),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_785),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_805),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_774),
.B(n_461),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_819),
.A2(n_203),
.B(n_202),
.C(n_221),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_785),
.Y(n_908)
);

NAND2x1_ASAP7_75t_L g909 ( 
.A(n_833),
.B(n_561),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_829),
.B(n_5),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_830),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_824),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_840),
.Y(n_913)
);

BUFx8_ASAP7_75t_L g914 ( 
.A(n_814),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_788),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_854),
.B(n_866),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_872),
.B(n_792),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_915),
.A2(n_452),
.B(n_575),
.Y(n_919)
);

CKINVDCx6p67_ASAP7_75t_R g920 ( 
.A(n_856),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_883),
.A2(n_792),
.B(n_410),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_873),
.B(n_806),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_863),
.A2(n_806),
.B1(n_452),
.B2(n_580),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_876),
.B(n_6),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_860),
.A2(n_814),
.B(n_561),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_849),
.A2(n_410),
.B(n_478),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_909),
.A2(n_561),
.B(n_544),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_916),
.A2(n_580),
.B(n_575),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_857),
.B(n_428),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_882),
.B(n_889),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_904),
.B(n_6),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_887),
.A2(n_466),
.B1(n_428),
.B2(n_440),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_853),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_843),
.A2(n_424),
.B(n_457),
.Y(n_935)
);

OR2x6_ASAP7_75t_SL g936 ( 
.A(n_850),
.B(n_457),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_871),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_842),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_843),
.A2(n_480),
.B(n_471),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_859),
.B(n_7),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_912),
.B(n_440),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_885),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_910),
.A2(n_466),
.B(n_481),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_879),
.A2(n_886),
.B(n_891),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_901),
.A2(n_439),
.B(n_414),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_914),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_861),
.B(n_8),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_890),
.A2(n_439),
.B1(n_456),
.B2(n_414),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_913),
.A2(n_439),
.B(n_495),
.C(n_414),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_879),
.A2(n_480),
.B(n_471),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_851),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_914),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_892),
.A2(n_485),
.B(n_484),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_908),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_865),
.A2(n_485),
.B(n_484),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_900),
.Y(n_956)
);

CKINVDCx10_ASAP7_75t_R g957 ( 
.A(n_881),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_844),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_865),
.A2(n_898),
.B(n_871),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_874),
.B(n_877),
.Y(n_960)
);

CKINVDCx6p67_ASAP7_75t_R g961 ( 
.A(n_906),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_896),
.A2(n_466),
.B1(n_464),
.B2(n_458),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_868),
.A2(n_899),
.B1(n_870),
.B2(n_867),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_894),
.B(n_440),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_858),
.B(n_893),
.C(n_911),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_895),
.B(n_8),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_864),
.A2(n_460),
.B1(n_456),
.B2(n_473),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_878),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_846),
.Y(n_969)
);

AO21x1_ASAP7_75t_L g970 ( 
.A1(n_847),
.A2(n_491),
.B(n_482),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_880),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_959),
.B(n_944),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_954),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_951),
.B(n_894),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_929),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_937),
.Y(n_976)
);

BUFx10_ASAP7_75t_L g977 ( 
.A(n_932),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_956),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_920),
.B(n_907),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_943),
.A2(n_933),
.B1(n_948),
.B2(n_965),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_942),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_917),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_931),
.B(n_885),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_930),
.B(n_204),
.C(n_200),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_952),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_921),
.A2(n_905),
.B(n_903),
.C(n_867),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_SL g987 ( 
.A(n_966),
.B(n_875),
.C(n_862),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_942),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_929),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_929),
.Y(n_990)
);

INVx5_ASAP7_75t_L g991 ( 
.A(n_946),
.Y(n_991)
);

AND3x2_ASAP7_75t_SL g992 ( 
.A(n_957),
.B(n_855),
.C(n_845),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_SL g993 ( 
.A(n_951),
.B(n_968),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_934),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_938),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_958),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_951),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_969),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_971),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_968),
.B(n_870),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_924),
.B(n_940),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_947),
.B(n_918),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_961),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_928),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_936),
.B(n_848),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_957),
.B(n_9),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_922),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_970),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_960),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_968),
.B(n_852),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_962),
.B(n_878),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_945),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_925),
.B(n_210),
.C(n_209),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_941),
.B(n_963),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_964),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_949),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_919),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_967),
.B(n_902),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_950),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_927),
.B(n_869),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_935),
.B(n_869),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_926),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_939),
.B(n_897),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_923),
.B(n_9),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_953),
.B(n_219),
.C(n_217),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_R g1026 ( 
.A(n_955),
.B(n_10),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_952),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_956),
.B(n_888),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_917),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_920),
.B(n_10),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_917),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_929),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_965),
.B(n_11),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_929),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_990),
.B(n_11),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_976),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1003),
.B(n_13),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_972),
.A2(n_494),
.B(n_493),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1023),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_978),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_1034),
.B(n_448),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_975),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_1006),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_993),
.B(n_203),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_985),
.A2(n_496),
.B(n_488),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_975),
.B(n_448),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_991),
.B(n_1033),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_982),
.B(n_13),
.Y(n_1049)
);

AO22x1_ASAP7_75t_L g1050 ( 
.A1(n_1033),
.A2(n_467),
.B1(n_464),
.B2(n_458),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_997),
.B(n_14),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1021),
.A2(n_499),
.B(n_498),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1040),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1040),
.Y(n_1056)
);

CKINVDCx8_ASAP7_75t_R g1057 ( 
.A(n_1042),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_991),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_1037),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1048),
.A2(n_1030),
.B(n_979),
.C(n_980),
.Y(n_1060)
);

BUFx8_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

AO221x2_ASAP7_75t_L g1062 ( 
.A1(n_1044),
.A2(n_992),
.B1(n_977),
.B2(n_1001),
.C(n_991),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1049),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_1042),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_1042),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_1035),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1039),
.A2(n_1027),
.B1(n_1016),
.B2(n_1008),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1052),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1035),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1036),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1047),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1050),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_1041),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1045),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1045),
.A2(n_1024),
.B1(n_1022),
.B2(n_1019),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1038),
.B(n_1029),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1047),
.B(n_1034),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_1067),
.A2(n_1017),
.B(n_1028),
.C(n_1015),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1058),
.B(n_1034),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1059),
.B(n_1031),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_1058),
.B(n_987),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1055),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1072),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1064),
.B(n_973),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1082),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1062),
.B1(n_1068),
.B2(n_1066),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1084),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1087),
.A2(n_1078),
.B(n_1060),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_1088),
.B(n_1066),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1090),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1089),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1094),
.B(n_1086),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1093),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1095),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1096),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1096),
.B(n_1079),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1100),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_1099),
.B(n_1097),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1101),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1102),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_1098),
.Y(n_1105)
);

NAND4xp25_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_1081),
.C(n_1069),
.D(n_1060),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_1106),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_1083),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1108),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1107),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1109),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1109),
.A2(n_1062),
.B1(n_1054),
.B2(n_1070),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1110),
.B(n_1062),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_1063),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1112),
.Y(n_1116)
);

OAI31xp33_ASAP7_75t_L g1117 ( 
.A1(n_1114),
.A2(n_1116),
.A3(n_1115),
.B(n_1065),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1114),
.B(n_1061),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1118),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1117),
.B(n_1070),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1120),
.B(n_1080),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_1061),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1122),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1121),
.B(n_977),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1124),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1123),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1126),
.A2(n_1125),
.B1(n_1057),
.B2(n_1032),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_L g1128 ( 
.A(n_1126),
.B(n_975),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1128),
.B(n_1127),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1128),
.Y(n_1130)
);

OAI32xp33_ASAP7_75t_L g1131 ( 
.A1(n_1127),
.A2(n_1073),
.A3(n_1074),
.B1(n_1072),
.B2(n_1077),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1130),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1129),
.B(n_203),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_1075),
.B(n_1032),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1133),
.B(n_14),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_1134),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1136),
.B(n_989),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_15),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1139),
.A2(n_203),
.B(n_989),
.C(n_1032),
.Y(n_1141)
);

NOR4xp75_ASAP7_75t_SL g1142 ( 
.A(n_1140),
.B(n_1076),
.C(n_1002),
.D(n_17),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1141),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1142),
.B(n_15),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1144),
.B(n_16),
.Y(n_1145)
);

INVxp67_ASAP7_75t_SL g1146 ( 
.A(n_1143),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_SL g1147 ( 
.A(n_1146),
.B(n_1075),
.C(n_1053),
.D(n_19),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1071),
.C(n_17),
.Y(n_1148)
);

NAND4xp25_ASAP7_75t_L g1149 ( 
.A(n_1145),
.B(n_18),
.C(n_19),
.D(n_20),
.Y(n_1149)
);

AOI211xp5_ASAP7_75t_L g1150 ( 
.A1(n_1149),
.A2(n_989),
.B(n_21),
.C(n_23),
.Y(n_1150)
);

AOI211xp5_ASAP7_75t_L g1151 ( 
.A1(n_1148),
.A2(n_18),
.B(n_21),
.C(n_24),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1147),
.B(n_272),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1152),
.Y(n_1153)
);

OAI31xp33_ASAP7_75t_SL g1154 ( 
.A1(n_1151),
.A2(n_1053),
.A3(n_25),
.B(n_26),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_1150),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1154),
.A2(n_1000),
.B1(n_272),
.B2(n_309),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1155),
.A2(n_984),
.B1(n_999),
.B2(n_1007),
.C(n_1013),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1156),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1158),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1157),
.A2(n_309),
.B1(n_1000),
.B2(n_988),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1159),
.A2(n_1047),
.B1(n_981),
.B2(n_988),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1160),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_1162),
.B(n_1025),
.C(n_981),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1161),
.B(n_309),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1164),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1163),
.B(n_24),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1164),
.Y(n_1167)
);

OAI222xp33_ASAP7_75t_L g1168 ( 
.A1(n_1166),
.A2(n_1167),
.B1(n_1165),
.B2(n_28),
.C1(n_29),
.C2(n_31),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1167),
.Y(n_1169)
);

NAND4xp25_ASAP7_75t_L g1170 ( 
.A(n_1166),
.B(n_25),
.C(n_27),
.D(n_28),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1169),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1168),
.A2(n_1010),
.B(n_27),
.Y(n_1172)
);

INVxp33_ASAP7_75t_L g1173 ( 
.A(n_1171),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1172),
.B(n_1170),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1173),
.B(n_974),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1174),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1176),
.B(n_1000),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1175),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1178),
.A2(n_29),
.B1(n_1000),
.B2(n_986),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1177),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1180),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_SL g1182 ( 
.A(n_1179),
.B(n_32),
.C(n_33),
.Y(n_1182)
);

AO22x2_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1182),
.A2(n_1014),
.B1(n_42),
.B2(n_43),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1181),
.A2(n_1011),
.B1(n_1020),
.B2(n_47),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1185),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1183),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1184),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1188),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_1186),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1189),
.A2(n_1187),
.B(n_1005),
.C(n_1011),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1190),
.A2(n_1011),
.B1(n_1018),
.B2(n_1012),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1192),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1191),
.A2(n_1011),
.B(n_983),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1192),
.A2(n_41),
.B(n_45),
.Y(n_1195)
);

OAI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1195),
.A2(n_1009),
.B1(n_56),
.B2(n_57),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1194),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1196),
.A2(n_62),
.B(n_64),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1198),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1197),
.A2(n_70),
.B(n_71),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1201),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1199),
.A2(n_1026),
.B(n_73),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1200),
.A2(n_72),
.B(n_74),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1201),
.A2(n_75),
.B(n_76),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1201),
.A2(n_77),
.B(n_78),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1201),
.A2(n_79),
.B(n_81),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1201),
.B(n_82),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1201),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1199),
.B(n_83),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1201),
.B(n_84),
.C(n_85),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1201),
.B(n_86),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1201),
.A2(n_87),
.B(n_88),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1201),
.A2(n_89),
.B(n_90),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1211),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1208),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1212),
.A2(n_1210),
.B1(n_1202),
.B2(n_1209),
.Y(n_1217)
);

AOI222xp33_ASAP7_75t_L g1218 ( 
.A1(n_1205),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.C1(n_105),
.C2(n_108),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1206),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1207),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_1220)
);

OAI221xp5_ASAP7_75t_R g1221 ( 
.A1(n_1213),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.C(n_121),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1214),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1203),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1217),
.A2(n_1204),
.B(n_131),
.Y(n_1224)
);

OAI222xp33_ASAP7_75t_L g1225 ( 
.A1(n_1219),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.C1(n_134),
.C2(n_137),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1221),
.A2(n_139),
.B(n_141),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1220),
.A2(n_998),
.B(n_995),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1218),
.A2(n_996),
.B(n_1004),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1216),
.A2(n_142),
.B(n_143),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_L g1230 ( 
.A1(n_1225),
.A2(n_1222),
.B1(n_1215),
.B2(n_1223),
.C(n_148),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1227),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.C(n_149),
.Y(n_1231)
);

AOI221x1_ASAP7_75t_L g1232 ( 
.A1(n_1229),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.C(n_156),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1224),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.C(n_161),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_1226),
.B1(n_1228),
.B2(n_166),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1234),
.A2(n_1231),
.B1(n_1232),
.B2(n_1230),
.Y(n_1235)
);

AOI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_162),
.B(n_164),
.C(n_167),
.Y(n_1236)
);

AOI211xp5_ASAP7_75t_L g1237 ( 
.A1(n_1236),
.A2(n_169),
.B(n_171),
.C(n_173),
.Y(n_1237)
);


endmodule