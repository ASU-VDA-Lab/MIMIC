module fake_jpeg_6693_n_86 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_58),
.B1(n_45),
.B2(n_37),
.Y(n_65)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_0),
.Y(n_56)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_52),
.B1(n_42),
.B2(n_49),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_47),
.A3(n_43),
.B1(n_51),
.B2(n_48),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_63),
.B1(n_64),
.B2(n_50),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_46),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_74),
.C(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_36),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_59),
.B1(n_13),
.B2(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_12),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_15),
.B(n_16),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_20),
.B(n_21),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_23),
.C(n_26),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_28),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_32),
.Y(n_86)
);


endmodule