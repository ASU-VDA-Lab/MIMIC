module fake_jpeg_24841_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_300;
wire n_294;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_247;
wire n_87;
wire n_46;
wire n_157;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_44),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_31),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_27),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_0),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_25),
.B1(n_30),
.B2(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_30),
.B1(n_18),
.B2(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_67),
.Y(n_109)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_75),
.Y(n_84)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_30),
.B1(n_38),
.B2(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_31),
.B1(n_18),
.B2(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_31),
.B1(n_18),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_77),
.B1(n_37),
.B2(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_19),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_20),
.Y(n_72)
);

OR2x2_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_76),
.Y(n_112)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_19),
.B1(n_37),
.B2(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_76),
.A2(n_42),
.B(n_27),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_1),
.C(n_2),
.Y(n_140)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_82),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_28),
.B1(n_27),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_104),
.B1(n_56),
.B2(n_54),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_90),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_15),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_3),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_92),
.B1(n_100),
.B2(n_90),
.Y(n_118)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_96),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_105),
.Y(n_139)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_108),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_22),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_115),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_34),
.B1(n_22),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_116),
.B1(n_74),
.B2(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_29),
.B1(n_34),
.B2(n_21),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_26),
.B1(n_1),
.B2(n_0),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_26),
.B(n_60),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_94),
.C(n_80),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_89),
.B1(n_88),
.B2(n_97),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_131),
.B1(n_110),
.B2(n_107),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_68),
.B1(n_73),
.B2(n_26),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_145),
.B1(n_11),
.B2(n_13),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_1),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_140),
.B(n_10),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_81),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_149),
.B1(n_113),
.B2(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_144),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_143),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_86),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_155),
.B(n_159),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_112),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_154),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_164),
.B(n_126),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_112),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_91),
.B1(n_81),
.B2(n_97),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_125),
.B1(n_127),
.B2(n_124),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_81),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_177),
.C(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_161),
.B(n_163),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_106),
.B1(n_88),
.B2(n_89),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_125),
.B1(n_146),
.B2(n_123),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_174),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_9),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_170),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_145),
.B(n_140),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_11),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.Y(n_209)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_137),
.B1(n_149),
.B2(n_119),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_11),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_17),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_198),
.B(n_201),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_192),
.B1(n_205),
.B2(n_155),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_156),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_144),
.B(n_121),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_191),
.B(n_204),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_133),
.B(n_142),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_167),
.B1(n_174),
.B2(n_166),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_120),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_199),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_123),
.B(n_129),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_141),
.B(n_15),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_14),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_14),
.B(n_15),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_16),
.B1(n_17),
.B2(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_175),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_182),
.C(n_183),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_219),
.C(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_161),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_191),
.C(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_178),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_193),
.B1(n_205),
.B2(n_201),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_180),
.C(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_195),
.B1(n_189),
.B2(n_194),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_173),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_186),
.C(n_208),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_246),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_236),
.B1(n_225),
.B2(n_231),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_192),
.B1(n_185),
.B2(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_184),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_211),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_250),
.B1(n_210),
.B2(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_247),
.C(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_204),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_218),
.C(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_212),
.B(n_222),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_233),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_208),
.B1(n_184),
.B2(n_157),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_257),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_231),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_222),
.B(n_213),
.C(n_225),
.D(n_218),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_261),
.C(n_265),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_250),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_223),
.B(n_220),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_260),
.A2(n_266),
.B(n_263),
.Y(n_271)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_266),
.B1(n_245),
.B2(n_240),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_246),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_247),
.C(n_242),
.Y(n_265)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_271),
.A2(n_259),
.B(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_234),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_265),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_274),
.B(n_270),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_258),
.B1(n_261),
.B2(n_254),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_279),
.C(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_293),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_300),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_294),
.CI(n_292),
.CON(n_303),
.SN(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_296),
.B(n_299),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_302),
.Y(n_306)
);


endmodule