module fake_jpeg_14014_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_8),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_2),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_3),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_25),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_19),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_38),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_74),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_11),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_12),
.Y(n_118)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_22),
.B1(n_21),
.B2(n_30),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_77),
.A2(n_98),
.B1(n_107),
.B2(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_83),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_25),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_42),
.B1(n_30),
.B2(n_24),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_90),
.B1(n_92),
.B2(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_42),
.B1(n_21),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_24),
.B1(n_21),
.B2(n_27),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_40),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_95),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_97),
.B(n_101),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_22),
.B1(n_24),
.B2(n_36),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_17),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_35),
.B1(n_34),
.B2(n_19),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_37),
.B1(n_17),
.B2(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_34),
.B1(n_3),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_83),
.B1(n_84),
.B2(n_116),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_34),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_13),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_14),
.B(n_15),
.C(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_144),
.Y(n_167)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_137),
.Y(n_177)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_40),
.Y(n_132)
);

OR2x6_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_80),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_93),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g187 ( 
.A(n_134),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_28),
.B(n_5),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_109),
.C(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_3),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_90),
.A2(n_60),
.B1(n_72),
.B2(n_28),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_153),
.B1(n_158),
.B2(n_120),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_152),
.B1(n_134),
.B2(n_141),
.Y(n_171)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_80),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_79),
.A2(n_13),
.B1(n_106),
.B2(n_112),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_95),
.A2(n_91),
.B1(n_100),
.B2(n_76),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_163),
.B1(n_142),
.B2(n_151),
.Y(n_196)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_85),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_109),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

CKINVDCx10_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_102),
.B1(n_76),
.B2(n_88),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_164),
.A2(n_188),
.B(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_166),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_123),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_85),
.B1(n_88),
.B2(n_78),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_126),
.A2(n_78),
.B1(n_120),
.B2(n_80),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_126),
.A2(n_147),
.B1(n_141),
.B2(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_141),
.C(n_144),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_129),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_122),
.B(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_124),
.B(n_133),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_197),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_128),
.B(n_145),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_159),
.B(n_132),
.C(n_156),
.D(n_149),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_201),
.A2(n_206),
.B(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_230),
.C(n_185),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_139),
.B(n_152),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_160),
.B1(n_157),
.B2(n_136),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_234)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_227),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_149),
.B(n_131),
.C(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_167),
.B(n_131),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_221),
.B(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_168),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_199),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_224),
.B(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_187),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_173),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_222),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_245),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_165),
.B1(n_174),
.B2(n_200),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_243),
.B1(n_244),
.B2(n_203),
.Y(n_267)
);

AOI32xp33_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_165),
.A3(n_174),
.B1(n_173),
.B2(n_184),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_207),
.B(n_214),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_178),
.B1(n_200),
.B2(n_194),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_178),
.B1(n_209),
.B2(n_216),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_231),
.B1(n_202),
.B2(n_224),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_202),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_251),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_204),
.A2(n_210),
.B1(n_206),
.B2(n_223),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_230),
.B1(n_221),
.B2(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_214),
.B1(n_201),
.B2(n_203),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_261),
.A2(n_267),
.B1(n_268),
.B2(n_274),
.Y(n_294)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_271),
.Y(n_291)
);

INVx2_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_219),
.B1(n_201),
.B2(n_205),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_240),
.C(n_255),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_235),
.B(n_220),
.CI(n_219),
.CON(n_271),
.SN(n_271)
);

OR2x2_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_220),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_281),
.B(n_239),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_211),
.B1(n_208),
.B2(n_212),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_279),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_280),
.B1(n_282),
.B2(n_260),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_247),
.B(n_249),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_249),
.B(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_240),
.C(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_253),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_236),
.C(n_271),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_297),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_253),
.B1(n_257),
.B2(n_251),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_275),
.B1(n_261),
.B2(n_272),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_246),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_265),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_242),
.B1(n_259),
.B2(n_234),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_238),
.C(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_217),
.B1(n_278),
.B2(n_280),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_263),
.B1(n_264),
.B2(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_270),
.B1(n_273),
.B2(n_282),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_266),
.B(n_265),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_287),
.B(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_293),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_284),
.C(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_288),
.C(n_297),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_286),
.C(n_294),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_301),
.C(n_303),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_289),
.B(n_290),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_309),
.A2(n_276),
.B(n_300),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_313),
.B1(n_306),
.B2(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_327),
.Y(n_336)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_332),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_306),
.C(n_310),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_319),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_318),
.B(n_315),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_314),
.B(n_320),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_302),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_333),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_340),
.B(n_341),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_338),
.C(n_336),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_342),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_343),
.C(n_326),
.Y(n_345)
);

AOI31xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_325),
.A3(n_328),
.B(n_323),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_323),
.Y(n_347)
);


endmodule