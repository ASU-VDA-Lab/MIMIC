module fake_aes_6955_n_754 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_754);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_754;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_105;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_102;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g83 ( .A(n_2), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_43), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_48), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_74), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_29), .Y(n_89) );
BUFx10_ASAP7_75t_L g90 ( .A(n_75), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_45), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_49), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_46), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_71), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_77), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_59), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_78), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_68), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_33), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_73), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_18), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_79), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_37), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_55), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_22), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_22), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_80), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_4), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_1), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_36), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_40), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_2), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_52), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_10), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_24), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_64), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_21), .Y(n_125) );
CKINVDCx14_ASAP7_75t_R g126 ( .A(n_53), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_17), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_1), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_57), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_39), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_62), .Y(n_131) );
INVxp33_ASAP7_75t_L g132 ( .A(n_60), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_23), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_101), .B(n_0), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_85), .B(n_0), .Y(n_137) );
NAND2x1_ASAP7_75t_L g138 ( .A(n_101), .B(n_3), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g139 ( .A(n_104), .B(n_30), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_101), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_103), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
BUFx8_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_83), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_103), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
NOR2xp33_ASAP7_75t_SL g152 ( .A(n_98), .B(n_31), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_117), .B(n_4), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_86), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_83), .B(n_5), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_90), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_88), .B(n_5), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_88), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_107), .B(n_6), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_87), .B(n_7), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_107), .B(n_7), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_132), .B(n_9), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_89), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_91), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_108), .B(n_10), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_92), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_92), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_93), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_96), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_96), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_99), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_108), .B(n_11), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_99), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_109), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_137), .B(n_116), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_168), .B(n_109), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_142), .B(n_100), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_142), .B(n_126), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_135), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
NAND3x1_ASAP7_75t_L g192 ( .A(n_137), .B(n_133), .C(n_110), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
OR2x2_ASAP7_75t_SL g199 ( .A(n_141), .B(n_133), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_146), .B(n_110), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_146), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_146), .B(n_122), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_136), .B(n_127), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_134), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_160), .B(n_127), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_153), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_140), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_146), .B(n_100), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_168), .B(n_131), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_150), .B(n_120), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_150), .B(n_94), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_150), .B(n_125), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_138), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_158), .B(n_130), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_139), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_158), .B(n_131), .Y(n_231) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_138), .B(n_115), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_158), .B(n_125), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_168), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_168), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_158), .B(n_114), .Y(n_237) );
NAND3x1_ASAP7_75t_L g238 ( .A(n_165), .B(n_111), .C(n_115), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_163), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_179), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_139), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_163), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_160), .B(n_119), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_143), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_241), .A2(n_230), .B1(n_226), .B2(n_224), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_204), .B(n_165), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_195), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_234), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_241), .A2(n_165), .B1(n_178), .B2(n_176), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_220), .Y(n_253) );
AND2x6_ASAP7_75t_SL g254 ( .A(n_182), .B(n_144), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_211), .B(n_222), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_211), .B(n_166), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_178), .B1(n_166), .B2(n_176), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_235), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_236), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_230), .B(n_179), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_244), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_182), .B(n_162), .Y(n_267) );
OAI21xp33_ASAP7_75t_L g268 ( .A1(n_245), .A2(n_156), .B(n_177), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_182), .B(n_162), .Y(n_269) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_230), .B(n_152), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_186), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_225), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_222), .B(n_167), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_186), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_239), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_182), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_189), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_181), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_190), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_239), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_238), .B(n_139), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_246), .B(n_152), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_186), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_194), .Y(n_288) );
AND2x6_ASAP7_75t_L g289 ( .A(n_197), .B(n_179), .Y(n_289) );
BUFx2_ASAP7_75t_R g290 ( .A(n_214), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_201), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_208), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_198), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_213), .B(n_143), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_200), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_184), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_203), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_184), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_226), .A2(n_167), .B1(n_171), .B2(n_179), .Y(n_299) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_208), .B(n_97), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_206), .Y(n_301) );
AOI22xp5_ASAP7_75t_SL g302 ( .A1(n_216), .A2(n_128), .B1(n_121), .B2(n_113), .Y(n_302) );
BUFx8_ASAP7_75t_L g303 ( .A(n_201), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_226), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_205), .B(n_143), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_188), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_219), .B(n_171), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_191), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_188), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_201), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_212), .Y(n_312) );
BUFx8_ASAP7_75t_L g313 ( .A(n_224), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_191), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_224), .B(n_143), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_233), .B(n_155), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_191), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_233), .B(n_144), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_232), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_260), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_250), .B(n_199), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_276), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_315), .A2(n_187), .B(n_202), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_276), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_318), .B(n_233), .Y(n_325) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_319), .B(n_278), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_271), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_277), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_302), .A2(n_223), .B1(n_215), .B2(n_185), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_318), .A2(n_238), .B1(n_192), .B2(n_231), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_319), .B(n_202), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_279), .Y(n_335) );
INVx5_ASAP7_75t_L g336 ( .A(n_260), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_294), .A2(n_229), .B(n_237), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_279), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_251), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_278), .B(n_183), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_271), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_247), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_300), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_247), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_310), .B(n_183), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_262), .A2(n_217), .B(n_192), .Y(n_348) );
AO32x2_ASAP7_75t_L g349 ( .A1(n_291), .A2(n_139), .A3(n_232), .B1(n_199), .B2(n_170), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_252), .A2(n_177), .B1(n_164), .B2(n_161), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_284), .A2(n_217), .B1(n_159), .B2(n_164), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_318), .B(n_156), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_260), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
BUFx8_ASAP7_75t_SL g356 ( .A(n_284), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_257), .B(n_159), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_300), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_258), .B(n_161), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_273), .B(n_169), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_292), .B(n_169), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_253), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_251), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_253), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_267), .A2(n_116), .B1(n_112), .B2(n_106), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_264), .B(n_155), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_289), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_255), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_261), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_274), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_260), .Y(n_373) );
INVx5_ASAP7_75t_L g374 ( .A(n_289), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_274), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_284), .A2(n_155), .B1(n_157), .B2(n_175), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_305), .A2(n_180), .B(n_193), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_374), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_333), .B(n_367), .C(n_352), .Y(n_380) );
CKINVDCx16_ASAP7_75t_R g381 ( .A(n_355), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_321), .A2(n_267), .B1(n_269), .B2(n_284), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_374), .B(n_287), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_350), .B(n_267), .Y(n_384) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_374), .B(n_269), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_350), .B(n_269), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_355), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_321), .A2(n_325), .B1(n_353), .B2(n_362), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_374), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_377), .A2(n_285), .B(n_264), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_325), .A2(n_311), .B1(n_291), .B2(n_270), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_353), .A2(n_311), .B1(n_270), .B2(n_304), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_333), .A2(n_259), .B1(n_248), .B2(n_264), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_346), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_304), .B1(n_289), .B2(n_268), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_357), .B(n_307), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_359), .B(n_254), .Y(n_400) );
AND2x6_ASAP7_75t_L g401 ( .A(n_334), .B(n_280), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_359), .A2(n_289), .B1(n_249), .B2(n_281), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
NAND3x1_ASAP7_75t_L g404 ( .A(n_356), .B(n_290), .C(n_118), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_376), .A2(n_293), .B1(n_282), .B2(n_312), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_289), .B1(n_280), .B2(n_282), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_340), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_336), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_361), .A2(n_289), .B1(n_281), .B2(n_312), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_365), .A2(n_293), .B1(n_295), .B2(n_301), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_345), .B(n_295), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_365), .A2(n_301), .B1(n_297), .B2(n_317), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_400), .A2(n_358), .B1(n_329), .B2(n_351), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_398), .B(n_360), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g416 ( .A1(n_406), .A2(n_348), .B(n_337), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_394), .A2(n_370), .B1(n_366), .B2(n_363), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_398), .B(n_338), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_388), .A2(n_363), .B1(n_366), .B2(n_370), .C1(n_297), .C2(n_324), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_412), .A2(n_347), .B1(n_341), .B2(n_334), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_406), .A2(n_323), .B(n_287), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_408), .A2(n_368), .B(n_340), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_378), .B(n_364), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_384), .A2(n_347), .B1(n_341), .B2(n_334), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_384), .A2(n_347), .B1(n_341), .B2(n_334), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_385), .B(n_368), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_380), .A2(n_368), .B1(n_341), .B2(n_331), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g429 ( .A1(n_401), .A2(n_368), .B1(n_369), .B2(n_347), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_378), .B(n_364), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_331), .B1(n_335), .B2(n_322), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_384), .A2(n_335), .B1(n_322), .B2(n_324), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_386), .A2(n_330), .B1(n_339), .B2(n_326), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_397), .A2(n_371), .B1(n_369), .B2(n_316), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_382), .A2(n_299), .B1(n_326), .B2(n_330), .C(n_339), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_386), .A2(n_375), .B1(n_342), .B2(n_372), .Y(n_436) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_391), .B(n_395), .C(n_405), .D(n_404), .Y(n_437) );
OAI21x1_ASAP7_75t_L g438 ( .A1(n_390), .A2(n_371), .B(n_372), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_386), .A2(n_375), .B1(n_372), .B2(n_327), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_411), .A2(n_157), .B1(n_175), .B2(n_255), .C(n_256), .Y(n_440) );
AOI22x1_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_320), .B1(n_354), .B2(n_343), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_391), .A2(n_157), .B1(n_175), .B2(n_256), .C(n_147), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_401), .A2(n_336), .B1(n_373), .B2(n_349), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_438), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_427), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_438), .A2(n_390), .B(n_395), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_415), .A2(n_381), .B1(n_397), .B2(n_387), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_420), .A2(n_386), .B1(n_401), .B2(n_392), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_420), .A2(n_401), .B1(n_404), .B2(n_393), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_430), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_414), .A2(n_413), .B1(n_396), .B2(n_402), .C(n_410), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_419), .A2(n_405), .B1(n_401), .B2(n_385), .C1(n_407), .C2(n_408), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
OAI221xp5_ASAP7_75t_SL g454 ( .A1(n_437), .A2(n_154), .B1(n_151), .B2(n_147), .C(n_145), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_427), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_421), .A2(n_401), .B1(n_409), .B2(n_327), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_437), .A2(n_129), .B(n_124), .C(n_154), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_424), .B(n_349), .Y(n_459) );
OAI221xp5_ASAP7_75t_SL g460 ( .A1(n_428), .A2(n_145), .B1(n_151), .B2(n_409), .C(n_111), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_443), .A2(n_123), .B(n_118), .C(n_119), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_434), .A2(n_123), .A3(n_148), .B1(n_149), .B2(n_349), .B3(n_193), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_418), .A2(n_409), .B1(n_401), .B2(n_399), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_425), .B(n_379), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_428), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_426), .A2(n_375), .B1(n_328), .B2(n_342), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_435), .A2(n_403), .A3(n_262), .B(n_263), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_427), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_441), .A2(n_403), .B1(n_399), .B2(n_389), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_423), .Y(n_473) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_422), .A2(n_148), .B(n_149), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_431), .B(n_432), .C(n_433), .D(n_442), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_429), .B(n_349), .Y(n_476) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_441), .B(n_399), .Y(n_477) );
AOI211xp5_ASAP7_75t_SL g478 ( .A1(n_440), .A2(n_379), .B(n_389), .C(n_349), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_436), .B(n_399), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_444), .Y(n_481) );
OAI33xp33_ASAP7_75t_L g482 ( .A1(n_447), .A2(n_148), .A3(n_149), .B1(n_180), .B2(n_14), .B3(n_15), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_449), .A2(n_389), .B1(n_379), .B2(n_403), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_453), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_463), .B(n_163), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_452), .A2(n_170), .B1(n_174), .B2(n_172), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_449), .B(n_210), .C(n_12), .D(n_13), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_450), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_454), .A2(n_172), .B1(n_174), .B2(n_170), .C(n_389), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_454), .A2(n_170), .B1(n_172), .B2(n_174), .C(n_379), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_448), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_463), .B(n_170), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
AND2x4_ASAP7_75t_SL g498 ( .A(n_445), .B(n_320), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_458), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_458), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_458), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_457), .B(n_102), .C(n_105), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_457), .A2(n_174), .B1(n_172), .B2(n_170), .C(n_263), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_475), .A2(n_174), .B1(n_172), .B2(n_170), .C(n_265), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_463), .B(n_172), .Y(n_505) );
AOI33xp33_ASAP7_75t_L g506 ( .A1(n_476), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_19), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_459), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_452), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_471), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_480), .B(n_466), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_465), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_476), .B(n_470), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_466), .B(n_172), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_465), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_174), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g517 ( .A1(n_478), .A2(n_174), .B(n_210), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_444), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_467), .B(n_16), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_475), .A2(n_373), .B1(n_342), .B2(n_327), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_467), .B(n_19), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_470), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_455), .B(n_20), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_462), .A2(n_265), .B1(n_243), .B2(n_242), .C(n_261), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_451), .A2(n_328), .B1(n_336), .B2(n_383), .C(n_194), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_445), .B(n_20), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_455), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_455), .B(n_21), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_455), .B(n_23), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_455), .B(n_336), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_507), .B(n_445), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_484), .B(n_445), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_490), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_498), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_513), .B(n_473), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_508), .B(n_455), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_513), .B(n_478), .Y(n_539) );
OAI211xp5_ASAP7_75t_SL g540 ( .A1(n_506), .A2(n_469), .B(n_451), .C(n_456), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
NAND4xp25_ASAP7_75t_SL g542 ( .A(n_506), .B(n_461), .C(n_469), .D(n_477), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_525), .B(n_479), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_498), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_491), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_528), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_487), .B(n_473), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_532), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_532), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_512), .B(n_479), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_528), .Y(n_551) );
AND4x1_ASAP7_75t_L g552 ( .A(n_482), .B(n_462), .C(n_477), .D(n_468), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_525), .B(n_479), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_515), .B(n_464), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_530), .B(n_464), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_499), .B(n_461), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
AND2x2_ASAP7_75t_SL g559 ( .A(n_530), .B(n_531), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_489), .B(n_460), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_502), .B(n_486), .C(n_504), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_510), .B(n_446), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_529), .B(n_444), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_509), .B(n_474), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_494), .B(n_460), .C(n_472), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_517), .A2(n_474), .B(n_336), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_520), .B(n_474), .Y(n_567) );
INVx3_ASAP7_75t_SL g568 ( .A(n_531), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
OAI31xp33_ASAP7_75t_SL g570 ( .A1(n_492), .A2(n_474), .A3(n_27), .B(n_28), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_505), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_511), .B(n_354), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_514), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_523), .B(n_25), .Y(n_575) );
AOI31xp33_ASAP7_75t_L g576 ( .A1(n_521), .A2(n_32), .A3(n_34), .B(n_35), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_522), .A2(n_328), .B1(n_336), .B2(n_343), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_503), .A2(n_317), .B(n_314), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_518), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_481), .Y(n_580) );
OA211x2_ASAP7_75t_L g581 ( .A1(n_526), .A2(n_41), .B(n_42), .C(n_44), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_519), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_524), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_493), .B(n_314), .C(n_274), .D(n_286), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_485), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_519), .B(n_354), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_47), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_488), .B(n_221), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_516), .B(n_50), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_485), .B(n_221), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_483), .B(n_51), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_488), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_495), .B(n_221), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_546), .B(n_496), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_551), .B(n_497), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_571), .B(n_497), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_495), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_568), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_537), .B(n_527), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_555), .B(n_221), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_539), .B(n_221), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_564), .B(n_209), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_593), .B(n_209), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_552), .B(n_209), .C(n_207), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_573), .B(n_209), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_534), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_541), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_560), .B(n_54), .Y(n_611) );
INVxp33_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_593), .B(n_209), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_582), .B(n_207), .Y(n_614) );
AND3x1_ASAP7_75t_L g615 ( .A(n_565), .B(n_56), .C(n_58), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_574), .B(n_207), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_557), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_536), .B(n_61), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_548), .Y(n_619) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_536), .B(n_354), .Y(n_620) );
NAND2x1_ASAP7_75t_L g621 ( .A(n_582), .B(n_354), .Y(n_621) );
AOI221x1_ASAP7_75t_L g622 ( .A1(n_565), .A2(n_540), .B1(n_591), .B2(n_575), .C(n_560), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_558), .Y(n_623) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_588), .A2(n_296), .B(n_309), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_569), .B(n_207), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_538), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_585), .B(n_207), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_540), .A2(n_343), .B1(n_320), .B2(n_194), .Y(n_630) );
INVx2_ASAP7_75t_R g631 ( .A(n_568), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_579), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_562), .B(n_194), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_570), .B(n_286), .C(n_308), .D(n_266), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_542), .B(n_343), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_561), .A2(n_343), .B1(n_320), .B2(n_194), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_582), .B(n_243), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_543), .B(n_243), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_553), .B(n_243), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_592), .B(n_63), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_544), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_533), .B(n_65), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_563), .B(n_242), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_548), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_563), .B(n_242), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_563), .B(n_242), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_541), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_559), .A2(n_320), .B1(n_243), .B2(n_242), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_554), .B(n_69), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_580), .B(n_70), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_627), .B(n_567), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_608), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_609), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_598), .B(n_579), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_612), .A2(n_559), .B1(n_549), .B2(n_550), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_612), .A2(n_584), .B(n_549), .C(n_587), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_598), .B(n_580), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_599), .B(n_594), .Y(n_658) );
XNOR2x2_ASAP7_75t_L g659 ( .A(n_641), .B(n_556), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_605), .A2(n_566), .B(n_576), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_625), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g662 ( .A(n_635), .B(n_589), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_632), .B(n_628), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_617), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_644), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_611), .A2(n_575), .B1(n_594), .B2(n_588), .C1(n_578), .C2(n_590), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_617), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_623), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_607), .B(n_577), .Y(n_670) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_619), .B(n_575), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_596), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_610), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_622), .A2(n_599), .B(n_648), .C(n_634), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_610), .Y(n_675) );
OA21x2_ASAP7_75t_SL g676 ( .A1(n_618), .A2(n_581), .B(n_572), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_595), .B(n_586), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_647), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_647), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_622), .B(n_72), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_615), .A2(n_286), .B(n_308), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_597), .B(n_76), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_620), .A2(n_308), .B(n_288), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_600), .A2(n_82), .B(n_266), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_626), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_602), .A2(n_272), .B(n_275), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_602), .A2(n_288), .B1(n_275), .B2(n_283), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_631), .B(n_288), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_603), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_631), .B(n_272), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_649), .B(n_288), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_640), .A2(n_283), .B(n_296), .C(n_298), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_649), .A2(n_288), .B1(n_298), .B2(n_306), .Y(n_693) );
XNOR2xp5_ASAP7_75t_L g694 ( .A(n_618), .B(n_306), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_630), .A2(n_309), .B1(n_642), .B2(n_636), .C(n_620), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_633), .Y(n_696) );
OAI21xp5_ASAP7_75t_SL g697 ( .A1(n_618), .A2(n_639), .B(n_638), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_601), .B(n_638), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_606), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_601), .B(n_639), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_624), .A2(n_604), .B(n_613), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_616), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_604), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_643), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_613), .Y(n_705) );
NOR3x1_ASAP7_75t_L g706 ( .A(n_621), .B(n_629), .C(n_633), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_643), .B(n_645), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_624), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_645), .A2(n_646), .B(n_650), .C(n_637), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_646), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_650), .Y(n_711) );
INVxp67_ASAP7_75t_L g712 ( .A(n_637), .Y(n_712) );
INVxp67_ASAP7_75t_L g713 ( .A(n_614), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_614), .B(n_621), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_608), .Y(n_715) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_674), .A2(n_697), .B(n_694), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_665), .A2(n_656), .B1(n_694), .B2(n_709), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_674), .A2(n_680), .B(n_655), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_676), .B(n_680), .C(n_666), .D(n_706), .Y(n_719) );
OA22x2_ASAP7_75t_L g720 ( .A1(n_659), .A2(n_654), .B1(n_701), .B2(n_663), .Y(n_720) );
INVxp67_ASAP7_75t_SL g721 ( .A(n_662), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_670), .A2(n_710), .B1(n_703), .B2(n_705), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_672), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_658), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_660), .A2(n_671), .B(n_670), .Y(n_725) );
OAI21xp33_ASAP7_75t_SL g726 ( .A1(n_660), .A2(n_714), .B(n_657), .Y(n_726) );
AO22x2_ASAP7_75t_SL g727 ( .A1(n_682), .A2(n_652), .B1(n_653), .B2(n_661), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g728 ( .A1(n_651), .A2(n_715), .B(n_684), .C(n_713), .Y(n_728) );
AO22x2_ASAP7_75t_L g729 ( .A1(n_664), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_729) );
XNOR2xp5_ASAP7_75t_L g730 ( .A(n_707), .B(n_704), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_718), .B(n_703), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_716), .A2(n_704), .B1(n_712), .B2(n_698), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_720), .A2(n_689), .B(n_691), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_721), .B(n_685), .Y(n_734) );
AOI211x1_ASAP7_75t_L g735 ( .A1(n_719), .A2(n_695), .B(n_700), .C(n_699), .Y(n_735) );
AND3x4_ASAP7_75t_L g736 ( .A(n_727), .B(n_673), .C(n_675), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_723), .Y(n_737) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_726), .A2(n_693), .B(n_702), .C(n_686), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_717), .A2(n_729), .B1(n_725), .B2(n_728), .C(n_722), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_738), .A2(n_730), .B(n_683), .Y(n_740) );
NAND5xp2_ASAP7_75t_L g741 ( .A(n_739), .B(n_691), .C(n_681), .D(n_683), .E(n_687), .Y(n_741) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_735), .B(n_724), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_732), .A2(n_729), .B1(n_711), .B2(n_696), .Y(n_743) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_736), .B(n_690), .C(n_692), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_742), .Y(n_745) );
OR4x2_ASAP7_75t_L g746 ( .A(n_741), .B(n_733), .C(n_731), .D(n_734), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_740), .B(n_737), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_747), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_745), .A2(n_743), .B1(n_744), .B2(n_708), .C(n_678), .Y(n_749) );
OAI222xp33_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_745), .B1(n_747), .B2(n_746), .C1(n_688), .C2(n_679), .Y(n_750) );
AO21x2_ASAP7_75t_L g751 ( .A1(n_749), .A2(n_746), .B(n_677), .Y(n_751) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_750), .A2(n_673), .B1(n_675), .B2(n_696), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_752), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_751), .B(n_745), .Y(n_754) );
endmodule