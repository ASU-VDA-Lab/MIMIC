module fake_netlist_6_2628_n_107 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_107);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_107;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_18;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVxp33_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVxp33_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_R g43 ( 
.A(n_18),
.B(n_2),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_29),
.C(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_45),
.B1(n_47),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_53),
.B1(n_23),
.B2(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_55),
.B1(n_34),
.B2(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_59),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_58),
.C(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_62),
.B1(n_59),
.B2(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_65),
.B(n_50),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_53),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_69),
.Y(n_77)
);

AO21x2_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_57),
.B(n_35),
.Y(n_78)
);

NAND2x1p5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_50),
.Y(n_79)
);

NAND4xp25_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_70),
.C(n_51),
.D(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_43),
.B1(n_34),
.B2(n_51),
.C(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_78),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_82),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_3),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_71),
.B(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_92),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_88),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_94),
.B(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_91),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_4),
.C(n_5),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);

OAI332xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_6),
.A3(n_8),
.B1(n_10),
.B2(n_14),
.B3(n_15),
.C1(n_53),
.C2(n_52),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_49),
.B(n_52),
.Y(n_107)
);


endmodule