module fake_jpeg_26486_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_58),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_30),
.B1(n_40),
.B2(n_39),
.Y(n_87)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_39),
.B1(n_27),
.B2(n_28),
.Y(n_95)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_45),
.B(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_72),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_40),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_64),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_84),
.B(n_67),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_43),
.B1(n_42),
.B2(n_35),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_87),
.B1(n_61),
.B2(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_41),
.B(n_45),
.C(n_36),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_94),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22x1_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_36),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_55),
.B1(n_38),
.B2(n_62),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_61),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_40),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_49),
.B1(n_54),
.B2(n_52),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_43),
.B1(n_42),
.B2(n_35),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_53),
.B1(n_38),
.B2(n_49),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_60),
.B(n_61),
.C(n_54),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_116),
.B1(n_76),
.B2(n_34),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_70),
.B(n_67),
.C(n_84),
.Y(n_107)
);

XOR2x1_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_23),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_47),
.C(n_65),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_38),
.C(n_33),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_120),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_49),
.B1(n_65),
.B2(n_63),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_52),
.B1(n_63),
.B2(n_56),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_33),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_93),
.B1(n_82),
.B2(n_71),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_128),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_133),
.Y(n_171)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_69),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_145),
.B1(n_117),
.B2(n_106),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_92),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_88),
.B1(n_69),
.B2(n_75),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_24),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_143),
.B(n_105),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_24),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_118),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_110),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_97),
.A2(n_90),
.B1(n_23),
.B2(n_12),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_8),
.Y(n_183)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_118),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_21),
.B1(n_20),
.B2(n_76),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_159),
.B(n_162),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_104),
.B(n_98),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_138),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_165),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_109),
.B(n_135),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_112),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_179),
.B1(n_183),
.B2(n_160),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_107),
.B(n_100),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_168),
.B(n_174),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_104),
.B(n_106),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_144),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_114),
.B1(n_117),
.B2(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_176),
.B1(n_185),
.B2(n_10),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_100),
.C(n_122),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_178),
.C(n_187),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_130),
.B(n_149),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_183),
.B(n_12),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_9),
.C(n_14),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_15),
.C(n_13),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_11),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_139),
.B1(n_132),
.B2(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_201),
.B1(n_187),
.B2(n_167),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_199),
.B(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_210),
.B(n_216),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_159),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_164),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_181),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_213),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_215),
.Y(n_235)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_218),
.B(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_202),
.B1(n_196),
.B2(n_210),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_198),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_197),
.B1(n_213),
.B2(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_238),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_191),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_207),
.B1(n_205),
.B2(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_238),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_165),
.C(n_161),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_234),
.C(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_162),
.C(n_159),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_181),
.C(n_160),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_195),
.C(n_196),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_233),
.C(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_251),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_250),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_257),
.B1(n_239),
.B2(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_226),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_190),
.B1(n_193),
.B2(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_232),
.A2(n_212),
.B(n_203),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_221),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_241),
.B(n_199),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_235),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_230),
.B1(n_227),
.B2(n_229),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_253),
.B1(n_271),
.B2(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_278),
.C(n_280),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_281),
.B(n_253),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_245),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_3),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_294),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_248),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_266),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_247),
.B(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_257),
.C(n_258),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.C(n_296),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_269),
.C(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_222),
.B1(n_236),
.B2(n_229),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_295),
.B1(n_277),
.B2(n_218),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_251),
.C(n_249),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_277),
.B1(n_268),
.B2(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_242),
.B1(n_201),
.B2(n_219),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_3),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_188),
.C(n_4),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_291),
.B(n_292),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_282),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_305),
.B(n_302),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_287),
.B(n_282),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_302),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_307),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_298),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_322),
.B(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_304),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_308),
.B(n_5),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_323),
.Y(n_326)
);

NAND4xp25_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_311),
.C(n_319),
.D(n_5),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_326),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_324),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_311),
.Y(n_331)
);


endmodule