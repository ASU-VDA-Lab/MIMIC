module fake_jpeg_1868_n_458 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_458);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_458;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_54),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_63),
.Y(n_119)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_56),
.Y(n_137)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_80),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_79),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_19),
.B(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_85),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_16),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_51),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_16),
.C(n_15),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_46),
.C(n_26),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_37),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_49),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_28),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_56),
.A2(n_38),
.B1(n_42),
.B2(n_51),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_132),
.B1(n_144),
.B2(n_163),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_54),
.A2(n_41),
.B(n_46),
.C(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_128),
.B(n_147),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_38),
.B1(n_42),
.B2(n_51),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_139),
.B(n_145),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_98),
.A2(n_38),
.B1(n_35),
.B2(n_47),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_35),
.B1(n_27),
.B2(n_33),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_35),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_150),
.B(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_48),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_87),
.B(n_20),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_159),
.B(n_166),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_58),
.A2(n_65),
.B1(n_113),
.B2(n_83),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_183),
.B1(n_106),
.B2(n_28),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_105),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_33),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_69),
.A2(n_44),
.B1(n_39),
.B2(n_36),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_167),
.A2(n_184),
.B1(n_144),
.B2(n_132),
.Y(n_230)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_73),
.B(n_27),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_186),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_97),
.A2(n_34),
.B1(n_20),
.B2(n_36),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_75),
.A2(n_34),
.B1(n_39),
.B2(n_44),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_81),
.A2(n_28),
.B1(n_24),
.B2(n_4),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_15),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_114),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_108),
.C(n_111),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_188),
.B(n_225),
.C(n_237),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_120),
.A2(n_100),
.B1(n_82),
.B2(n_107),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_189),
.A2(n_193),
.B1(n_224),
.B2(n_134),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_190),
.B(n_233),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_191),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_125),
.B(n_28),
.C(n_109),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_194),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_121),
.A2(n_2),
.B(n_3),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_200),
.B(n_213),
.Y(n_263)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_129),
.A2(n_28),
.B(n_15),
.C(n_13),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_202),
.A2(n_242),
.B(n_134),
.Y(n_275)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_28),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_109),
.B(n_78),
.C(n_4),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

OR2x4_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_78),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_205),
.A2(n_208),
.B(n_151),
.Y(n_259)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

OR2x4_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_2),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_2),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_210),
.B(n_220),
.Y(n_256)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_11),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_115),
.B(n_3),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_214),
.Y(n_274)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_5),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_184),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_222),
.A2(n_230),
.B1(n_231),
.B2(n_246),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_123),
.B(n_10),
.C(n_136),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_119),
.B(n_133),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_227),
.B(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_167),
.A2(n_163),
.B1(n_116),
.B2(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_126),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_165),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_235),
.B(n_248),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g236 ( 
.A1(n_155),
.A2(n_164),
.B1(n_171),
.B2(n_142),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_231),
.B1(n_200),
.B2(n_246),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_154),
.B(n_179),
.Y(n_237)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_117),
.Y(n_239)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_158),
.A2(n_154),
.B1(n_146),
.B2(n_179),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_243),
.B1(n_151),
.B2(n_160),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_180),
.A2(n_158),
.B(n_124),
.C(n_122),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_180),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_245),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_118),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_122),
.A2(n_130),
.B1(n_157),
.B2(n_140),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_130),
.B(n_157),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_279),
.B1(n_281),
.B2(n_288),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_259),
.A2(n_261),
.B(n_263),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_205),
.A2(n_160),
.B(n_173),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_173),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_292),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_275),
.A2(n_195),
.B1(n_207),
.B2(n_243),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_234),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_291),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_217),
.A2(n_193),
.B1(n_208),
.B2(n_199),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_280),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_217),
.A2(n_214),
.B1(n_203),
.B2(n_196),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_222),
.A2(n_202),
.B1(n_213),
.B2(n_242),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_215),
.B1(n_244),
.B2(n_218),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_214),
.A2(n_229),
.B1(n_224),
.B2(n_213),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_200),
.A2(n_191),
.B1(n_204),
.B2(n_237),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_264),
.B1(n_258),
.B2(n_267),
.Y(n_324)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_238),
.A2(n_194),
.A3(n_236),
.B1(n_206),
.B2(n_211),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_188),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_262),
.B1(n_289),
.B2(n_266),
.Y(n_351)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_272),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_298),
.B(n_308),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_212),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_302),
.C(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_303),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_237),
.C(n_236),
.Y(n_302)
);

XNOR2x2_ASAP7_75t_SL g303 ( 
.A(n_250),
.B(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_198),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_256),
.B(n_201),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_310),
.B(n_316),
.Y(n_349)
);

INVx4_ASAP7_75t_SL g312 ( 
.A(n_273),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_312),
.A2(n_321),
.B1(n_324),
.B2(n_262),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_223),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_315),
.Y(n_342)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_256),
.B(n_219),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_320),
.B(n_285),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_239),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_289),
.C(n_265),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_259),
.A2(n_223),
.B(n_197),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_254),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_258),
.B(n_276),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_328),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_337),
.C(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_304),
.B(n_288),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_341),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_322),
.A2(n_269),
.B1(n_284),
.B2(n_264),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_351),
.B1(n_353),
.B2(n_356),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_282),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_261),
.B(n_282),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_339),
.A2(n_350),
.B(n_296),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_282),
.C(n_269),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_319),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_314),
.B1(n_325),
.B2(n_323),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_355),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_320),
.A2(n_271),
.B(n_267),
.Y(n_350)
);

OAI32xp33_ASAP7_75t_L g352 ( 
.A1(n_294),
.A2(n_280),
.A3(n_266),
.B1(n_265),
.B2(n_287),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_307),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_280),
.B1(n_253),
.B2(n_273),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_253),
.C(n_277),
.Y(n_355)
);

AO32x1_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_303),
.A3(n_318),
.B1(n_301),
.B2(n_317),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_339),
.A2(n_332),
.B1(n_353),
.B2(n_345),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_370),
.B1(n_371),
.B2(n_373),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_365),
.Y(n_385)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_347),
.A2(n_303),
.A3(n_310),
.B1(n_305),
.B2(n_300),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_367),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_365),
.B(n_379),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_346),
.A2(n_314),
.B1(n_312),
.B2(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_340),
.Y(n_367)
);

AO32x1_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_306),
.A3(n_297),
.B1(n_277),
.B2(n_278),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_369),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_312),
.B1(n_316),
.B2(n_326),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_372),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_295),
.B1(n_321),
.B2(n_273),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_376),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_342),
.B(n_278),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_377),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_251),
.B1(n_347),
.B2(n_355),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_378),
.A2(n_350),
.B1(n_342),
.B2(n_349),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g379 ( 
.A(n_341),
.B(n_251),
.CI(n_333),
.CON(n_379),
.SN(n_379)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_385),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_335),
.C(n_331),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_395),
.C(n_357),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_335),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_392),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_352),
.B1(n_351),
.B2(n_348),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_390),
.A2(n_378),
.B1(n_377),
.B2(n_361),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_341),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_337),
.C(n_343),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_370),
.A2(n_343),
.B1(n_354),
.B2(n_338),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_396),
.A2(n_360),
.B1(n_369),
.B2(n_354),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_404),
.Y(n_420)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_388),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_405),
.Y(n_415)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_380),
.B(n_367),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_329),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_406),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_412),
.Y(n_419)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_393),
.Y(n_408)
);

INVx13_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_409),
.A2(n_410),
.B1(n_411),
.B2(n_413),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_384),
.A2(n_375),
.B1(n_358),
.B2(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_391),
.Y(n_411)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_390),
.B1(n_394),
.B2(n_384),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_424),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_399),
.A2(n_398),
.B(n_385),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_412),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_399),
.A2(n_382),
.B(n_363),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_397),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_402),
.A2(n_413),
.B1(n_411),
.B2(n_382),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_391),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_427),
.B(n_392),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_431),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_SL g427 ( 
.A(n_419),
.B(n_407),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_428),
.A2(n_415),
.B1(n_420),
.B2(n_403),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_414),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_372),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_386),
.C(n_383),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_400),
.Y(n_437)
);

BUFx24_ASAP7_75t_SL g433 ( 
.A(n_418),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_387),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_425),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_440),
.B1(n_441),
.B2(n_415),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_439),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_438),
.C(n_389),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_400),
.C(n_416),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_443),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_435),
.A2(n_421),
.B(n_414),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_446),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_440),
.A2(n_420),
.B(n_364),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_424),
.C(n_381),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_381),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_449),
.B(n_451),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_450),
.B(n_439),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_453),
.B(n_448),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_452),
.C(n_408),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_404),
.C(n_369),
.Y(n_456)
);

OAI221xp5_ASAP7_75t_L g457 ( 
.A1(n_456),
.A2(n_422),
.B1(n_379),
.B2(n_389),
.C(n_338),
.Y(n_457)
);

OAI321xp33_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_251),
.A3(n_357),
.B1(n_379),
.B2(n_422),
.C(n_398),
.Y(n_458)
);


endmodule