module fake_netlist_1_3777_n_33 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_5), .B(n_2), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_12), .B(n_5), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_10), .B(n_7), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_1), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx4_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AO32x2_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_16), .A3(n_14), .B1(n_15), .B2(n_18), .Y(n_21) );
AOI221xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_13), .B1(n_17), .B2(n_15), .C(n_3), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_0), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
OAI21xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .B(n_17), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_0), .Y(n_26) );
XOR2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_1), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_2), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_30), .B(n_29), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_25), .B1(n_15), .B2(n_19), .Y(n_32) );
OAI221xp5_ASAP7_75t_R g33 ( .A1(n_32), .A2(n_4), .B1(n_6), .B2(n_9), .C(n_11), .Y(n_33) );
endmodule