module fake_jpeg_14663_n_25 (n_3, n_2, n_1, n_0, n_4, n_5, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_5),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_L g8 ( 
.A1(n_1),
.A2(n_5),
.B1(n_4),
.B2(n_3),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_SL g9 ( 
.A1(n_2),
.A2(n_4),
.B1(n_0),
.B2(n_3),
.Y(n_9)
);

INVx6_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_SL g11 ( 
.A1(n_4),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

AO21x1_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_2),
.B(n_0),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_16),
.B1(n_10),
.B2(n_7),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_6),
.A2(n_1),
.B(n_8),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_9),
.B(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_11),
.B1(n_8),
.B2(n_7),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_8),
.B1(n_11),
.B2(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_9),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_14),
.B2(n_7),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_22),
.B1(n_10),
.B2(n_20),
.Y(n_24)
);

AO221x1_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_10),
.B1(n_13),
.B2(n_7),
.C(n_16),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_21),
.C(n_23),
.Y(n_25)
);


endmodule