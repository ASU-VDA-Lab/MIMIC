module real_aes_2374_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_794, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_794;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g207 ( .A(n_0), .B(n_129), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_1), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_2), .B(n_135), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_3), .B(n_125), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_4), .B(n_135), .Y(n_148) );
INVx1_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
NAND2xp33_ASAP7_75t_SL g199 ( .A(n_6), .B(n_133), .Y(n_199) );
INVx1_ASAP7_75t_L g180 ( .A(n_7), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_8), .A2(n_42), .B1(n_103), .B2(n_104), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_8), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g762 ( .A(n_9), .Y(n_762) );
AND2x2_ASAP7_75t_L g146 ( .A(n_10), .B(n_139), .Y(n_146) );
AND2x2_ASAP7_75t_L g491 ( .A(n_11), .B(n_173), .Y(n_491) );
AND2x2_ASAP7_75t_L g499 ( .A(n_12), .B(n_196), .Y(n_499) );
INVx2_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_14), .B(n_125), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_15), .Y(n_434) );
AOI221x1_ASAP7_75t_L g193 ( .A1(n_16), .A2(n_117), .B1(n_194), .B2(n_196), .C(n_198), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_17), .B(n_135), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_18), .B(n_135), .Y(n_472) );
INVx1_ASAP7_75t_L g437 ( .A(n_19), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_20), .A2(n_89), .B1(n_135), .B2(n_181), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_21), .A2(n_117), .B(n_150), .Y(n_149) );
AOI221xp5_ASAP7_75t_SL g160 ( .A1(n_22), .A2(n_37), .B1(n_117), .B2(n_135), .C(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_23), .B(n_129), .Y(n_151) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_24), .A2(n_101), .B1(n_755), .B2(n_766), .C1(n_782), .C2(n_786), .Y(n_100) );
AOI22xp5_ASAP7_75t_SL g773 ( .A1(n_24), .A2(n_77), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_24), .Y(n_775) );
OR2x2_ASAP7_75t_L g141 ( .A(n_25), .B(n_88), .Y(n_141) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_25), .A2(n_88), .B(n_140), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_26), .B(n_125), .Y(n_172) );
INVxp67_ASAP7_75t_L g192 ( .A(n_27), .Y(n_192) );
AND2x2_ASAP7_75t_L g223 ( .A(n_28), .B(n_138), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_29), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_30), .A2(n_117), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_31), .A2(n_196), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_32), .B(n_125), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_33), .A2(n_117), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_34), .B(n_125), .Y(n_458) );
AND2x2_ASAP7_75t_L g118 ( .A(n_35), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g133 ( .A(n_35), .B(n_122), .Y(n_133) );
INVx1_ASAP7_75t_L g188 ( .A(n_35), .Y(n_188) );
OR2x6_ASAP7_75t_L g435 ( .A(n_36), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_38), .B(n_135), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_39), .A2(n_81), .B1(n_117), .B2(n_186), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_40), .B(n_125), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_41), .B(n_135), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_42), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_43), .B(n_129), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_44), .A2(n_117), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g210 ( .A(n_45), .B(n_138), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_46), .B(n_129), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_47), .B(n_138), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_48), .B(n_135), .Y(n_447) );
INVx1_ASAP7_75t_L g121 ( .A(n_49), .Y(n_121) );
INVx1_ASAP7_75t_L g131 ( .A(n_49), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_50), .B(n_125), .Y(n_497) );
AND2x2_ASAP7_75t_L g463 ( .A(n_51), .B(n_138), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_52), .B(n_135), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_53), .B(n_129), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_54), .B(n_129), .Y(n_457) );
AND2x2_ASAP7_75t_L g142 ( .A(n_55), .B(n_138), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_56), .B(n_135), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_57), .B(n_125), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_58), .B(n_135), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_59), .A2(n_117), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_60), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_61), .B(n_139), .Y(n_175) );
AND2x2_ASAP7_75t_L g478 ( .A(n_62), .B(n_139), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_63), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_64), .A2(n_117), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_65), .B(n_125), .Y(n_152) );
AND2x2_ASAP7_75t_SL g260 ( .A(n_66), .B(n_173), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_67), .B(n_129), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_68), .B(n_129), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_69), .A2(n_92), .B1(n_117), .B2(n_186), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_70), .B(n_125), .Y(n_475) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
INVx1_ASAP7_75t_L g127 ( .A(n_71), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_72), .B(n_129), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_73), .A2(n_117), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_74), .A2(n_117), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_75), .A2(n_117), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g460 ( .A(n_76), .B(n_139), .Y(n_460) );
INVx1_ASAP7_75t_L g774 ( .A(n_77), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_78), .B(n_138), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_79), .B(n_135), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_80), .A2(n_83), .B1(n_135), .B2(n_181), .Y(n_258) );
INVx1_ASAP7_75t_L g438 ( .A(n_82), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_84), .B(n_129), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_85), .B(n_129), .Y(n_163) );
AND2x2_ASAP7_75t_L g529 ( .A(n_86), .B(n_173), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_87), .A2(n_117), .B(n_123), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_90), .B(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_91), .A2(n_117), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_93), .B(n_125), .Y(n_527) );
INVxp67_ASAP7_75t_L g195 ( .A(n_94), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_95), .B(n_135), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_96), .B(n_125), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_97), .A2(n_117), .B(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g477 ( .A(n_98), .Y(n_477) );
BUFx2_ASAP7_75t_L g763 ( .A(n_99), .Y(n_763) );
BUFx2_ASAP7_75t_SL g790 ( .A(n_99), .Y(n_790) );
AO221x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_105), .B1(n_741), .B2(n_749), .C(n_750), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_102), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_432), .B1(n_439), .B2(n_739), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_106), .B(n_747), .Y(n_746) );
AOI22x1_ASAP7_75t_L g770 ( .A1(n_106), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
INVx4_ASAP7_75t_L g771 ( .A(n_106), .Y(n_771) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_371), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_264), .C(n_315), .Y(n_107) );
OAI211xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_154), .B(n_211), .C(n_242), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_143), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_113), .B(n_216), .Y(n_379) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g224 ( .A(n_114), .B(n_145), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_114), .B(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g241 ( .A(n_114), .B(n_231), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_114), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g278 ( .A(n_114), .B(n_254), .Y(n_278) );
INVx2_ASAP7_75t_L g304 ( .A(n_114), .Y(n_304) );
AND2x4_ASAP7_75t_L g313 ( .A(n_114), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g418 ( .A(n_114), .B(n_285), .Y(n_418) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_137), .B(n_142), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_134), .Y(n_115) );
AND2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
BUFx3_ASAP7_75t_L g185 ( .A(n_118), .Y(n_185) );
AND2x6_ASAP7_75t_L g129 ( .A(n_119), .B(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g190 ( .A(n_119), .Y(n_190) );
AND2x4_ASAP7_75t_L g186 ( .A(n_120), .B(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g125 ( .A(n_121), .B(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g183 ( .A(n_121), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_122), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_128), .B(n_132), .Y(n_123) );
AND2x4_ASAP7_75t_L g136 ( .A(n_126), .B(n_130), .Y(n_136) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_129), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_132), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_132), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_132), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_132), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_132), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_132), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_132), .A2(n_457), .B(n_458), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_132), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_132), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_132), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_132), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_132), .A2(n_527), .B(n_528), .Y(n_526) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g135 ( .A(n_133), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_137), .A2(n_217), .B(n_223), .Y(n_216) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_137), .A2(n_217), .B(n_223), .Y(n_231) );
AOI21x1_ASAP7_75t_L g484 ( .A1(n_137), .A2(n_485), .B(n_491), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_138), .Y(n_137) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_138), .A2(n_160), .B(n_164), .Y(n_159) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_138), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_138), .A2(n_524), .B(n_525), .Y(n_523) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g153 ( .A(n_140), .B(n_141), .Y(n_153) );
AND2x2_ASAP7_75t_L g302 ( .A(n_143), .B(n_303), .Y(n_302) );
OAI32xp33_ASAP7_75t_L g385 ( .A1(n_143), .A2(n_307), .A3(n_311), .B1(n_318), .B2(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_143), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g239 ( .A(n_144), .B(n_240), .Y(n_239) );
NAND3xp33_ASAP7_75t_L g312 ( .A(n_144), .B(n_234), .C(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g338 ( .A(n_144), .B(n_241), .Y(n_338) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_145), .Y(n_228) );
INVx5_ASAP7_75t_L g263 ( .A(n_145), .Y(n_263) );
AND2x4_ASAP7_75t_L g319 ( .A(n_145), .B(n_231), .Y(n_319) );
OR2x2_ASAP7_75t_L g334 ( .A(n_145), .B(n_254), .Y(n_334) );
OR2x2_ASAP7_75t_L g360 ( .A(n_145), .B(n_216), .Y(n_360) );
AND2x2_ASAP7_75t_L g368 ( .A(n_145), .B(n_314), .Y(n_368) );
AND2x4_ASAP7_75t_SL g393 ( .A(n_145), .B(n_313), .Y(n_393) );
OR2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_153), .B(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_153), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_153), .B(n_195), .Y(n_194) );
NOR3xp33_ASAP7_75t_L g198 ( .A(n_153), .B(n_199), .C(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_153), .A2(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_153), .A2(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_155), .B(n_313), .Y(n_389) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_165), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_156), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OR2x6_ASAP7_75t_SL g213 ( .A(n_157), .B(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_158), .B(n_273), .Y(n_291) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_158), .Y(n_429) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g246 ( .A(n_159), .Y(n_246) );
AND2x2_ASAP7_75t_L g271 ( .A(n_159), .B(n_202), .Y(n_271) );
INVx2_ASAP7_75t_L g299 ( .A(n_159), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_159), .B(n_166), .Y(n_340) );
BUFx3_ASAP7_75t_L g364 ( .A(n_159), .Y(n_364) );
OR2x2_ASAP7_75t_L g376 ( .A(n_159), .B(n_166), .Y(n_376) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_159), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_165), .A2(n_407), .B1(n_410), .B2(n_411), .Y(n_406) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_176), .Y(n_165) );
INVx1_ASAP7_75t_L g234 ( .A(n_166), .Y(n_234) );
OR2x2_ASAP7_75t_L g245 ( .A(n_166), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g252 ( .A(n_166), .Y(n_252) );
AND2x4_ASAP7_75t_SL g269 ( .A(n_166), .B(n_177), .Y(n_269) );
AND2x4_ASAP7_75t_L g274 ( .A(n_166), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g283 ( .A(n_166), .Y(n_283) );
OR2x2_ASAP7_75t_L g289 ( .A(n_166), .B(n_177), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_166), .B(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_166), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_166), .B(n_271), .Y(n_405) );
OR2x2_ASAP7_75t_L g421 ( .A(n_166), .B(n_324), .Y(n_421) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_175), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
INVx2_ASAP7_75t_SL g256 ( .A(n_173), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_173), .A2(n_472), .B(n_473), .Y(n_471) );
BUFx4f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx3_ASAP7_75t_L g197 ( .A(n_174), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_176), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g247 ( .A(n_176), .Y(n_247) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_176), .B(n_238), .Y(n_354) );
AND2x4_ASAP7_75t_L g176 ( .A(n_177), .B(n_201), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_177), .B(n_202), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_177), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_177), .B(n_246), .Y(n_250) );
INVx3_ASAP7_75t_L g275 ( .A(n_177), .Y(n_275) );
INVx1_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
AND2x2_ASAP7_75t_L g388 ( .A(n_177), .B(n_252), .Y(n_388) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B1(n_186), .B2(n_191), .Y(n_178) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_185), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g453 ( .A(n_196), .Y(n_453) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21x1_ASAP7_75t_L g203 ( .A1(n_197), .A2(n_204), .B(n_210), .Y(n_203) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_197), .A2(n_493), .B(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_202), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
AND2x2_ASAP7_75t_L g298 ( .A(n_202), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g324 ( .A(n_202), .B(n_246), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_202), .B(n_275), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_202), .Y(n_347) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AOI222xp33_ASAP7_75t_SL g211 ( .A1(n_212), .A2(n_215), .B1(n_225), .B2(n_232), .C1(n_235), .C2(n_239), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_224), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_216), .B(n_285), .Y(n_336) );
AND2x4_ASAP7_75t_L g352 ( .A(n_216), .B(n_263), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_222), .Y(n_217) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_227), .B(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g277 ( .A(n_228), .B(n_278), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g242 ( .A1(n_229), .A2(n_243), .B1(n_248), .B2(n_253), .C1(n_261), .C2(n_794), .Y(n_242) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g381 ( .A(n_230), .B(n_285), .Y(n_381) );
OR2x2_ASAP7_75t_L g424 ( .A(n_230), .B(n_330), .Y(n_424) );
AND2x2_ASAP7_75t_L g253 ( .A(n_231), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g314 ( .A(n_231), .Y(n_314) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_231), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_232), .A2(n_343), .B(n_348), .C(n_349), .Y(n_342) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g370 ( .A(n_234), .Y(n_370) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g300 ( .A(n_239), .Y(n_300) );
AND2x2_ASAP7_75t_L g284 ( .A(n_240), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_240), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OAI31xp33_ASAP7_75t_L g335 ( .A1(n_243), .A2(n_261), .A3(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_244), .A2(n_294), .B(n_338), .C(n_339), .Y(n_337) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
OR2x2_ASAP7_75t_L g326 ( .A(n_245), .B(n_275), .Y(n_326) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
BUFx2_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
AND2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
AOI21x1_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_260), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_263), .B(n_320), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_276), .B(n_279), .C(n_301), .Y(n_264) );
INVxp33_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_272), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g305 ( .A(n_269), .B(n_298), .Y(n_305) );
OR2x2_ASAP7_75t_L g281 ( .A(n_270), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g311 ( .A(n_270), .B(n_285), .Y(n_311) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g387 ( .A(n_271), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g410 ( .A(n_272), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_274), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_274), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g422 ( .A(n_274), .B(n_298), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_274), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g365 ( .A(n_275), .B(n_347), .Y(n_365) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AOI322xp5_ASAP7_75t_L g419 ( .A1(n_278), .A2(n_298), .A3(n_352), .B1(n_377), .B2(n_420), .C1(n_422), .C2(n_423), .Y(n_419) );
AOI211xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_284), .B(n_286), .C(n_295), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_282), .B(n_310), .Y(n_332) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_298), .Y(n_297) );
NOR2x1p5_ASAP7_75t_L g363 ( .A(n_283), .B(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_283), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_284), .A2(n_302), .B(n_305), .C(n_306), .Y(n_301) );
AND2x4_ASAP7_75t_L g320 ( .A(n_285), .B(n_304), .Y(n_320) );
INVx2_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_285), .B(n_319), .Y(n_350) );
AND2x2_ASAP7_75t_L g392 ( .A(n_285), .B(n_393), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_285), .B(n_409), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_285), .B(n_313), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B(n_292), .Y(n_286) );
AND2x2_ASAP7_75t_L g382 ( .A(n_288), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_303), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g397 ( .A(n_303), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_309), .B(n_311), .C(n_312), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_310), .Y(n_394) );
INVx3_ASAP7_75t_SL g409 ( .A(n_313), .Y(n_409) );
NAND5xp2_ASAP7_75t_L g315 ( .A(n_316), .B(n_335), .C(n_342), .D(n_355), .E(n_366), .Y(n_315) );
AOI222xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_325), .B2(n_327), .C1(n_331), .C2(n_333), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_318), .A2(n_399), .B1(n_403), .B2(n_404), .Y(n_398) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g348 ( .A(n_319), .B(n_320), .Y(n_348) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_329), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_330), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g367 ( .A(n_330), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g378 ( .A(n_330), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g408 ( .A(n_334), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g356 ( .A(n_341), .Y(n_356) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B(n_353), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_352), .A2(n_356), .B1(n_357), .B2(n_361), .Y(n_355) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_352), .Y(n_403) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g369 ( .A(n_354), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g374 ( .A(n_356), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_SL g402 ( .A(n_365), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_390), .C(n_413), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_389), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_380), .B2(n_382), .C(n_385), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g414 ( .A(n_376), .B(n_402), .Y(n_414) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OAI321xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .A3(n_395), .B1(n_397), .B2(n_398), .C(n_406), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_404), .A2(n_426), .B1(n_430), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B(n_419), .C(n_425), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_433), .Y(n_748) );
AND2x6_ASAP7_75t_SL g433 ( .A(n_434), .B(n_435), .Y(n_433) );
OR2x6_ASAP7_75t_SL g739 ( .A(n_434), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g754 ( .A(n_434), .B(n_435), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_434), .B(n_740), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_435), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx4_ASAP7_75t_L g745 ( .A(n_439), .Y(n_745) );
AND3x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_617), .C(n_713), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_559), .C(n_586), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_479), .B(n_508), .C(n_532), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_461), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_443), .A2(n_510), .B(n_514), .C(n_520), .Y(n_509) );
OR2x2_ASAP7_75t_L g632 ( .A(n_443), .B(n_569), .Y(n_632) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g599 ( .A(n_444), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_444), .B(n_570), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_444), .B(n_715), .Y(n_730) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
AND2x2_ASAP7_75t_L g516 ( .A(n_445), .B(n_462), .Y(n_516) );
INVx1_ASAP7_75t_L g536 ( .A(n_445), .Y(n_536) );
OR2x2_ASAP7_75t_L g551 ( .A(n_445), .B(n_470), .Y(n_551) );
INVx2_ASAP7_75t_L g557 ( .A(n_445), .Y(n_557) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_445), .Y(n_612) );
INVx1_ASAP7_75t_L g689 ( .A(n_445), .Y(n_689) );
NOR2x1_ASAP7_75t_SL g538 ( .A(n_452), .B(n_470), .Y(n_538) );
AND2x2_ASAP7_75t_L g568 ( .A(n_452), .B(n_557), .Y(n_568) );
AO21x1_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B(n_460), .Y(n_452) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_453), .A2(n_454), .B(n_460), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
OR2x2_ASAP7_75t_L g562 ( .A(n_461), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_461), .B(n_669), .Y(n_668) );
INVx3_ASAP7_75t_L g690 ( .A(n_461), .Y(n_690) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_470), .Y(n_461) );
OR2x2_ASAP7_75t_SL g550 ( .A(n_462), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g554 ( .A(n_462), .Y(n_554) );
INVx4_ASAP7_75t_L g570 ( .A(n_462), .Y(n_570) );
OR2x2_ASAP7_75t_L g585 ( .A(n_462), .B(n_518), .Y(n_585) );
AND2x2_ASAP7_75t_L g624 ( .A(n_462), .B(n_538), .Y(n_624) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_462), .Y(n_636) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AND2x2_ASAP7_75t_L g517 ( .A(n_470), .B(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g569 ( .A(n_470), .B(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g584 ( .A(n_470), .Y(n_584) );
AND2x2_ASAP7_75t_L g600 ( .A(n_470), .B(n_570), .Y(n_600) );
AND2x2_ASAP7_75t_L g613 ( .A(n_470), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g645 ( .A(n_470), .B(n_557), .Y(n_645) );
INVx2_ASAP7_75t_SL g715 ( .A(n_470), .Y(n_715) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_478), .Y(n_470) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp67_ASAP7_75t_L g480 ( .A(n_481), .B(n_500), .Y(n_480) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_481), .A2(n_587), .B(n_591), .C(n_607), .Y(n_586) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g682 ( .A(n_482), .B(n_521), .Y(n_682) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx2_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_483), .B(n_522), .Y(n_542) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_483), .Y(n_546) );
AND2x2_ASAP7_75t_L g604 ( .A(n_483), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g678 ( .A(n_483), .Y(n_678) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_484), .Y(n_580) );
AND2x2_ASAP7_75t_L g623 ( .A(n_484), .B(n_492), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_490), .Y(n_485) );
INVx2_ASAP7_75t_L g513 ( .A(n_492), .Y(n_513) );
AND2x2_ASAP7_75t_L g573 ( .A(n_492), .B(n_522), .Y(n_573) );
INVx2_ASAP7_75t_L g605 ( .A(n_492), .Y(n_605) );
OR2x2_ASAP7_75t_L g628 ( .A(n_492), .B(n_503), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_500), .B(n_545), .Y(n_652) );
AND2x2_ASAP7_75t_L g686 ( .A(n_500), .B(n_622), .Y(n_686) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI31xp33_ASAP7_75t_SL g607 ( .A1(n_501), .A2(n_588), .A3(n_608), .B(n_615), .Y(n_607) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_502), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g541 ( .A(n_503), .Y(n_541) );
AND2x2_ASAP7_75t_L g558 ( .A(n_503), .B(n_521), .Y(n_558) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g548 ( .A(n_504), .B(n_505), .Y(n_548) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g693 ( .A(n_511), .Y(n_693) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_513), .B(n_522), .Y(n_575) );
AND2x2_ASAP7_75t_L g616 ( .A(n_513), .B(n_531), .Y(n_616) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_554), .Y(n_596) );
AND2x2_ASAP7_75t_L g555 ( .A(n_518), .B(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_518), .Y(n_564) );
INVx2_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
AND2x2_ASAP7_75t_L g704 ( .A(n_518), .B(n_689), .Y(n_704) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g710 ( .A(n_520), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_521), .B(n_580), .Y(n_649) );
AND2x2_ASAP7_75t_L g697 ( .A(n_521), .B(n_623), .Y(n_697) );
INVx4_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g606 ( .A(n_522), .B(n_578), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_522), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g627 ( .A(n_522), .Y(n_627) );
BUFx2_ASAP7_75t_L g643 ( .A(n_522), .Y(n_643) );
AND2x4_ASAP7_75t_L g677 ( .A(n_522), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g722 ( .A(n_522), .B(n_623), .Y(n_722) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .Y(n_522) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_539), .B1(n_543), .B2(n_549), .C1(n_552), .C2(n_558), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_534), .A2(n_598), .B1(n_601), .B2(n_606), .Y(n_597) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
AND2x2_ASAP7_75t_L g581 ( .A(n_535), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_535), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_535), .B(n_600), .Y(n_733) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g694 ( .A(n_536), .B(n_600), .Y(n_694) );
OR2x2_ASAP7_75t_L g671 ( .A(n_537), .B(n_553), .Y(n_671) );
OR2x2_ASAP7_75t_L g679 ( .A(n_537), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g663 ( .A(n_538), .B(n_556), .Y(n_663) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g571 ( .A(n_541), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g721 ( .A(n_541), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g672 ( .A(n_542), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_542), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g707 ( .A(n_542), .Y(n_707) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
INVx2_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g594 ( .A(n_546), .B(n_573), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_547), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g593 ( .A(n_547), .Y(n_593) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_547), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g696 ( .A(n_547), .B(n_568), .Y(n_696) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g630 ( .A(n_548), .B(n_616), .Y(n_630) );
AND2x2_ASAP7_75t_L g673 ( .A(n_548), .B(n_605), .Y(n_673) );
AND2x4_ASAP7_75t_L g588 ( .A(n_549), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g729 ( .A(n_551), .B(n_585), .Y(n_729) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_553), .B(n_568), .Y(n_712) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_554), .B(n_568), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_554), .A2(n_595), .B(n_696), .C(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g726 ( .A(n_554), .B(n_704), .Y(n_726) );
INVx1_ASAP7_75t_L g637 ( .A(n_555), .Y(n_637) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_558), .B(n_622), .Y(n_621) );
OAI21xp33_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_571), .B(n_574), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_565), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_562), .A2(n_715), .B1(n_716), .B2(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g590 ( .A(n_564), .Y(n_590) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_570), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g662 ( .A(n_570), .Y(n_662) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_581), .Y(n_574) );
INVx1_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_595), .B(n_597), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g638 ( .A(n_593), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g675 ( .A(n_593), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_593), .B(n_623), .Y(n_711) );
INVx1_ASAP7_75t_L g731 ( .A(n_594), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_596), .A2(n_699), .B1(n_702), .B2(n_705), .C(n_708), .Y(n_698) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI321xp33_ASAP7_75t_L g719 ( .A1(n_601), .A2(n_636), .A3(n_720), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g660 ( .A(n_605), .Y(n_660) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g654 ( .A(n_610), .Y(n_654) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g680 ( .A(n_611), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_613), .A2(n_641), .B1(n_645), .B2(n_646), .C(n_651), .Y(n_640) );
INVxp67_ASAP7_75t_L g669 ( .A(n_614), .Y(n_669) );
INVx1_ASAP7_75t_L g639 ( .A(n_616), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_618), .B(n_664), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_640), .C(n_655), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_624), .B1(n_625), .B2(n_631), .C(n_633), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g738 ( .A(n_623), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_629), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_627), .B(n_673), .Y(n_718) );
INVx2_ASAP7_75t_SL g650 ( .A(n_628), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_629), .A2(n_634), .B1(n_635), .B2(n_638), .Y(n_633) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_637), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_638), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g644 ( .A(n_639), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_641), .A2(n_684), .B1(n_686), .B2(n_687), .C1(n_691), .C2(n_694), .Y(n_683) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_642), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g717 ( .A(n_642), .B(n_696), .Y(n_717) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_650), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_650), .B(n_710), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_654), .Y(n_651) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_661), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND4xp25_ASAP7_75t_SL g664 ( .A(n_665), .B(n_683), .C(n_695), .D(n_698), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B(n_672), .C(n_674), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_671), .A2(n_675), .B1(n_679), .B2(n_681), .Y(n_674) );
INVx1_ASAP7_75t_L g701 ( .A(n_673), .Y(n_701) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_690), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_707), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_712), .Y(n_708) );
NOR4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_719), .C(n_732), .D(n_734), .Y(n_713) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx11_ASAP7_75t_R g744 ( .A(n_739), .Y(n_744) );
OAI21x1_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_745), .B(n_746), .Y(n_741) );
BUFx4f_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_764), .Y(n_757) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_760), .B(n_763), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_SL g785 ( .A(n_761), .B(n_763), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_761), .A2(n_788), .B(n_791), .Y(n_787) );
INVx1_ASAP7_75t_SL g769 ( .A(n_764), .Y(n_769) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx3_ASAP7_75t_L g780 ( .A(n_765), .Y(n_780) );
BUFx2_ASAP7_75t_L g792 ( .A(n_765), .Y(n_792) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AOI21xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_770), .B(n_776), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVxp33_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_SL g776 ( .A(n_777), .B(n_781), .Y(n_776) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
CKINVDCx9p33_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
endmodule