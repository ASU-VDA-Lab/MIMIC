module fake_jpeg_12091_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_378;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_54),
.Y(n_114)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_9),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_74),
.Y(n_126)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g119 ( 
.A(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_79),
.Y(n_156)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_82),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_88),
.B(n_92),
.Y(n_145)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_29),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

BUFx2_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_47),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_12),
.Y(n_152)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_32),
.C(n_34),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_105),
.B(n_46),
.C(n_45),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_39),
.B1(n_22),
.B2(n_44),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_110),
.A2(n_123),
.B1(n_136),
.B2(n_39),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_44),
.B1(n_46),
.B2(n_45),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_65),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_132),
.Y(n_175)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_142),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_79),
.A2(n_39),
.B1(n_22),
.B2(n_27),
.Y(n_136)
);

CKINVDCx12_ASAP7_75t_R g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_51),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_101),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_77),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_163),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_62),
.B1(n_61),
.B2(n_72),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_166),
.A2(n_87),
.B1(n_84),
.B2(n_112),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_167),
.B(n_173),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_186),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_43),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_20),
.B(n_1),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_178),
.A2(n_196),
.B(n_198),
.Y(n_246)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_43),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_182),
.B(n_184),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_187),
.B1(n_81),
.B2(n_85),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_33),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_33),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_136),
.A2(n_94),
.B1(n_93),
.B2(n_83),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_135),
.B(n_40),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_188),
.B(n_202),
.Y(n_212)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_22),
.B1(n_80),
.B2(n_75),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_40),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_121),
.B(n_0),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_110),
.A2(n_20),
.B(n_89),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

NAND2x1p5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_20),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_11),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_120),
.Y(n_203)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_113),
.B(n_86),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_89),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_196),
.B(n_163),
.C(n_206),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_226),
.B1(n_106),
.B2(n_125),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_175),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_223),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_229),
.B1(n_199),
.B2(n_200),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_111),
.B1(n_112),
.B2(n_129),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_118),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_116),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_155),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_178),
.B1(n_210),
.B2(n_198),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_255),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_172),
.B(n_164),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_252),
.A2(n_261),
.B(n_272),
.Y(n_318)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_269),
.B1(n_275),
.B2(n_222),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_171),
.B(n_150),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_267),
.Y(n_291)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_185),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_192),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_120),
.B1(n_129),
.B2(n_157),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_214),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_273),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_176),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_274),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_106),
.B1(n_154),
.B2(n_141),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_218),
.B(n_148),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_177),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_218),
.A2(n_157),
.B1(n_122),
.B2(n_201),
.Y(n_275)
);

HAxp5_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_205),
.CON(n_276),
.SN(n_276)
);

OAI21xp33_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_162),
.B(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_168),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_212),
.B(n_148),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_211),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_181),
.C(n_171),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_284),
.C(n_248),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_204),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_285),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_240),
.B(n_169),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_287),
.B(n_266),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_236),
.B1(n_212),
.B2(n_222),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_288),
.A2(n_300),
.B1(n_303),
.B2(n_309),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_252),
.A2(n_239),
.B(n_248),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_294),
.A2(n_315),
.B(n_261),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_162),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_307),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_243),
.B1(n_230),
.B2(n_216),
.Y(n_300)
);

XNOR2x2_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_119),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_301),
.A2(n_251),
.B(n_268),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_239),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_304),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_254),
.A2(n_243),
.B1(n_216),
.B2(n_232),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_215),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_232),
.B1(n_189),
.B2(n_203),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_179),
.B1(n_197),
.B2(n_165),
.Y(n_311)
);

AO21x2_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_266),
.B(n_285),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_258),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_316),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_314),
.B(n_317),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_273),
.A2(n_244),
.B(n_238),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_250),
.B(n_247),
.CI(n_228),
.CON(n_316),
.SN(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_244),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_274),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_250),
.B1(n_267),
.B2(n_271),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_325),
.A2(n_339),
.B1(n_309),
.B2(n_303),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_258),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_327),
.B(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_320),
.Y(n_329)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_329),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_253),
.B1(n_272),
.B2(n_257),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_312),
.B(n_296),
.Y(n_374)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_332),
.A2(n_343),
.B(n_349),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_336),
.B(n_347),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_256),
.Y(n_337)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_260),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_346),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_318),
.A2(n_266),
.B(n_280),
.Y(n_343)
);

OR2x4_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_266),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_302),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_286),
.B(n_270),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_348),
.A2(n_355),
.B1(n_305),
.B2(n_308),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_320),
.A2(n_280),
.B(n_265),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_351),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_253),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_354),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_305),
.A2(n_283),
.B(n_247),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_264),
.B(n_259),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_228),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_286),
.A2(n_234),
.B1(n_122),
.B2(n_238),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_356),
.A2(n_374),
.B1(n_339),
.B2(n_326),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_333),
.B(n_304),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_368),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_316),
.B1(n_301),
.B2(n_287),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_361),
.A2(n_381),
.B1(n_345),
.B2(n_351),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_294),
.C(n_315),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_375),
.C(n_334),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_288),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_306),
.Y(n_370)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_371),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_316),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_328),
.B1(n_355),
.B2(n_350),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_321),
.A2(n_308),
.B(n_289),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_377),
.A2(n_383),
.B(n_386),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_234),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_380),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_169),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_300),
.B1(n_312),
.B2(n_296),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_343),
.A2(n_264),
.B(n_259),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_180),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_387),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_349),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_398),
.Y(n_429)
);

XOR2x1_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_361),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_393),
.B(n_401),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_370),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_400),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_329),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_365),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_364),
.A2(n_339),
.B1(n_326),
.B2(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_339),
.B1(n_347),
.B2(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_388),
.A2(n_339),
.B1(n_323),
.B2(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_408),
.Y(n_430)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_383),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_335),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_415),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_354),
.C(n_346),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_413),
.C(n_414),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_412),
.A2(n_356),
.B1(n_374),
.B2(n_376),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_353),
.C(n_340),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_372),
.C(n_382),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_328),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_174),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_417),
.C(n_418),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_174),
.C(n_133),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_133),
.C(n_151),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_360),
.Y(n_420)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_388),
.B1(n_379),
.B2(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_424),
.B(n_426),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_377),
.C(n_389),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_414),
.B(n_363),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_428),
.B(n_439),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_440),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_407),
.B(n_366),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_434),
.B(n_398),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_396),
.B(n_416),
.Y(n_452)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_366),
.C(n_358),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_386),
.B1(n_371),
.B2(n_369),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_419),
.A2(n_413),
.B1(n_409),
.B2(n_393),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_133),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_415),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_445),
.B(n_453),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_446),
.B(n_452),
.Y(n_466)
);

OA21x2_ASAP7_75t_SL g447 ( 
.A1(n_436),
.A2(n_401),
.B(n_391),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_447),
.A2(n_427),
.B(n_420),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_430),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_411),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_459),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_443),
.A2(n_396),
.B1(n_417),
.B2(n_418),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_457),
.B1(n_438),
.B2(n_442),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_435),
.A2(n_76),
.B(n_59),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_435),
.B(n_425),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_45),
.C(n_46),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_461),
.C(n_462),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_151),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_180),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_425),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_151),
.C(n_49),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_64),
.C(n_60),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_448),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_465),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_431),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_426),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_474),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_421),
.Y(n_469)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_463),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_478),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_434),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_437),
.B1(n_441),
.B2(n_443),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_476),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_480),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_429),
.B(n_64),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_463),
.A2(n_27),
.B1(n_26),
.B2(n_48),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_460),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_485),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_469),
.A2(n_457),
.B1(n_452),
.B2(n_456),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_27),
.B1(n_26),
.B2(n_4),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_452),
.C(n_459),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_477),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_446),
.C(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_488),
.B(n_495),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_462),
.B(n_1),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_489),
.A2(n_478),
.B(n_474),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_48),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_467),
.B(n_50),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_496),
.B(n_11),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_497),
.A2(n_502),
.B1(n_505),
.B2(n_506),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_492),
.A2(n_477),
.B(n_466),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_498),
.B(n_500),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_48),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_504),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_483),
.A2(n_491),
.B(n_482),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_486),
.A2(n_26),
.B1(n_41),
.B2(n_4),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_50),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_508),
.C(n_41),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_484),
.A2(n_50),
.B1(n_47),
.B2(n_6),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_493),
.A3(n_489),
.B1(n_494),
.B2(n_485),
.C1(n_488),
.C2(n_41),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_513),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_11),
.B(n_3),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_511),
.C(n_508),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_50),
.C(n_47),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_515),
.B(n_507),
.Y(n_517)
);

AOI31xp67_ASAP7_75t_SL g521 ( 
.A1(n_517),
.A2(n_510),
.A3(n_3),
.B(n_6),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_519),
.B(n_512),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_50),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

AOI322xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_516),
.A3(n_3),
.B1(n_8),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_0),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_0),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_0),
.Y(n_526)
);


endmodule