module fake_jpeg_25649_n_296 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_20),
.B1(n_26),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_26),
.B1(n_20),
.B2(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_26),
.B1(n_27),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_25),
.B1(n_24),
.B2(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_60),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_36),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_28),
.B(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_33),
.B1(n_50),
.B2(n_47),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_47),
.Y(n_81)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_46),
.C(n_42),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_52),
.C(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_83),
.B1(n_90),
.B2(n_92),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_62),
.B1(n_67),
.B2(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_59),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_34),
.B1(n_35),
.B2(n_14),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_45),
.B1(n_29),
.B2(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_96),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_33),
.B1(n_29),
.B2(n_45),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_39),
.B1(n_47),
.B2(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_57),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_118),
.C(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_113),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_29),
.B1(n_45),
.B2(n_33),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_110),
.Y(n_148)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_95),
.B1(n_106),
.B2(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_66),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_71),
.B1(n_33),
.B2(n_66),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_29),
.B1(n_33),
.B2(n_55),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_27),
.B(n_18),
.C(n_22),
.D(n_13),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_120),
.C(n_90),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_68),
.C(n_72),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_22),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_27),
.C(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_68),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_74),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_74),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_130),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_134),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_85),
.B(n_77),
.C(n_91),
.D(n_94),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_149),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_78),
.B(n_80),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_142),
.B(n_22),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_146),
.B1(n_151),
.B2(n_56),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_80),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_75),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_104),
.B1(n_107),
.B2(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_92),
.B1(n_89),
.B2(n_71),
.Y(n_151)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_89),
.B(n_70),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_157),
.B(n_169),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_19),
.B(n_17),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_11),
.B(n_12),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_171),
.B1(n_145),
.B2(n_150),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_72),
.C(n_21),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_174),
.C(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_185),
.B(n_6),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_72),
.C(n_21),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_13),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_17),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_23),
.C(n_36),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_23),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_144),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_23),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_23),
.C(n_36),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_23),
.C(n_36),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_131),
.B1(n_136),
.B2(n_123),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_189),
.B1(n_196),
.B2(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_135),
.B1(n_132),
.B2(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_205),
.B1(n_176),
.B2(n_206),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_133),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_122),
.B1(n_137),
.B2(n_126),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_36),
.B1(n_22),
.B2(n_19),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_36),
.C(n_19),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_208),
.C(n_210),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_22),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_7),
.C(n_12),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_165),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_155),
.B1(n_160),
.B2(n_159),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_181),
.B1(n_157),
.B2(n_170),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_6),
.B1(n_11),
.B2(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_156),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_6),
.CI(n_11),
.CON(n_209),
.SN(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_5),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_174),
.C(n_177),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_213),
.C(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_162),
.C(n_183),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_158),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_5),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_162),
.C(n_182),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_167),
.B1(n_185),
.B2(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_229),
.B1(n_192),
.B2(n_154),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_166),
.C(n_163),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.C(n_12),
.Y(n_238)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_184),
.C(n_172),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_186),
.B1(n_188),
.B2(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_198),
.B1(n_197),
.B2(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_237),
.B1(n_224),
.B2(n_221),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_209),
.A3(n_210),
.B1(n_197),
.B2(n_199),
.C1(n_153),
.C2(n_171),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_243),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_209),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_238),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_0),
.C(n_1),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_4),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_4),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_236),
.B1(n_211),
.B2(n_237),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_223),
.C(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_227),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_220),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_234),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_233),
.B(n_242),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_260),
.B(n_3),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_233),
.B(n_230),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_3),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_245),
.B1(n_211),
.B2(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_245),
.B1(n_8),
.B2(n_2),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_8),
.B1(n_10),
.B2(n_2),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_0),
.C(n_1),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_247),
.C(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_249),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_276),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_251),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_278),
.B(n_3),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_265),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_3),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_282),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_265),
.B(n_259),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_283),
.B(n_286),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_266),
.C(n_269),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_9),
.C(n_10),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_8),
.C(n_9),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_290),
.B(n_10),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_284),
.B(n_11),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_289),
.C(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_0),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_1),
.Y(n_296)
);


endmodule