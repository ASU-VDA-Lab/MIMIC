module fake_jpeg_17952_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_241;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_29),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_13),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_66),
.B1(n_34),
.B2(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_21),
.B1(n_19),
.B2(n_14),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_12),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_30),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_86),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_80),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_37),
.B1(n_40),
.B2(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_56),
.B1(n_40),
.B2(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_43),
.C(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.C(n_69),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_48),
.C(n_65),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_97),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_92),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_96),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_11),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_72),
.A3(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_105),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_24),
.B(n_18),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_22),
.B1(n_44),
.B2(n_14),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_44),
.B1(n_14),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_77),
.B1(n_76),
.B2(n_71),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_77),
.B1(n_71),
.B2(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_83),
.B1(n_14),
.B2(n_16),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_44),
.B1(n_83),
.B2(n_22),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_128),
.B(n_24),
.Y(n_149)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

AND2x4_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_18),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_105),
.B1(n_94),
.B2(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_80),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_97),
.B(n_93),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_107),
.B(n_116),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_42),
.C(n_36),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_28),
.C(n_35),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_96),
.B1(n_16),
.B2(n_24),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_13),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_24),
.A3(n_12),
.B1(n_23),
.B2(n_25),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_23),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_23),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

NOR4xp25_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_117),
.C(n_119),
.D(n_112),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_52),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_108),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_162),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_173),
.B(n_149),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_127),
.B1(n_117),
.B2(n_68),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_161),
.A2(n_150),
.B1(n_134),
.B2(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_25),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_144),
.B(n_146),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_176),
.C(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_52),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_148),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_29),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_144),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_187),
.A2(n_194),
.B1(n_161),
.B2(n_171),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_147),
.B1(n_142),
.B2(n_131),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_166),
.B1(n_168),
.B2(n_144),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_142),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_130),
.C(n_141),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.C(n_164),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_140),
.C(n_129),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_172),
.B(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_129),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_144),
.B(n_17),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_196),
.B(n_17),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_153),
.B1(n_165),
.B2(n_168),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_185),
.B1(n_187),
.B2(n_189),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_203),
.C(n_211),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_162),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_213),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_54),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_29),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_184),
.B(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_177),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_185),
.B1(n_188),
.B2(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_220),
.A2(n_222),
.B1(n_197),
.B2(n_201),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_182),
.B1(n_181),
.B2(n_187),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_196),
.B(n_186),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_0),
.B(n_1),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_68),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_207),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_230),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_206),
.B1(n_199),
.B2(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_25),
.C(n_15),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_220),
.C(n_222),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_238),
.C(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_236),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_10),
.B(n_2),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_227),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_0),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_35),
.C(n_33),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_239),
.B(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_238),
.C(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_10),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_25),
.B(n_4),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_5),
.B(n_6),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_253),
.C(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_228),
.B(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_25),
.B(n_4),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_5),
.B(n_6),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_257),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_262),
.C(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_28),
.C(n_15),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_265),
.A3(n_258),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_5),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_15),
.C(n_20),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_20),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_267),
.B(n_6),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_15),
.C1(n_20),
.C2(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_9),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_20),
.B(n_15),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_15),
.C(n_20),
.Y(n_272)
);


endmodule