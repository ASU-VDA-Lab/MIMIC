module fake_jpeg_24617_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_22),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_17),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_14),
.B1(n_13),
.B2(n_9),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_28),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_20),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.C(n_21),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_36),
.B(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_12),
.B2(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_37),
.Y(n_53)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_41),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_37),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_10),
.C(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_57),
.B(n_44),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_62),
.C(n_10),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_43),
.A3(n_46),
.B1(n_47),
.B2(n_23),
.C1(n_3),
.C2(n_8),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_42),
.A3(n_56),
.B1(n_17),
.B2(n_25),
.C1(n_2),
.C2(n_7),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_62),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_67),
.C(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_60),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_69),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.C(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_2),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_1),
.C(n_75),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_1),
.Y(n_78)
);


endmodule