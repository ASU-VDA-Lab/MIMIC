module real_aes_1724_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_782, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_782;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g519 ( .A(n_0), .B(n_145), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_1), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_2), .B(n_127), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_3), .B(n_143), .Y(n_190) );
INVx1_ASAP7_75t_L g134 ( .A(n_4), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_5), .B(n_127), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g511 ( .A(n_6), .B(n_133), .Y(n_511) );
INVx1_ASAP7_75t_L g504 ( .A(n_7), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_8), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_9), .Y(n_756) );
AND2x2_ASAP7_75t_L g473 ( .A(n_10), .B(n_158), .Y(n_473) );
AND2x2_ASAP7_75t_L g192 ( .A(n_11), .B(n_177), .Y(n_192) );
AND2x2_ASAP7_75t_L g200 ( .A(n_12), .B(n_121), .Y(n_200) );
INVx2_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_14), .B(n_143), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_15), .Y(n_107) );
AOI221x1_ASAP7_75t_L g507 ( .A1(n_16), .A2(n_121), .B1(n_136), .B2(n_508), .C(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_17), .B(n_127), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_18), .B(n_127), .Y(n_171) );
INVx1_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_20), .A2(n_86), .B1(n_127), .B2(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_21), .A2(n_136), .B(n_477), .Y(n_476) );
AOI221xp5_ASAP7_75t_SL g486 ( .A1(n_22), .A2(n_36), .B1(n_127), .B2(n_136), .C(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_23), .B(n_145), .Y(n_478) );
OA21x2_ASAP7_75t_L g123 ( .A1(n_24), .A2(n_85), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g148 ( .A(n_24), .B(n_85), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_25), .B(n_143), .Y(n_498) );
INVxp67_ASAP7_75t_L g506 ( .A(n_26), .Y(n_506) );
AND2x2_ASAP7_75t_L g535 ( .A(n_27), .B(n_162), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_28), .A2(n_136), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_29), .A2(n_121), .B(n_125), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_30), .B(n_143), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_31), .A2(n_136), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_32), .B(n_143), .Y(n_155) );
AND2x2_ASAP7_75t_L g133 ( .A(n_33), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g137 ( .A(n_33), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g216 ( .A(n_33), .Y(n_216) );
OR2x6_ASAP7_75t_L g109 ( .A(n_34), .B(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_35), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_37), .B(n_127), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_38), .A2(n_78), .B1(n_136), .B2(n_214), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_39), .B(n_143), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_40), .B(n_127), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_41), .B(n_145), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_42), .A2(n_136), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_43), .B(n_145), .Y(n_239) );
AND2x2_ASAP7_75t_L g522 ( .A(n_44), .B(n_162), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_45), .B(n_162), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_46), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g130 ( .A(n_47), .Y(n_130) );
INVx1_ASAP7_75t_L g140 ( .A(n_47), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_48), .B(n_143), .Y(n_198) );
AND2x2_ASAP7_75t_L g161 ( .A(n_49), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_50), .B(n_127), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_51), .B(n_145), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_52), .B(n_145), .Y(n_154) );
AND2x2_ASAP7_75t_L g469 ( .A(n_53), .B(n_162), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_54), .B(n_127), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_55), .B(n_143), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_56), .B(n_127), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_57), .A2(n_136), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_58), .B(n_145), .Y(n_467) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_59), .B(n_158), .Y(n_499) );
AND2x2_ASAP7_75t_L g178 ( .A(n_60), .B(n_158), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_61), .A2(n_136), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_62), .B(n_143), .Y(n_479) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_63), .B(n_177), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_64), .B(n_145), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_65), .B(n_145), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_66), .A2(n_89), .B1(n_136), .B2(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_67), .B(n_143), .Y(n_174) );
INVx1_ASAP7_75t_L g132 ( .A(n_68), .Y(n_132) );
INVx1_ASAP7_75t_L g138 ( .A(n_68), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_69), .B(n_145), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_70), .A2(n_136), .B(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_71), .A2(n_136), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_72), .A2(n_136), .B(n_141), .Y(n_135) );
AND2x2_ASAP7_75t_L g157 ( .A(n_73), .B(n_158), .Y(n_157) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_74), .A2(n_99), .B1(n_749), .B2(n_760), .C1(n_772), .C2(n_774), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_74), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_74), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_75), .B(n_162), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_76), .B(n_127), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_77), .A2(n_80), .B1(n_127), .B2(n_208), .Y(n_570) );
INVx1_ASAP7_75t_L g112 ( .A(n_79), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_81), .B(n_145), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_82), .B(n_145), .Y(n_489) );
AND2x2_ASAP7_75t_L g240 ( .A(n_83), .B(n_177), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_84), .A2(n_136), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_87), .B(n_143), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_88), .A2(n_136), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_90), .B(n_143), .Y(n_238) );
BUFx2_ASAP7_75t_L g176 ( .A(n_91), .Y(n_176) );
INVxp67_ASAP7_75t_L g509 ( .A(n_92), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_93), .B(n_127), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_94), .A2(n_136), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_95), .B(n_143), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_96), .A2(n_100), .B1(n_745), .B2(n_747), .Y(n_744) );
BUFx2_ASAP7_75t_L g757 ( .A(n_97), .Y(n_757) );
BUFx2_ASAP7_75t_SL g778 ( .A(n_97), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_101), .B(n_744), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI21x1_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_113), .B(n_450), .Y(n_102) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx11_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_106), .A2(n_114), .B1(n_454), .B2(n_746), .Y(n_745) );
OR2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x6_ASAP7_75t_SL g453 ( .A(n_107), .B(n_109), .Y(n_453) );
OR2x2_ASAP7_75t_L g748 ( .A(n_107), .B(n_109), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_107), .B(n_108), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx4_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND3x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_328), .C(n_424), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_270), .C(n_297), .Y(n_115) );
OAI211xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_179), .B(n_219), .C(n_243), .Y(n_116) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_159), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_118), .A2(n_221), .B(n_225), .C(n_231), .Y(n_220) );
OR2x2_ASAP7_75t_L g343 ( .A(n_118), .B(n_280), .Y(n_343) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g310 ( .A(n_119), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_119), .B(n_281), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_119), .B(n_426), .Y(n_441) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_149), .Y(n_119) );
AND2x2_ASAP7_75t_L g227 ( .A(n_120), .B(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g247 ( .A(n_120), .Y(n_247) );
OR2x2_ASAP7_75t_L g262 ( .A(n_120), .B(n_169), .Y(n_262) );
INVx2_ASAP7_75t_L g268 ( .A(n_120), .Y(n_268) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_120), .Y(n_323) );
INVx1_ASAP7_75t_L g400 ( .A(n_120), .Y(n_400) );
INVx3_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_122), .A2(n_194), .B(n_200), .Y(n_193) );
AOI21x1_ASAP7_75t_L g515 ( .A1(n_122), .A2(n_516), .B(n_522), .Y(n_515) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_123), .Y(n_177) );
AND2x4_ASAP7_75t_L g147 ( .A(n_124), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_124), .B(n_148), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_135), .B(n_147), .Y(n_125) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_133), .Y(n_127) );
INVx1_ASAP7_75t_L g512 ( .A(n_128), .Y(n_512) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
AND2x6_ASAP7_75t_L g145 ( .A(n_129), .B(n_138), .Y(n_145) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g143 ( .A(n_131), .B(n_140), .Y(n_143) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx5_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
AND2x2_ASAP7_75t_L g139 ( .A(n_134), .B(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_134), .Y(n_211) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx3_ASAP7_75t_L g212 ( .A(n_137), .Y(n_212) );
INVx2_ASAP7_75t_L g218 ( .A(n_138), .Y(n_218) );
AND2x4_ASAP7_75t_L g214 ( .A(n_139), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_146), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_145), .B(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_146), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_146), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_146), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_146), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_146), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_146), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_146), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_146), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_146), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_146), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_146), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_146), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_147), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_147), .A2(n_475), .B(n_476), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_147), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_147), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_147), .B(n_509), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_147), .B(n_511), .C(n_512), .Y(n_510) );
NOR2x1_ASAP7_75t_SL g249 ( .A(n_149), .B(n_169), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_149), .B(n_268), .Y(n_279) );
AO21x1_ASAP7_75t_SL g149 ( .A1(n_150), .A2(n_151), .B(n_157), .Y(n_149) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_150), .A2(n_151), .B(n_157), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_158), .Y(n_162) );
OR2x2_ASAP7_75t_L g273 ( .A(n_159), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_159), .B(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g401 ( .A(n_159), .Y(n_401) );
NAND2x1_ASAP7_75t_L g159 ( .A(n_160), .B(n_169), .Y(n_159) );
OR2x2_ASAP7_75t_SL g261 ( .A(n_160), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g265 ( .A(n_160), .Y(n_265) );
INVx4_ASAP7_75t_L g281 ( .A(n_160), .Y(n_281) );
OR2x2_ASAP7_75t_L g296 ( .A(n_160), .B(n_229), .Y(n_296) );
AND2x2_ASAP7_75t_L g335 ( .A(n_160), .B(n_249), .Y(n_335) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_160), .Y(n_347) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_162), .Y(n_185) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_162), .A2(n_207), .B(n_213), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_162), .A2(n_235), .B(n_236), .Y(n_234) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_162), .A2(n_486), .B(n_490), .Y(n_485) );
AND2x2_ASAP7_75t_L g228 ( .A(n_169), .B(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g280 ( .A(n_169), .B(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g295 ( .A(n_169), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_169), .B(n_281), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_169), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g356 ( .A(n_169), .B(n_268), .Y(n_356) );
INVx2_ASAP7_75t_SL g426 ( .A(n_169), .Y(n_426) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_178), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_177), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_177), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_SL g568 ( .A(n_177), .Y(n_568) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp67_ASAP7_75t_L g180 ( .A(n_181), .B(n_201), .Y(n_180) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_181), .A2(n_298), .B(n_302), .C(n_318), .Y(n_297) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g393 ( .A(n_182), .B(n_232), .Y(n_393) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
INVx2_ASAP7_75t_L g242 ( .A(n_183), .Y(n_242) );
AND2x4_ASAP7_75t_SL g253 ( .A(n_183), .B(n_233), .Y(n_253) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_183), .Y(n_257) );
AND2x2_ASAP7_75t_L g315 ( .A(n_183), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g389 ( .A(n_183), .Y(n_389) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_184), .Y(n_291) );
AND2x2_ASAP7_75t_L g334 ( .A(n_184), .B(n_193), .Y(n_334) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_192), .Y(n_184) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_185), .A2(n_463), .B(n_469), .Y(n_462) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_185), .A2(n_529), .B(n_535), .Y(n_528) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_185), .A2(n_529), .B(n_535), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
INVx2_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
AND2x2_ASAP7_75t_L g284 ( .A(n_193), .B(n_233), .Y(n_284) );
INVx2_ASAP7_75t_L g316 ( .A(n_193), .Y(n_316) );
OR2x2_ASAP7_75t_L g339 ( .A(n_193), .B(n_204), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_201), .B(n_256), .Y(n_363) );
AND2x2_ASAP7_75t_L g397 ( .A(n_201), .B(n_333), .Y(n_397) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OAI31xp33_ASAP7_75t_SL g318 ( .A1(n_202), .A2(n_299), .A3(n_319), .B(n_326), .Y(n_318) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_203), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx3_ASAP7_75t_L g252 ( .A(n_204), .Y(n_252) );
AND2x2_ASAP7_75t_L g269 ( .A(n_204), .B(n_232), .Y(n_269) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x4_ASAP7_75t_L g259 ( .A(n_205), .B(n_206), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_208), .A2(n_214), .B1(n_503), .B2(n_505), .Y(n_502) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g404 ( .A(n_222), .Y(n_404) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2x1_ASAP7_75t_L g286 ( .A(n_224), .B(n_233), .Y(n_286) );
AND2x2_ASAP7_75t_L g327 ( .A(n_224), .B(n_242), .Y(n_327) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g307 ( .A(n_228), .B(n_265), .Y(n_307) );
AND2x2_ASAP7_75t_L g266 ( .A(n_229), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_229), .Y(n_275) );
INVx2_ASAP7_75t_L g325 ( .A(n_229), .Y(n_325) );
AND2x2_ASAP7_75t_L g415 ( .A(n_229), .B(n_400), .Y(n_415) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g421 ( .A(n_231), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_232), .B(n_241), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_232), .B(n_291), .Y(n_360) );
AND2x2_ASAP7_75t_L g408 ( .A(n_232), .B(n_334), .Y(n_408) );
INVx4_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g317 ( .A(n_233), .B(n_289), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_233), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g338 ( .A(n_233), .Y(n_338) );
BUFx2_ASAP7_75t_L g354 ( .A(n_233), .Y(n_354) );
AND2x4_ASAP7_75t_L g388 ( .A(n_233), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g433 ( .A(n_233), .B(n_334), .Y(n_433) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AOI222xp33_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_250), .B1(n_254), .B2(n_260), .C1(n_263), .C2(n_269), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_245), .A2(n_309), .B1(n_312), .B2(n_317), .Y(n_308) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g292 ( .A(n_246), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_SL g306 ( .A(n_246), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_246), .B(n_311), .Y(n_444) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g405 ( .A(n_247), .B(n_311), .Y(n_405) );
OR2x2_ASAP7_75t_L g382 ( .A(n_248), .B(n_264), .Y(n_382) );
OR2x2_ASAP7_75t_L g390 ( .A(n_248), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g374 ( .A(n_249), .B(n_267), .Y(n_374) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OR2x2_ASAP7_75t_L g282 ( .A(n_252), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g432 ( .A(n_252), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g383 ( .A(n_253), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_253), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g418 ( .A(n_253), .Y(n_418) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx2_ASAP7_75t_L g403 ( .A(n_256), .Y(n_403) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g305 ( .A(n_257), .B(n_284), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_258), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_258), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g407 ( .A(n_258), .B(n_279), .Y(n_407) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g341 ( .A(n_259), .B(n_327), .Y(n_341) );
AND2x2_ASAP7_75t_L g384 ( .A(n_259), .B(n_316), .Y(n_384) );
AND2x4_ASAP7_75t_L g299 ( .A(n_260), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g440 ( .A(n_262), .B(n_296), .Y(n_440) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_264), .B(n_279), .Y(n_423) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_265), .B(n_279), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_265), .A2(n_306), .B(n_407), .C(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_L g437 ( .A(n_265), .B(n_415), .Y(n_437) );
INVx1_ASAP7_75t_L g348 ( .A(n_266), .Y(n_348) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_269), .B(n_333), .Y(n_332) );
OAI21xp33_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_282), .B(n_285), .Y(n_270) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_273), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_281), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g373 ( .A(n_281), .Y(n_373) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_292), .Y(n_285) );
INVx1_ASAP7_75t_L g364 ( .A(n_286), .Y(n_364) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B(n_308), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
OR2x2_ASAP7_75t_L g349 ( .A(n_304), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g386 ( .A(n_304), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_304), .B(n_334), .Y(n_422) );
INVx1_ASAP7_75t_L g442 ( .A(n_305), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_307), .A2(n_410), .B1(n_413), .B2(n_416), .C(n_419), .Y(n_409) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI321xp33_ASAP7_75t_L g430 ( .A1(n_312), .A2(n_347), .A3(n_431), .B1(n_434), .B2(n_436), .C(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g371 ( .A(n_316), .Y(n_371) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g391 ( .A(n_322), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_352), .B1(n_356), .B2(n_357), .C(n_362), .Y(n_351) );
INVxp67_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
INVx1_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
NOR2xp67_ASAP7_75t_L g328 ( .A(n_329), .B(n_375), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_351), .C(n_366), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_336), .B2(n_342), .C(n_344), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g449 ( .A(n_334), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_337), .B(n_340), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_338), .B(n_384), .Y(n_429) );
INVx2_ASAP7_75t_SL g361 ( .A(n_339), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_340), .A2(n_345), .B1(n_346), .B2(n_349), .Y(n_344) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_348), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_349), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g355 ( .A(n_350), .Y(n_355) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_352), .A2(n_395), .B1(n_397), .B2(n_398), .C1(n_402), .C2(n_405), .Y(n_394) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_353), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g428 ( .A(n_353), .B(n_407), .Y(n_428) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_361), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_361), .B(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_365), .Y(n_362) );
NAND2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_372), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND4xp25_ASAP7_75t_SL g375 ( .A(n_376), .B(n_394), .C(n_406), .D(n_409), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B(n_383), .C(n_385), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_382), .A2(n_386), .B1(n_390), .B2(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_401), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_418), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_423), .Y(n_419) );
NOR4xp25_ASAP7_75t_L g424 ( .A(n_425), .B(n_430), .C(n_443), .D(n_445), .Y(n_424) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx3_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
CKINVDCx11_ASAP7_75t_R g746 ( .A(n_453), .Y(n_746) );
INVx4_ASAP7_75t_L g764 ( .A(n_454), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_454), .Y(n_765) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_683), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_576), .C(n_627), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_480), .B(n_523), .C(n_554), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_461), .B(n_528), .Y(n_691) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g536 ( .A(n_462), .B(n_472), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_462), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g553 ( .A(n_462), .B(n_543), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_462), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g590 ( .A(n_462), .B(n_566), .Y(n_590) );
INVx2_ASAP7_75t_L g616 ( .A(n_462), .Y(n_616) );
AND2x4_ASAP7_75t_L g625 ( .A(n_462), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g730 ( .A(n_462), .B(n_597), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .Y(n_463) );
AND2x2_ASAP7_75t_L g614 ( .A(n_470), .B(n_615), .Y(n_614) );
OAI32xp33_ASAP7_75t_L g697 ( .A1(n_470), .A2(n_619), .A3(n_623), .B1(n_630), .B2(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_470), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_552), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_471), .B(n_546), .C(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g650 ( .A(n_471), .B(n_553), .Y(n_650) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
INVx5_ASAP7_75t_L g575 ( .A(n_472), .Y(n_575) );
AND2x4_ASAP7_75t_L g631 ( .A(n_472), .B(n_543), .Y(n_631) );
OR2x2_ASAP7_75t_L g646 ( .A(n_472), .B(n_566), .Y(n_646) );
OR2x2_ASAP7_75t_L g672 ( .A(n_472), .B(n_528), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_472), .B(n_626), .Y(n_680) );
AND2x4_ASAP7_75t_SL g705 ( .A(n_472), .B(n_625), .Y(n_705) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_481), .B(n_625), .Y(n_701) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_482), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x6_ASAP7_75t_SL g525 ( .A(n_483), .B(n_526), .Y(n_525) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_484), .B(n_585), .Y(n_603) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_484), .Y(n_741) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g558 ( .A(n_485), .Y(n_558) );
AND2x2_ASAP7_75t_L g583 ( .A(n_485), .B(n_514), .Y(n_583) );
INVx2_ASAP7_75t_L g611 ( .A(n_485), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_485), .B(n_492), .Y(n_652) );
BUFx3_ASAP7_75t_L g676 ( .A(n_485), .Y(n_676) );
OR2x2_ASAP7_75t_L g688 ( .A(n_485), .B(n_492), .Y(n_688) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_485), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_491), .A2(n_719), .B1(n_722), .B2(n_723), .Y(n_718) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_500), .Y(n_491) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
OR2x2_ASAP7_75t_L g557 ( .A(n_492), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g564 ( .A(n_492), .Y(n_564) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_492), .B(n_501), .Y(n_581) );
AND2x4_ASAP7_75t_L g586 ( .A(n_492), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g595 ( .A(n_492), .Y(n_595) );
OR2x2_ASAP7_75t_L g601 ( .A(n_492), .B(n_501), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_492), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_492), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_492), .B(n_583), .Y(n_717) );
OR2x2_ASAP7_75t_L g733 ( .A(n_492), .B(n_636), .Y(n_733) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_500), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g559 ( .A(n_500), .Y(n_559) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_500), .B(n_550), .Y(n_666) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_501), .B(n_514), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_501), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_501), .B(n_558), .Y(n_562) );
INVx3_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
INVx1_ASAP7_75t_L g620 ( .A(n_501), .Y(n_620) );
AND2x2_ASAP7_75t_L g700 ( .A(n_501), .B(n_564), .Y(n_700) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_514), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g585 ( .A(n_514), .Y(n_585) );
AND2x2_ASAP7_75t_L g610 ( .A(n_514), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g636 ( .A(n_514), .B(n_558), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_514), .B(n_587), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_514), .Y(n_659) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
AOI222xp33_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_527), .B1(n_537), .B2(n_544), .C1(n_547), .C2(n_551), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_536), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_528), .B(n_597), .Y(n_648) );
AND2x4_ASAP7_75t_L g664 ( .A(n_528), .B(n_575), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_590), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g554 ( .A1(n_541), .A2(n_555), .B1(n_560), .B2(n_565), .C1(n_573), .C2(n_782), .Y(n_554) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g693 ( .A(n_542), .B(n_597), .Y(n_693) );
OR2x2_ASAP7_75t_L g736 ( .A(n_542), .B(n_642), .Y(n_736) );
AND2x2_ASAP7_75t_L g565 ( .A(n_543), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g626 ( .A(n_543), .Y(n_626) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_543), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_544), .A2(n_655), .B(n_660), .C(n_661), .Y(n_654) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g682 ( .A(n_546), .Y(n_682) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g612 ( .A(n_551), .Y(n_612) );
AND2x2_ASAP7_75t_L g596 ( .A(n_552), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g605 ( .A(n_552), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_555), .A2(n_573), .A3(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_556), .A2(n_606), .B(n_650), .C(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
OR2x2_ASAP7_75t_L g638 ( .A(n_557), .B(n_587), .Y(n_638) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
BUFx2_ASAP7_75t_L g606 ( .A(n_566), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_566), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_567), .Y(n_597) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_572), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_575), .B(n_632), .Y(n_724) );
OAI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_588), .B(n_591), .C(n_613), .Y(n_576) );
INVxp33_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_584), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_610), .Y(n_617) );
OR2x2_ASAP7_75t_L g593 ( .A(n_582), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g623 ( .A(n_582), .B(n_597), .Y(n_623) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g699 ( .A(n_583), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g722 ( .A(n_584), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_586), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_586), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g734 ( .A(n_586), .B(n_610), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_586), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g677 ( .A(n_587), .B(n_659), .Y(n_677) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AOI322xp5_ASAP7_75t_L g731 ( .A1(n_590), .A2(n_610), .A3(n_664), .B1(n_689), .B2(n_732), .C1(n_734), .C2(n_735), .Y(n_731) );
AOI211xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_596), .B(n_598), .C(n_607), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_594), .B(n_622), .Y(n_644) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g609 ( .A(n_595), .B(n_610), .Y(n_609) );
NOR2x1p5_ASAP7_75t_L g675 ( .A(n_595), .B(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_595), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_596), .A2(n_614), .B(n_617), .C(n_618), .Y(n_613) );
AND2x4_ASAP7_75t_L g632 ( .A(n_597), .B(n_616), .Y(n_632) );
INVx2_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_597), .B(n_631), .Y(n_662) );
AND2x2_ASAP7_75t_L g704 ( .A(n_597), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_597), .B(n_721), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_597), .B(n_625), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_604), .Y(n_598) );
AND2x2_ASAP7_75t_L g694 ( .A(n_600), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g622 ( .A(n_603), .Y(n_622) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_615), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g709 ( .A(n_615), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_621), .B(n_623), .C(n_624), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_622), .Y(n_706) );
INVx3_ASAP7_75t_SL g721 ( .A(n_625), .Y(n_721) );
NAND5xp2_ASAP7_75t_L g627 ( .A(n_628), .B(n_647), .C(n_654), .D(n_667), .E(n_678), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_633), .B1(n_637), .B2(n_639), .C1(n_643), .C2(n_645), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_630), .A2(n_711), .B1(n_715), .B2(n_716), .Y(n_710) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g660 ( .A(n_631), .B(n_632), .Y(n_660) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_641), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_642), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g679 ( .A(n_642), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g690 ( .A(n_642), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g720 ( .A(n_646), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g668 ( .A(n_653), .Y(n_668) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B(n_665), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_664), .A2(n_668), .B1(n_669), .B2(n_673), .Y(n_667) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_664), .Y(n_715) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g681 ( .A(n_666), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g686 ( .A(n_668), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_SL g714 ( .A(n_677), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_702), .C(n_725), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_701), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g726 ( .A(n_688), .B(n_714), .Y(n_726) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OAI321xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_706), .A3(n_707), .B1(n_709), .B2(n_710), .C(n_718), .Y(n_702) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_716), .A2(n_738), .B1(n_742), .B2(n_743), .Y(n_737) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI211xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_727), .B(n_731), .C(n_737), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_758), .Y(n_751) );
INVxp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_757), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_SL g773 ( .A(n_755), .B(n_757), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_755), .A2(n_776), .B(n_779), .Y(n_775) );
INVx1_ASAP7_75t_SL g767 ( .A(n_758), .Y(n_767) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx3_ASAP7_75t_L g770 ( .A(n_759), .Y(n_770) );
BUFx2_ASAP7_75t_L g780 ( .A(n_759), .Y(n_780) );
INVxp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_766), .B(n_768), .Y(n_761) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_769), .B(n_771), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
CKINVDCx8_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
endmodule