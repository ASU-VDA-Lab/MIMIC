module fake_jpeg_13630_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_5),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_47),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_55),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_17),
.B1(n_22),
.B2(n_13),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_21),
.Y(n_55)
);

FAx1_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_38),
.CI(n_32),
.CON(n_63),
.SN(n_63)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_20),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_74),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_40),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2x1_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_41),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_57),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_35),
.B1(n_45),
.B2(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_47),
.B1(n_54),
.B2(n_37),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_87),
.B(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_39),
.B1(n_31),
.B2(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_20),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_73),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_18),
.B1(n_3),
.B2(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_64),
.C(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_99),
.C(n_100),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_63),
.B(n_62),
.Y(n_95)
);

OAI211xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_89),
.B(n_92),
.C(n_80),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_82),
.B(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_84),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_77),
.C(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_68),
.C(n_18),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_67),
.C(n_66),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_86),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

XOR2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_111),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_95),
.C(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_6),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_119),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_105),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_104),
.B(n_106),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_114),
.B1(n_119),
.B2(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_128),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_12),
.B(n_6),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_121),
.B(n_124),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_125),
.A3(n_127),
.B1(n_128),
.B2(n_11),
.C1(n_12),
.C2(n_129),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_1),
.B(n_3),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_3),
.Y(n_133)
);


endmodule