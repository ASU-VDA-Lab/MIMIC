module fake_jpeg_14620_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_3),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_29),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_37),
.B1(n_30),
.B2(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_21),
.B1(n_14),
.B2(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_32),
.B1(n_31),
.B2(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_17),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_50),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_56),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_19),
.C(n_28),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_37),
.B1(n_36),
.B2(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_61),
.B1(n_67),
.B2(n_69),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_28),
.B1(n_15),
.B2(n_13),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_0),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_24),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_24),
.B(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_55),
.C(n_46),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_87),
.C(n_88),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_1),
.B(n_4),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_58),
.B1(n_18),
.B2(n_12),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_84),
.B1(n_65),
.B2(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_12),
.B1(n_19),
.B2(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_61),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_65),
.C(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_75),
.B(n_63),
.C(n_69),
.D(n_60),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_103),
.B(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_79),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_1),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_82),
.Y(n_109)
);

BUFx12f_ASAP7_75t_SL g105 ( 
.A(n_103),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_112),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_89),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_89),
.B(n_113),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_106),
.B1(n_105),
.B2(n_86),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_100),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_80),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_117),
.C(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_114),
.B(n_109),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_98),
.B(n_102),
.C(n_84),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_6),
.A3(n_8),
.B1(n_11),
.B2(n_117),
.C1(n_129),
.C2(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_131),
.C(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule