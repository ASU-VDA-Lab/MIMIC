module fake_jpeg_11308_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_54),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_56),
.Y(n_131)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_18),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_59),
.B(n_35),
.Y(n_169)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_79),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_22),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_78),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_0),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_97),
.Y(n_130)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_16),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_0),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_20),
.Y(n_134)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_21),
.B1(n_35),
.B2(n_27),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_23),
.B1(n_31),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_109),
.A2(n_163),
.B1(n_166),
.B2(n_27),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_68),
.A2(n_49),
.B1(n_37),
.B2(n_45),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_133),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_70),
.A2(n_49),
.B1(n_37),
.B2(n_45),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_49),
.B1(n_37),
.B2(n_42),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_59),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_136),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_46),
.B1(n_21),
.B2(n_53),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_161),
.B1(n_38),
.B2(n_36),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_84),
.A2(n_23),
.B1(n_42),
.B2(n_38),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_134),
.B(n_148),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_47),
.B(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_47),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_29),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_39),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_94),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_63),
.A2(n_33),
.B1(n_29),
.B2(n_40),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_58),
.A2(n_42),
.B1(n_23),
.B2(n_31),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_20),
.Y(n_189)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_177),
.Y(n_270)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_180),
.B(n_214),
.Y(n_266)
);

BUFx4f_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_185),
.B1(n_193),
.B2(n_232),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_75),
.B1(n_73),
.B2(n_90),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_183),
.A2(n_172),
.B1(n_138),
.B2(n_158),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_95),
.B1(n_87),
.B2(n_76),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_117),
.A2(n_41),
.B(n_39),
.C(n_20),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_187),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_264)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_188),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_190),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_116),
.B(n_33),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_191),
.B(n_201),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_117),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_192),
.B(n_205),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_194),
.Y(n_251)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_197),
.B(n_224),
.Y(n_267)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_131),
.B(n_31),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_200),
.A2(n_9),
.B(n_10),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_26),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_133),
.A2(n_26),
.B(n_109),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_207),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_279)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_221),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_111),
.B(n_38),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_164),
.A2(n_81),
.B1(n_36),
.B2(n_103),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_159),
.B1(n_124),
.B2(n_149),
.Y(n_245)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_137),
.B(n_36),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_227),
.B(n_236),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_118),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_119),
.A2(n_2),
.B(n_3),
.Y(n_229)
);

MAJx3_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_234),
.C(n_11),
.Y(n_274)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_113),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_233),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_121),
.A2(n_107),
.B1(n_104),
.B2(n_41),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_139),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_237),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_120),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_238),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_113),
.B1(n_122),
.B2(n_138),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_243),
.B1(n_271),
.B2(n_221),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_143),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_255),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_151),
.C(n_140),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_248),
.B(n_254),
.C(n_265),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_158),
.B1(n_143),
.B2(n_139),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_250),
.A2(n_262),
.B1(n_213),
.B2(n_211),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_146),
.C(n_123),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_185),
.B(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_175),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_293),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_261),
.B(n_192),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_184),
.A2(n_120),
.B1(n_5),
.B2(n_7),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_4),
.CI(n_5),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_234),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_264),
.B(n_233),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_9),
.C(n_10),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_268),
.A2(n_279),
.B(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_184),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_187),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_282),
.A2(n_263),
.B1(n_281),
.B2(n_249),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_196),
.B(n_14),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_217),
.B(n_14),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_246),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_303),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_183),
.B1(n_225),
.B2(n_230),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_297),
.A2(n_324),
.B1(n_328),
.B2(n_331),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_298),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

O2A1O1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_222),
.B(n_231),
.C(n_194),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_259),
.B(n_199),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_306),
.B(n_319),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_203),
.B(n_215),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_186),
.B1(n_208),
.B2(n_218),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_308),
.A2(n_316),
.B1(n_317),
.B2(n_326),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_266),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_254),
.C(n_261),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_242),
.C(n_294),
.Y(n_353)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_334),
.Y(n_347)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_210),
.B1(n_202),
.B2(n_198),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_244),
.A2(n_223),
.B1(n_181),
.B2(n_16),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_273),
.B(n_15),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_252),
.Y(n_320)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_321),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_329),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_181),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_332),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_244),
.A2(n_16),
.B1(n_250),
.B2(n_279),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_247),
.A2(n_16),
.B(n_268),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_325),
.A2(n_278),
.B(n_277),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_240),
.A2(n_267),
.B1(n_274),
.B2(n_272),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_264),
.B1(n_282),
.B2(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_264),
.A2(n_282),
.B1(n_293),
.B2(n_288),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_239),
.C(n_290),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_252),
.A2(n_282),
.B1(n_264),
.B2(n_275),
.Y(n_333)
);

AO21x2_ASAP7_75t_L g378 ( 
.A1(n_333),
.A2(n_258),
.B(n_253),
.Y(n_378)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_284),
.C(n_280),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_341),
.Y(n_373)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_241),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_345),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_286),
.A2(n_263),
.B1(n_284),
.B2(n_265),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_337),
.A2(n_340),
.B1(n_303),
.B2(n_307),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_275),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_342),
.Y(n_350)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_326),
.B1(n_316),
.B2(n_305),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_269),
.A2(n_258),
.B1(n_276),
.B2(n_253),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_246),
.B(n_292),
.C(n_249),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_257),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_344),
.Y(n_351)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_332),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_356),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_377),
.C(n_359),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_341),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_277),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_382),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_304),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_362),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_335),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_311),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_369),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_330),
.B(n_278),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_387),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_318),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_372),
.A2(n_299),
.B(n_320),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_321),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_375),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_242),
.C(n_294),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_378),
.A2(n_338),
.B1(n_314),
.B2(n_343),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_304),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_359),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_323),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_327),
.A2(n_317),
.B1(n_296),
.B2(n_297),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_312),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_324),
.A2(n_312),
.B1(n_337),
.B2(n_325),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_386),
.A2(n_299),
.B1(n_339),
.B2(n_312),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_313),
.B(n_344),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_350),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_391),
.A2(n_403),
.B1(n_407),
.B2(n_424),
.Y(n_442)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_379),
.B(n_308),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_394),
.B(n_398),
.Y(n_429)
);

NAND4xp25_ASAP7_75t_SL g395 ( 
.A(n_351),
.B(n_322),
.C(n_345),
.D(n_338),
.Y(n_395)
);

INVx8_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_350),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_382),
.B(n_339),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_399),
.A2(n_404),
.B(n_416),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_423),
.B1(n_378),
.B2(n_380),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_351),
.A2(n_334),
.B(n_354),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_353),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_386),
.B1(n_364),
.B2(n_378),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_408),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_411),
.B(n_398),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_413),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_366),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_418),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_357),
.B(n_371),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_415),
.B(n_417),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_354),
.A2(n_347),
.B(n_384),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_372),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_420),
.B(n_421),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_348),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_347),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_422),
.A2(n_389),
.B1(n_396),
.B2(n_391),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_360),
.A2(n_364),
.B1(n_349),
.B2(n_381),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_378),
.A2(n_360),
.B1(n_370),
.B2(n_349),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_431),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_419),
.A2(n_378),
.B1(n_370),
.B2(n_360),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_427),
.A2(n_444),
.B1(n_403),
.B2(n_409),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_373),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_373),
.C(n_377),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_433),
.B(n_435),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_370),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_438),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_380),
.C(n_352),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_436),
.A2(n_427),
.B1(n_424),
.B2(n_407),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_404),
.A2(n_367),
.B(n_352),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_388),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_410),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_446),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_388),
.C(n_376),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_448),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_423),
.A2(n_376),
.B1(n_408),
.B2(n_402),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_421),
.B(n_406),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_420),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_394),
.B(n_406),
.C(n_398),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_416),
.A2(n_422),
.B(n_397),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_450),
.A2(n_414),
.B(n_418),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_451),
.A2(n_412),
.B(n_415),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_455),
.B(n_431),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_400),
.Y(n_464)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_428),
.B(n_434),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_467),
.A2(n_468),
.B1(n_479),
.B2(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_445),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_478),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_413),
.B1(n_409),
.B2(n_390),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_471),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_395),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_399),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_473),
.A2(n_430),
.B(n_429),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_444),
.A2(n_450),
.B1(n_437),
.B2(n_442),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_480),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_392),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_455),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_477),
.B(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_451),
.A2(n_393),
.B1(n_432),
.B2(n_443),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_426),
.Y(n_494)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_448),
.CI(n_429),
.CON(n_485),
.SN(n_485)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_485),
.B(n_494),
.CI(n_489),
.CON(n_520),
.SN(n_520)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_428),
.B(n_441),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_489),
.A2(n_490),
.B(n_495),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_438),
.C(n_435),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_493),
.B(n_501),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_471),
.Y(n_498)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_449),
.C(n_475),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_503),
.B1(n_469),
.B2(n_461),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_476),
.B(n_465),
.Y(n_503)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_502),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_504),
.B(n_505),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_456),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_487),
.A2(n_476),
.B1(n_478),
.B2(n_459),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_506),
.B(n_507),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_474),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_515),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_458),
.C(n_462),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_516),
.C(n_514),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_487),
.A2(n_486),
.B1(n_491),
.B2(n_484),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_458),
.C(n_462),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_484),
.B(n_481),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_517),
.A2(n_521),
.B(n_485),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_500),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_520),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_496),
.B(n_482),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_509),
.A2(n_486),
.B1(n_491),
.B2(n_498),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_526),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_482),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_526),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_486),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_490),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_531),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_518),
.A2(n_495),
.B(n_499),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_529),
.A2(n_530),
.B(n_535),
.Y(n_536)
);

OAI221xp5_ASAP7_75t_L g530 ( 
.A1(n_517),
.A2(n_496),
.B1(n_492),
.B2(n_499),
.C(n_483),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_483),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_514),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_511),
.A2(n_498),
.B(n_492),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_534),
.B(n_518),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_539),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_533),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_541),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_515),
.Y(n_541)
);

INVx11_ASAP7_75t_L g543 ( 
.A(n_529),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_543),
.B(n_544),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_512),
.C(n_516),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_528),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_532),
.C(n_527),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_549),
.B(n_550),
.Y(n_553)
);

MAJx2_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_512),
.C(n_520),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_543),
.Y(n_552)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_552),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_546),
.Y(n_554)
);

AOI31xp33_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_553),
.A3(n_547),
.B(n_548),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_555),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_556),
.C(n_547),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_558),
.Y(n_559)
);

OAI321xp33_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_542),
.A3(n_536),
.B1(n_539),
.B2(n_523),
.C(n_544),
.Y(n_560)
);

NOR3xp33_ASAP7_75t_SL g561 ( 
.A(n_560),
.B(n_520),
.C(n_485),
.Y(n_561)
);


endmodule