module real_jpeg_17487_n_25 (n_17, n_8, n_0, n_157, n_21, n_168, n_2, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_159, n_161, n_162, n_169, n_167, n_23, n_11, n_14, n_160, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_25);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_159;
input n_161;
input n_162;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_131;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g103 ( 
.A(n_0),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_0),
.B(n_100),
.C(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_1),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_2),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_44),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_4),
.B(n_81),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_98),
.B(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_78),
.A3(n_90),
.B1(n_93),
.B2(n_126),
.C1(n_128),
.C2(n_168),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_8),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_10),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_96),
.C(n_119),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_16),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_17),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_18),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_19),
.B(n_67),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_20),
.B(n_74),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_22),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_31),
.B(n_94),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_149),
.B(n_155),
.Y(n_35)
);

OAI31xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_63),
.A3(n_131),
.B(n_135),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_49),
.C(n_56),
.Y(n_37)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_38),
.A2(n_49),
.A3(n_136),
.B1(n_137),
.B2(n_140),
.C(n_169),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

OAI322xp33_ASAP7_75t_L g140 ( 
.A1(n_39),
.A2(n_50),
.A3(n_141),
.B1(n_146),
.B2(n_147),
.C1(n_148),
.C2(n_170),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_42),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_43),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_47),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_102),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_56),
.B(n_142),
.C(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_62),
.Y(n_136)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI31xp67_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_72),
.A3(n_95),
.B(n_122),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.C(n_84),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_86),
.C(n_127),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_84),
.A3(n_123),
.B1(n_124),
.B2(n_125),
.C(n_167),
.Y(n_122)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_114),
.C(n_115),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_157),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_158),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_159),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_160),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_161),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_162),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_163),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_164),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_165),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_166),
.Y(n_120)
);


endmodule