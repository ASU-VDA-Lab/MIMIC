module fake_netlist_5_2241_n_1108 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1108);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1108;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_579;
wire n_204;
wire n_394;
wire n_250;
wire n_341;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1095;
wire n_976;
wire n_1096;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_482;
wire n_517;
wire n_342;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_599;
wire n_334;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_31),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_159),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_99),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_68),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_62),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_20),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_108),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_123),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_122),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_105),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_106),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_38),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_119),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_13),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_117),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_64),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_45),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_157),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_36),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_53),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_107),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_142),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_152),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_184),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_126),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_23),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_146),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_22),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_180),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_208),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_252),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_232),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_267),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_212),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_217),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_259),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_232),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_202),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_214),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_221),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_223),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_224),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_201),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_201),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_207),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_204),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_237),
.B1(n_205),
.B2(n_206),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_219),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_274),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OA22x2_ASAP7_75t_SL g328 ( 
.A1(n_280),
.A2(n_213),
.B1(n_222),
.B2(n_220),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_204),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_228),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_230),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_231),
.Y(n_338)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_234),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_207),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_294),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_205),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_271),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_240),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

AOI22x1_ASAP7_75t_L g363 ( 
.A1(n_313),
.A2(n_244),
.B1(n_256),
.B2(n_260),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_289),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_276),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

BUFx6f_ASAP7_75t_SL g377 ( 
.A(n_348),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_331),
.B(n_278),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_349),
.Y(n_381)
);

BUFx6f_ASAP7_75t_SL g382 ( 
.A(n_349),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_278),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_298),
.B1(n_311),
.B2(n_293),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_292),
.B1(n_270),
.B2(n_275),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_284),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_347),
.B(n_284),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_347),
.B(n_285),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_331),
.B(n_207),
.Y(n_398)
);

BUFx6f_ASAP7_75t_SL g399 ( 
.A(n_323),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_285),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_329),
.B(n_302),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_332),
.B(n_207),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_371),
.B(n_312),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_371),
.B(n_315),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_367),
.A2(n_273),
.B1(n_364),
.B2(n_322),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_371),
.B(n_206),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_350),
.A2(n_269),
.B1(n_266),
.B2(n_263),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_339),
.A2(n_233),
.B(n_226),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_353),
.B(n_236),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_327),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_332),
.B(n_238),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_336),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_353),
.B(n_332),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_374),
.B(n_209),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_374),
.B(n_209),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_374),
.A2(n_269),
.B1(n_266),
.B2(n_263),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_359),
.B(n_48),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_239),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_325),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_330),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_367),
.A2(n_210),
.B1(n_261),
.B2(n_258),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_326),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_359),
.B(n_242),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_320),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_326),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_320),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_373),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_372),
.C(n_362),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_373),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_428),
.B(n_400),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_373),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_373),
.C(n_372),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_373),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_353),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_379),
.B(n_330),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_353),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_352),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_321),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_385),
.A2(n_366),
.B1(n_359),
.B2(n_321),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_380),
.B(n_323),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_358),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_434),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_322),
.Y(n_471)
);

AND2x6_ASAP7_75t_SL g472 ( 
.A(n_425),
.B(n_328),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_395),
.B(n_352),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_358),
.Y(n_476)
);

INVx8_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NOR3xp33_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_358),
.C(n_339),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_403),
.B(n_368),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_403),
.B(n_358),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_363),
.C(n_352),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_403),
.B(n_358),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_422),
.B(n_323),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_425),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_437),
.B(n_323),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_425),
.B(n_323),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_443),
.B(n_383),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_443),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_423),
.A2(n_338),
.B(n_354),
.C(n_360),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_423),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_366),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_443),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_401),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_429),
.B(n_366),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_432),
.B(n_210),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_433),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_377),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_338),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_338),
.Y(n_501)
);

NOR3xp33_ASAP7_75t_L g502 ( 
.A(n_407),
.B(n_357),
.C(n_351),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_375),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_338),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_351),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_410),
.B(n_357),
.Y(n_507)
);

BUFx6f_ASAP7_75t_SL g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_378),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_386),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_441),
.B(n_245),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_383),
.B(n_338),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_390),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_393),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_399),
.A2(n_249),
.B1(n_254),
.B2(n_250),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_406),
.A2(n_333),
.B(n_324),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_384),
.B(n_355),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_384),
.B(n_355),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_399),
.A2(n_377),
.B1(n_436),
.B2(n_382),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_388),
.B(n_355),
.Y(n_527)
);

INVx8_ASAP7_75t_L g528 ( 
.A(n_382),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_388),
.B(n_355),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_414),
.B(n_361),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_389),
.B(n_355),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_389),
.B(n_355),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_523),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_455),
.B(n_463),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_504),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_467),
.Y(n_537)
);

AO22x2_ASAP7_75t_L g538 ( 
.A1(n_507),
.A2(n_451),
.B1(n_457),
.B2(n_481),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_361),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_414),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_457),
.A2(n_328),
.B1(n_363),
.B2(n_436),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_484),
.B(n_436),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_469),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_361),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_497),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_494),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_509),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_489),
.B(n_436),
.Y(n_553)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_499),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_513),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_454),
.B(n_405),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_493),
.B(n_503),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_454),
.B(n_405),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_519),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_464),
.B(n_408),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_519),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_461),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_471),
.A2(n_377),
.B1(n_399),
.B2(n_354),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_450),
.B(n_408),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_458),
.B(n_419),
.Y(n_570)
);

NOR4xp25_ASAP7_75t_SL g571 ( 
.A(n_514),
.B(n_262),
.C(n_419),
.D(n_397),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_498),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_475),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_458),
.B(n_406),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_453),
.B(n_365),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_453),
.B(n_426),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_511),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_512),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_521),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_468),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_476),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_502),
.B(n_488),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_480),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

BUFx8_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_478),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_460),
.Y(n_591)
);

OAI221xp5_ASAP7_75t_L g592 ( 
.A1(n_471),
.A2(n_354),
.B1(n_346),
.B2(n_360),
.C(n_365),
.Y(n_592)
);

AO22x2_ASAP7_75t_L g593 ( 
.A1(n_502),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_517),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_417),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_473),
.A2(n_376),
.B1(n_418),
.B2(n_415),
.Y(n_598)
);

OAI221xp5_ASAP7_75t_L g599 ( 
.A1(n_496),
.A2(n_346),
.B1(n_360),
.B2(n_365),
.C(n_324),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_540),
.B(n_496),
.C(n_495),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_540),
.A2(n_508),
.B1(n_487),
.B2(n_466),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_563),
.A2(n_452),
.B(n_483),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_578),
.B(n_559),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_578),
.A2(n_462),
.B(n_483),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_535),
.B(n_492),
.Y(n_606)
);

BUFx12f_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_563),
.A2(n_486),
.B(n_487),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_547),
.B(n_492),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_549),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_562),
.B(n_495),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_570),
.A2(n_486),
.B(n_479),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_479),
.B(n_459),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_565),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_465),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_478),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_522),
.B1(n_518),
.B2(n_466),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_573),
.B(n_499),
.Y(n_619)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_575),
.A2(n_530),
.B(n_532),
.Y(n_620)
);

NOR2x1_ASAP7_75t_L g621 ( 
.A(n_567),
.B(n_527),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_575),
.A2(n_525),
.B(n_524),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_539),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_594),
.A2(n_531),
.B(n_529),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_538),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_591),
.B(n_477),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_597),
.A2(n_490),
.B(n_527),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_538),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_534),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_543),
.B(n_477),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_587),
.A2(n_528),
.B(n_477),
.C(n_472),
.Y(n_632)
);

OA22x2_ASAP7_75t_L g633 ( 
.A1(n_537),
.A2(n_545),
.B1(n_544),
.B2(n_546),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_553),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_548),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_583),
.B(n_528),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_595),
.B(n_528),
.Y(n_637)
);

AO21x1_ASAP7_75t_L g638 ( 
.A1(n_541),
.A2(n_447),
.B(n_439),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_596),
.A2(n_404),
.B(n_396),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_568),
.A2(n_416),
.B(n_392),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_553),
.A2(n_404),
.B(n_412),
.C(n_396),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_558),
.A2(n_430),
.B(n_417),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_567),
.A2(n_396),
.B1(n_404),
.B2(n_424),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_558),
.B(n_412),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_560),
.B(n_412),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_554),
.B(n_344),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_555),
.Y(n_649)
);

O2A1O1Ixp33_ASAP7_75t_SL g650 ( 
.A1(n_560),
.A2(n_424),
.B(n_430),
.C(n_427),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_589),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_589),
.B(n_344),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_566),
.B(n_569),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_576),
.A2(n_427),
.B1(n_426),
.B2(n_424),
.Y(n_655)
);

BUFx8_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_542),
.A2(n_355),
.B(n_342),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_599),
.A2(n_596),
.B(n_561),
.C(n_557),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_568),
.B(n_577),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_610),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_609),
.A2(n_599),
.B1(n_598),
.B2(n_542),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_579),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_621),
.B(n_550),
.Y(n_663)
);

BUFx4f_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_626),
.B(n_629),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_601),
.B(n_580),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_633),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_630),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_635),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_604),
.A2(n_590),
.B1(n_593),
.B2(n_581),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_606),
.B(n_582),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_642),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_649),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_612),
.B(n_533),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_611),
.B(n_551),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_652),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_624),
.B(n_618),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_659),
.B(n_593),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_624),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_634),
.Y(n_682)
);

INVx3_ASAP7_75t_SL g683 ( 
.A(n_624),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_651),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_617),
.B(n_592),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_636),
.B(n_592),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_616),
.B(n_590),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_637),
.B(n_590),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_600),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_656),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_602),
.A2(n_541),
.B1(n_571),
.B2(n_426),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_SL g692 ( 
.A1(n_605),
.A2(n_571),
.B(n_427),
.C(n_446),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_615),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_634),
.B(n_344),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_619),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_654),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_648),
.B(n_392),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_656),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_627),
.Y(n_700)
);

AND3x1_ASAP7_75t_SL g701 ( 
.A(n_632),
.B(n_3),
.C(n_4),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_658),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_646),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_L g704 ( 
.A1(n_653),
.A2(n_342),
.B1(n_333),
.B2(n_343),
.C(n_345),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_643),
.B(n_608),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_631),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_608),
.B(n_345),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_655),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_644),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_622),
.B(n_345),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_620),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_641),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_613),
.B(n_343),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_639),
.B(n_392),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_706),
.A2(n_603),
.B(n_613),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_680),
.B(n_670),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_702),
.A2(n_603),
.B1(n_614),
.B2(n_628),
.Y(n_718)
);

BUFx2_ASAP7_75t_SL g719 ( 
.A(n_667),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_660),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_665),
.B(n_689),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_657),
.B(n_650),
.C(n_638),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_685),
.B(n_628),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_665),
.B(n_3),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_689),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_670),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_698),
.A2(n_614),
.B(n_625),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_664),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_705),
.B(n_625),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_675),
.B(n_622),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_666),
.B(n_640),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_683),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_678),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_700),
.A2(n_640),
.B1(n_421),
.B2(n_416),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_673),
.B(n_4),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_693),
.B(n_5),
.Y(n_737)
);

O2A1O1Ixp5_ASAP7_75t_SL g738 ( 
.A1(n_691),
.A2(n_340),
.B(n_334),
.C(n_7),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_683),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_706),
.A2(n_421),
.B(n_416),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_667),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_711),
.A2(n_421),
.B(n_416),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_678),
.Y(n_743)
);

CKINVDCx11_ASAP7_75t_R g744 ( 
.A(n_696),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_690),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_700),
.A2(n_421),
.B1(n_416),
.B2(n_392),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_678),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_671),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_688),
.A2(n_340),
.B(n_326),
.C(n_334),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_671),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_710),
.A2(n_421),
.B1(n_392),
.B2(n_369),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_693),
.B(n_5),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_664),
.B(n_334),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_668),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_664),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_695),
.B(n_6),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_674),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_681),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_710),
.A2(n_369),
.B1(n_340),
.B2(n_334),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_336),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_681),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_684),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_682),
.B(n_49),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_703),
.B(n_6),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_692),
.A2(n_661),
.B(n_712),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_672),
.A2(n_369),
.B1(n_340),
.B2(n_334),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_703),
.B(n_7),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_712),
.A2(n_340),
.B(n_336),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_669),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_682),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_663),
.A2(n_676),
.B(n_714),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_663),
.A2(n_341),
.B(n_336),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_682),
.B(n_713),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_682),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_662),
.B(n_8),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_690),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_663),
.A2(n_341),
.B(n_336),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_669),
.B(n_8),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_687),
.B(n_10),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_677),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_677),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_720),
.B(n_697),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_732),
.B(n_713),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_721),
.B(n_714),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_748),
.B(n_708),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_731),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_717),
.B(n_707),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_782),
.B(n_708),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_725),
.A2(n_699),
.B1(n_713),
.B2(n_709),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_750),
.B(n_677),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_758),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_739),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_764),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_733),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_724),
.B(n_694),
.Y(n_798)
);

AOI211xp5_ASAP7_75t_L g799 ( 
.A1(n_781),
.A2(n_701),
.B(n_699),
.C(n_704),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_SL g801 ( 
.A1(n_727),
.A2(n_694),
.B(n_715),
.C(n_12),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_777),
.B(n_10),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_751),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_723),
.A2(n_761),
.B(n_736),
.C(n_766),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_726),
.B(n_715),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_772),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_730),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_751),
.B(n_715),
.Y(n_808)
);

INVx3_ASAP7_75t_SL g809 ( 
.A(n_745),
.Y(n_809)
);

O2A1O1Ixp5_ASAP7_75t_L g810 ( 
.A1(n_767),
.A2(n_773),
.B(n_716),
.C(n_768),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_723),
.B(n_11),
.Y(n_811)
);

BUFx2_ASAP7_75t_R g812 ( 
.A(n_745),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_755),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_769),
.B(n_11),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_761),
.A2(n_341),
.B(n_336),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_755),
.B(n_12),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_771),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_783),
.B(n_771),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_729),
.B(n_13),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_783),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_780),
.B(n_14),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_742),
.A2(n_341),
.B(n_14),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_SL g823 ( 
.A1(n_718),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_737),
.B(n_15),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_753),
.B(n_16),
.Y(n_825)
);

AND2x4_ASAP7_75t_SL g826 ( 
.A(n_728),
.B(n_341),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_744),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_734),
.B(n_369),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_782),
.B(n_17),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_SL g830 ( 
.A1(n_718),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_759),
.B(n_18),
.Y(n_831)
);

OA21x2_ASAP7_75t_L g832 ( 
.A1(n_740),
.A2(n_341),
.B(n_19),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_722),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_734),
.B(n_50),
.Y(n_834)
);

O2A1O1Ixp5_ASAP7_75t_L g835 ( 
.A1(n_735),
.A2(n_752),
.B(n_760),
.C(n_746),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_757),
.B(n_51),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_749),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_756),
.A2(n_369),
.B1(n_341),
.B2(n_26),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_765),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_756),
.A2(n_369),
.B1(n_28),
.B2(n_29),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_744),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_741),
.A2(n_369),
.B1(n_29),
.B2(n_30),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_799),
.A2(n_747),
.B1(n_743),
.B2(n_741),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_833),
.A2(n_747),
.B1(n_775),
.B2(n_728),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_811),
.A2(n_778),
.B1(n_728),
.B2(n_765),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_833),
.A2(n_728),
.B1(n_765),
.B2(n_754),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_794),
.Y(n_848)
);

OAI21xp33_ASAP7_75t_L g849 ( 
.A1(n_839),
.A2(n_738),
.B(n_772),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_811),
.A2(n_763),
.B1(n_776),
.B2(n_762),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_786),
.B(n_788),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_834),
.A2(n_776),
.B1(n_762),
.B2(n_763),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_SL g854 ( 
.A1(n_809),
.A2(n_754),
.B1(n_30),
.B2(n_31),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_802),
.A2(n_770),
.B1(n_32),
.B2(n_33),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_814),
.A2(n_791),
.B1(n_827),
.B2(n_841),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_785),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_785),
.B(n_779),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_804),
.B(n_774),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_807),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_786),
.B(n_27),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_798),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_798),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_788),
.B(n_39),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_819),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_818),
.B(n_40),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_793),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_793),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_789),
.B(n_41),
.Y(n_869)
);

AOI21xp33_ASAP7_75t_L g870 ( 
.A1(n_823),
.A2(n_42),
.B(n_43),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_839),
.A2(n_369),
.B1(n_44),
.B2(n_43),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_800),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_837),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_837),
.A2(n_797),
.B1(n_795),
.B2(n_784),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_818),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_842),
.A2(n_840),
.B1(n_821),
.B2(n_824),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_831),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_809),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_803),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_836),
.A2(n_199),
.B1(n_63),
.B2(n_65),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_806),
.Y(n_881)
);

OAI22xp33_ASAP7_75t_L g882 ( 
.A1(n_825),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_SL g883 ( 
.A1(n_821),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_806),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_824),
.A2(n_816),
.B1(n_817),
.B2(n_829),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_SL g887 ( 
.A1(n_829),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_792),
.B(n_198),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_816),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_852),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_866),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_854),
.A2(n_812),
.B1(n_832),
.B2(n_843),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_845),
.A2(n_857),
.B(n_873),
.C(n_871),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_875),
.B(n_792),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_867),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_851),
.B(n_843),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_848),
.Y(n_897)
);

OAI211xp5_ASAP7_75t_SL g898 ( 
.A1(n_857),
.A2(n_810),
.B(n_830),
.C(n_823),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_865),
.A2(n_830),
.B1(n_801),
.B2(n_838),
.C(n_787),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_860),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_867),
.B(n_790),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_SL g902 ( 
.A1(n_874),
.A2(n_801),
.B(n_815),
.C(n_813),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_884),
.Y(n_903)
);

AO32x2_ASAP7_75t_L g904 ( 
.A1(n_844),
.A2(n_832),
.A3(n_822),
.B1(n_805),
.B2(n_787),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_877),
.B(n_805),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_870),
.A2(n_835),
.B(n_828),
.C(n_790),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_881),
.Y(n_907)
);

OA21x2_ASAP7_75t_L g908 ( 
.A1(n_859),
.A2(n_808),
.B(n_813),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_879),
.Y(n_909)
);

AO21x1_ASAP7_75t_L g910 ( 
.A1(n_856),
.A2(n_790),
.B(n_808),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_855),
.A2(n_832),
.B(n_822),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_855),
.A2(n_822),
.B(n_803),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_868),
.B(n_826),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_858),
.A2(n_826),
.B(n_80),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_79),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_885),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_889),
.A2(n_82),
.B(n_83),
.C(n_84),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_885),
.B(n_85),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_886),
.B(n_86),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_896),
.B(n_858),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_908),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_897),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_900),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_890),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_905),
.B(n_886),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_903),
.Y(n_926)
);

OAI222xp33_ASAP7_75t_L g927 ( 
.A1(n_919),
.A2(n_846),
.B1(n_876),
.B2(n_850),
.C1(n_863),
.C2(n_862),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_890),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_916),
.B(n_850),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_916),
.B(n_861),
.Y(n_931)
);

CKINVDCx14_ASAP7_75t_R g932 ( 
.A(n_895),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_908),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_894),
.B(n_888),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_907),
.B(n_853),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_909),
.B(n_916),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_901),
.B(n_864),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_916),
.B(n_869),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_910),
.B(n_849),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_904),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_911),
.B(n_862),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_904),
.B(n_863),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_921),
.A2(n_912),
.B(n_893),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_921),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_929),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_921),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_930),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_941),
.A2(n_893),
.B(n_917),
.C(n_906),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_933),
.A2(n_914),
.B(n_913),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_928),
.Y(n_950)
);

OA21x2_ASAP7_75t_L g951 ( 
.A1(n_928),
.A2(n_940),
.B(n_939),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_940),
.A2(n_902),
.B(n_898),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_933),
.A2(n_914),
.B(n_847),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_928),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_924),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_941),
.A2(n_902),
.B(n_917),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_933),
.A2(n_904),
.B(n_899),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_933),
.B(n_895),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_924),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_927),
.A2(n_906),
.B(n_889),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_947),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_960),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_947),
.B(n_935),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_951),
.B(n_942),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_947),
.B(n_935),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_956),
.B(n_938),
.Y(n_968)
);

NOR2x1_ASAP7_75t_L g969 ( 
.A(n_956),
.B(n_922),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_944),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_961),
.B(n_892),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_945),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_953),
.B(n_930),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_944),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_962),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_971),
.A2(n_961),
.B1(n_932),
.B2(n_943),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_972),
.Y(n_977)
);

OR2x2_ASAP7_75t_SL g978 ( 
.A(n_971),
.B(n_943),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_963),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_969),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_971),
.A2(n_943),
.B1(n_942),
.B2(n_952),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_965),
.B(n_952),
.Y(n_982)
);

OAI322xp33_ASAP7_75t_L g983 ( 
.A1(n_976),
.A2(n_966),
.A3(n_964),
.B1(n_958),
.B2(n_954),
.C1(n_974),
.C2(n_970),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_977),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_967),
.Y(n_985)
);

AND2x4_ASAP7_75t_SL g986 ( 
.A(n_980),
.B(n_931),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_981),
.B(n_968),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_979),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_986),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_985),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_987),
.B(n_981),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_984),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_988),
.Y(n_993)
);

NOR2x1p5_ASAP7_75t_L g994 ( 
.A(n_983),
.B(n_982),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_983),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_984),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_987),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_988),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_990),
.Y(n_999)
);

AOI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_995),
.A2(n_980),
.B1(n_966),
.B2(n_948),
.C(n_978),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_991),
.A2(n_948),
.B(n_973),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_990),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_998),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_997),
.A2(n_943),
.B(n_957),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

OAI32xp33_ASAP7_75t_L g1006 ( 
.A1(n_989),
.A2(n_958),
.A3(n_974),
.B1(n_970),
.B2(n_946),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_992),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_993),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1005),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1003),
.B(n_994),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1006),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_1000),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1001),
.B(n_996),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_1004),
.B(n_996),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1009),
.B(n_973),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_1013),
.B(n_958),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_952),
.B1(n_954),
.B2(n_882),
.C(n_872),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_1007),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1010),
.A2(n_957),
.B(n_951),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1011),
.A2(n_952),
.B1(n_946),
.B2(n_944),
.C(n_950),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1008),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1018),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1021),
.B(n_1014),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1015),
.B(n_951),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_943),
.B1(n_957),
.B2(n_952),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1016),
.B(n_951),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_1020),
.Y(n_1027)
);

AND2x2_ASAP7_75t_SL g1028 ( 
.A(n_1019),
.B(n_915),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_SL g1029 ( 
.A(n_1018),
.B(n_951),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1018),
.A2(n_950),
.B(n_946),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1018),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1029),
.Y(n_1032)
);

AOI222xp33_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_891),
.B1(n_950),
.B2(n_925),
.C1(n_878),
.C2(n_953),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1022),
.B(n_883),
.C(n_887),
.Y(n_1034)
);

AOI211xp5_ASAP7_75t_L g1035 ( 
.A1(n_1031),
.A2(n_918),
.B(n_953),
.C(n_949),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_1023),
.A2(n_955),
.B(n_918),
.C(n_959),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1025),
.B(n_880),
.C(n_918),
.D(n_930),
.Y(n_1037)
);

OAI211xp5_ASAP7_75t_L g1038 ( 
.A1(n_1025),
.A2(n_949),
.B(n_955),
.C(n_920),
.Y(n_1038)
);

AOI211x1_ASAP7_75t_SL g1039 ( 
.A1(n_1026),
.A2(n_1030),
.B(n_1028),
.C(n_1024),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1029),
.Y(n_1040)
);

OAI221xp5_ASAP7_75t_SL g1041 ( 
.A1(n_1025),
.A2(n_936),
.B1(n_959),
.B2(n_945),
.C(n_937),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1032),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1038),
.A2(n_949),
.B(n_937),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1041),
.B(n_959),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1034),
.A2(n_891),
.B1(n_936),
.B2(n_931),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1033),
.B(n_931),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1048),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_1047),
.B(n_1037),
.Y(n_1050)
);

AOI31xp33_ASAP7_75t_L g1051 ( 
.A1(n_1042),
.A2(n_1035),
.A3(n_1036),
.B(n_930),
.Y(n_1051)
);

XOR2xp5_ASAP7_75t_L g1052 ( 
.A(n_1043),
.B(n_931),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1046),
.A2(n_926),
.B1(n_923),
.B2(n_922),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1045),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_923),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_1047),
.B(n_926),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1042),
.Y(n_1057)
);

XNOR2xp5_ASAP7_75t_L g1058 ( 
.A(n_1048),
.B(n_87),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1058),
.A2(n_1049),
.B(n_1052),
.Y(n_1059)
);

NOR2x1p5_ASAP7_75t_L g1060 ( 
.A(n_1057),
.B(n_934),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1050),
.B(n_934),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_1054),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1051),
.A2(n_88),
.B(n_90),
.C(n_91),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_1056),
.Y(n_1064)
);

AND2x2_ASAP7_75t_SL g1065 ( 
.A(n_1055),
.B(n_93),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1053),
.A2(n_94),
.B(n_96),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1058),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1062),
.A2(n_904),
.B1(n_98),
.B2(n_100),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1061),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1065),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1064),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1067),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1063),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1059),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_1066),
.B(n_103),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1061),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1064),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_1062),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1061),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1069),
.Y(n_1082)
);

NAND5xp2_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_113),
.C(n_114),
.D(n_115),
.E(n_118),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1077),
.A2(n_120),
.B(n_125),
.C(n_127),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_1070),
.A2(n_128),
.B(n_129),
.Y(n_1085)
);

OAI211xp5_ASAP7_75t_L g1086 ( 
.A1(n_1078),
.A2(n_1072),
.B(n_1075),
.C(n_1073),
.Y(n_1086)
);

OAI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1071),
.A2(n_197),
.B1(n_131),
.B2(n_132),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1076),
.Y(n_1088)
);

AOI311xp33_ASAP7_75t_L g1089 ( 
.A1(n_1086),
.A2(n_1074),
.A3(n_1082),
.B(n_1088),
.C(n_1084),
.Y(n_1089)
);

AND3x4_ASAP7_75t_L g1090 ( 
.A(n_1083),
.B(n_1068),
.C(n_134),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_1085),
.B(n_1081),
.C(n_1087),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1082),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_1086),
.B(n_137),
.C(n_139),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_1086),
.B(n_140),
.C(n_141),
.Y(n_1094)
);

AOI221xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1089),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.C(n_147),
.Y(n_1095)
);

NAND4xp25_ASAP7_75t_SL g1096 ( 
.A(n_1094),
.B(n_148),
.C(n_149),
.D(n_150),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1093),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_1097)
);

AO22x2_ASAP7_75t_L g1098 ( 
.A1(n_1095),
.A2(n_1091),
.B1(n_1090),
.B2(n_1092),
.Y(n_1098)
);

AOI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_1097),
.B(n_1096),
.Y(n_1099)
);

XOR2xp5_ASAP7_75t_L g1100 ( 
.A(n_1099),
.B(n_158),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_160),
.B(n_161),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1101),
.B(n_162),
.Y(n_1102)
);

XOR2xp5_ASAP7_75t_L g1103 ( 
.A(n_1100),
.B(n_164),
.Y(n_1103)
);

OAI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_1100),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.C1(n_168),
.C2(n_170),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1102),
.A2(n_172),
.B(n_173),
.Y(n_1105)
);

OA22x2_ASAP7_75t_L g1106 ( 
.A1(n_1103),
.A2(n_1104),
.B1(n_176),
.B2(n_177),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1106),
.A2(n_175),
.B1(n_179),
.B2(n_181),
.Y(n_1107)
);

AOI211xp5_ASAP7_75t_L g1108 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_182),
.C(n_183),
.Y(n_1108)
);


endmodule