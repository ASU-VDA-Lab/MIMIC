module fake_netlist_6_837_n_2334 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2334);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2334;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_1159;
wire n_276;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g226 ( 
.A(n_93),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_80),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_16),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_224),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_5),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_100),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_75),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_68),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_15),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_69),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_40),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_164),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_27),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_93),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_183),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_179),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_14),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_13),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_181),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_125),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_111),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_101),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_118),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_191),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_155),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_148),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_83),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_182),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_104),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_126),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_63),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_30),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_35),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_129),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_10),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_85),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_67),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_0),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_116),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_23),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_39),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_204),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_134),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_186),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_223),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_176),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_168),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_58),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_219),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_117),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_163),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_112),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_105),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_71),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_77),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_79),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_141),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_76),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_24),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_121),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_75),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_61),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_8),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_120),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_173),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_86),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_71),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_20),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_203),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_81),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_130),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_82),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_137),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_3),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_149),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_68),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_153),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_208),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_113),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_42),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_24),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_212),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_199),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_88),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_85),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_184),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_90),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_6),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_160),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_218),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_177),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_142),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_33),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_139),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_198),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_202),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_215),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_18),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_72),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_23),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_81),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_84),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_154),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_147),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_98),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_73),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_64),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_30),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_96),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_16),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_190),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_48),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_108),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_150),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_9),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_79),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_217),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_17),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_59),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_9),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_80),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_89),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_124),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_77),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_7),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_37),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_67),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_2),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_169),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_66),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_46),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_57),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_143),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_56),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_86),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_3),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_140),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_103),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_26),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_172),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_152),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_11),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_25),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_161),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_52),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_28),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_6),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_1),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_48),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_127),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_166),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_162),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_200),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_88),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_22),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_157),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_38),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_43),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_171),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_72),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_41),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_33),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_110),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_151),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_44),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_205),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_45),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_195),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_158),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_42),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_57),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_7),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_174),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_29),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_180),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_69),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_193),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_102),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_95),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_58),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_13),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_66),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_228),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_229),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_241),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_235),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_241),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_250),
.B(n_0),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_241),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_249),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_241),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_354),
.B(n_2),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_241),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_249),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_236),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_280),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_241),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_328),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_247),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_300),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_351),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_304),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_354),
.B(n_4),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_304),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_252),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_301),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_338),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_256),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_257),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_304),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_304),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_258),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_388),
.B(n_4),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_259),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_321),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_304),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_262),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_304),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_368),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_265),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_10),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_414),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_314),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_314),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_269),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_337),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_250),
.B(n_12),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_321),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_427),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_376),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_250),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_250),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_337),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_270),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_261),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_261),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_261),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_295),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_230),
.B(n_12),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_437),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_273),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_274),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_276),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_249),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_295),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_295),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_376),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_R g515 ( 
.A(n_411),
.B(n_15),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_268),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_281),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_411),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_419),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_246),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_282),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_312),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_289),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_294),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_312),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_297),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_437),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_299),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_302),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_226),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_312),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_418),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_335),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_307),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_335),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_244),
.B(n_17),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_308),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_335),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_392),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_392),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_244),
.B(n_19),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_392),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_407),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_319),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_268),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_266),
.B(n_19),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_330),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_418),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_332),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_334),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_438),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_266),
.B(n_21),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_342),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_345),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_268),
.B(n_21),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_226),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_233),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_233),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_237),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_447),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_493),
.B(n_278),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_451),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_457),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_278),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_497),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_532),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_498),
.B(n_278),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_461),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_467),
.B(n_349),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_539),
.B(n_230),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

CKINVDCx11_ASAP7_75t_R g584 ( 
.A(n_487),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_471),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_453),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_489),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_452),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_455),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_459),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_474),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_498),
.B(n_254),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_464),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_452),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_476),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_446),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_551),
.B(n_357),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_475),
.B(n_246),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_499),
.B(n_254),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_472),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_499),
.B(n_364),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_479),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_448),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_458),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_490),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_462),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_501),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_508),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_509),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_500),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_483),
.B(n_365),
.Y(n_621)
);

AND2x4_ASAP7_75t_SL g622 ( 
.A(n_549),
.B(n_231),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_468),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_473),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_478),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_456),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_517),
.B(n_521),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_523),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_511),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_482),
.B(n_352),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_478),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_524),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_480),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_540),
.B(n_374),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_511),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_526),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_528),
.B(n_378),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_485),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_529),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_486),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_486),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_248),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_534),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_507),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_537),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_527),
.B(n_242),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_488),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_511),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_469),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_545),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_488),
.B(n_364),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_552),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_632),
.A2(n_553),
.B1(n_460),
.B2(n_463),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_652),
.B(n_541),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_652),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_652),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_567),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_565),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_628),
.B(n_583),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_584),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_565),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_572),
.B(n_364),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_568),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_572),
.B(n_543),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_621),
.B(n_254),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_626),
.B(n_450),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_656),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_567),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_572),
.A2(n_450),
.B1(n_465),
.B2(n_454),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_572),
.A2(n_559),
.B1(n_542),
.B2(n_548),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_607),
.A2(n_575),
.B1(n_477),
.B2(n_518),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_570),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_577),
.B(n_557),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_581),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_569),
.Y(n_684)
);

BUFx4f_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_581),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_569),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_571),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_575),
.B(n_543),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_621),
.B(n_254),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_596),
.B(n_254),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_571),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_580),
.B(n_558),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_646),
.B(n_544),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_573),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_573),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_575),
.B(n_372),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_582),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_576),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_574),
.B(n_481),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_589),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_589),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_566),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_606),
.B(n_492),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_646),
.B(n_544),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_600),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_637),
.B(n_547),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_589),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_650),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_587),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_606),
.B(n_492),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_637),
.B(n_547),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_640),
.B(n_495),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_592),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_589),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_578),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_579),
.B(n_519),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_589),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_585),
.B(n_494),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_595),
.B(n_506),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_598),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

XNOR2xp5_ASAP7_75t_L g730 ( 
.A(n_650),
.B(n_484),
.Y(n_730)
);

INVx4_ASAP7_75t_SL g731 ( 
.A(n_596),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_593),
.B(n_495),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_578),
.B(n_550),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_593),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_599),
.B(n_514),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_578),
.B(n_372),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_598),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_596),
.B(n_254),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_598),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_598),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_611),
.B(n_506),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_642),
.A2(n_536),
.B1(n_556),
.B2(n_275),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_594),
.B(n_496),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_614),
.B(n_555),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_594),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_578),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_602),
.B(n_496),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_602),
.B(n_352),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_603),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_620),
.B(n_555),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_656),
.Y(n_751)
);

CKINVDCx16_ASAP7_75t_R g752 ( 
.A(n_620),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_603),
.B(n_426),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_591),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_598),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_610),
.B(n_426),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_617),
.B(n_231),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_604),
.B(n_336),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_605),
.B(n_550),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_605),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_598),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_601),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_656),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_612),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_618),
.B(n_554),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_601),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_591),
.B(n_554),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_624),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_613),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_624),
.B(n_625),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_625),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_610),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_656),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_648),
.B(n_248),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_641),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_SL g777 ( 
.A1(n_615),
.A2(n_344),
.B1(n_377),
.B2(n_263),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_623),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_641),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_643),
.B(n_560),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_643),
.Y(n_781)
);

BUFx10_ASAP7_75t_L g782 ( 
.A(n_619),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_601),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_601),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_645),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_645),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_654),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_629),
.B(n_231),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_610),
.A2(n_239),
.B1(n_243),
.B2(n_237),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_634),
.B(n_560),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_651),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_586),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_601),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_639),
.B(n_530),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_586),
.B(n_502),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_647),
.B(n_231),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_601),
.Y(n_799)
);

AND3x4_ASAP7_75t_L g800 ( 
.A(n_622),
.B(n_515),
.C(n_393),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_586),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_627),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_627),
.B(n_372),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_649),
.B(n_384),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_590),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_627),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_627),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_590),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_622),
.A2(n_405),
.B1(n_429),
.B2(n_380),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_590),
.B(n_502),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_627),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_622),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_597),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_655),
.B(n_563),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_597),
.B(n_516),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_597),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_627),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_685),
.B(n_657),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_682),
.B(n_227),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_797),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_711),
.B(n_271),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_669),
.A2(n_699),
.B1(n_676),
.B2(n_677),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_725),
.B(n_361),
.C(n_346),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_671),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_671),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_768),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_664),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_685),
.B(n_390),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_664),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_711),
.B(n_271),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_764),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_723),
.B(n_358),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_792),
.B(n_346),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_717),
.B(n_277),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_685),
.A2(n_305),
.B1(n_285),
.B2(n_298),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_683),
.B(n_399),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_674),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_681),
.B(n_436),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_669),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_797),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_744),
.B(n_361),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_717),
.B(n_277),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_679),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_683),
.B(n_686),
.Y(n_845)
);

AND2x4_ASAP7_75t_SL g846 ( 
.A(n_681),
.B(n_293),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_796),
.B(n_395),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_679),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_686),
.B(n_400),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_395),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_789),
.B(n_659),
.Y(n_851)
);

INVx8_ASAP7_75t_L g852 ( 
.A(n_669),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_814),
.B(n_403),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_696),
.B(n_561),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_707),
.B(n_285),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_810),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_814),
.B(n_404),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_764),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_742),
.A2(n_243),
.B(n_255),
.C(n_239),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_810),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_764),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_735),
.B(n_404),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_751),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_684),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_716),
.B(n_298),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_756),
.B(n_406),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_718),
.B(n_306),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_684),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_706),
.B(n_768),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_751),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_756),
.B(n_412),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_661),
.B(n_306),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_661),
.B(n_323),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_662),
.B(n_323),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_774),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_681),
.B(n_782),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_756),
.B(n_413),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_669),
.A2(n_324),
.B1(n_348),
.B2(n_341),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_561),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_708),
.B(n_421),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_774),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_669),
.B(n_596),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_662),
.B(n_722),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_777),
.B(n_410),
.C(n_234),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_722),
.B(n_324),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_746),
.B(n_341),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_706),
.B(n_410),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_666),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_746),
.B(n_348),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_678),
.A2(n_439),
.B1(n_440),
.B2(n_431),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_669),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_773),
.B(n_350),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_782),
.B(n_293),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_773),
.B(n_350),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_678),
.A2(n_394),
.B1(n_402),
.B2(n_375),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_671),
.B(n_375),
.Y(n_896)
);

INVx8_ASAP7_75t_L g897 ( 
.A(n_669),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_678),
.A2(n_402),
.B1(n_415),
.B2(n_394),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_688),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_690),
.A2(n_425),
.B(n_428),
.C(n_415),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_771),
.A2(n_638),
.B(n_653),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_702),
.B(n_106),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_708),
.B(n_690),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_688),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_689),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_699),
.A2(n_425),
.B1(n_428),
.B2(n_430),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_690),
.B(n_430),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_776),
.B(n_630),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_708),
.B(n_562),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_689),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_693),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_660),
.B(n_309),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_719),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_693),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_776),
.B(n_630),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_660),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_699),
.A2(n_309),
.B1(n_355),
.B2(n_608),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_666),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_781),
.B(n_630),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_660),
.B(n_727),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_697),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_733),
.B(n_562),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_741),
.B(n_759),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_699),
.A2(n_309),
.B1(n_355),
.B2(n_596),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_697),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_719),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_781),
.B(n_630),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_786),
.B(n_630),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_698),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_786),
.B(n_630),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_793),
.B(n_631),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_733),
.B(n_748),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_665),
.B(n_255),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_733),
.B(n_564),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_721),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_793),
.B(n_631),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_699),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_699),
.A2(n_309),
.B1(n_355),
.B2(n_596),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_668),
.B(n_631),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_809),
.B(n_800),
.C(n_812),
.Y(n_940)
);

BUFx8_ASAP7_75t_L g941 ( 
.A(n_754),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_678),
.A2(n_596),
.B1(n_608),
.B2(n_355),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_698),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_753),
.B(n_309),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_782),
.Y(n_945)
);

INVx8_ASAP7_75t_L g946 ( 
.A(n_699),
.Y(n_946)
);

NAND2x1_ASAP7_75t_L g947 ( 
.A(n_736),
.B(n_596),
.Y(n_947)
);

NOR2x2_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_293),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_765),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_754),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_670),
.B(n_631),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_710),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_715),
.B(n_631),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_675),
.B(n_309),
.Y(n_954)
);

AND2x6_ASAP7_75t_SL g955 ( 
.A(n_775),
.B(n_264),
.Y(n_955)
);

NOR2x1p5_ASAP7_75t_L g956 ( 
.A(n_750),
.B(n_710),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_672),
.A2(n_272),
.B(n_264),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_720),
.B(n_631),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_758),
.B(n_355),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_736),
.A2(n_355),
.B1(n_608),
.B2(n_636),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_SL g961 ( 
.A(n_752),
.B(n_750),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_804),
.B(n_232),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_673),
.A2(n_608),
.B1(n_516),
.B2(n_546),
.Y(n_963)
);

INVx8_ASAP7_75t_L g964 ( 
.A(n_736),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_673),
.B(n_238),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_700),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_700),
.Y(n_967)
);

AOI22x1_ASAP7_75t_L g968 ( 
.A1(n_701),
.A2(n_546),
.B1(n_373),
.B2(n_292),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_766),
.B(n_564),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_701),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_745),
.B(n_609),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_673),
.B(n_503),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_736),
.A2(n_608),
.B1(n_644),
.B2(n_636),
.Y(n_973)
);

NAND2x1_ASAP7_75t_L g974 ( 
.A(n_736),
.B(n_608),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_SL g975 ( 
.A1(n_800),
.A2(n_367),
.B1(n_291),
.B2(n_287),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_709),
.B(n_609),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_798),
.B(n_240),
.Y(n_977)
);

AND2x2_ASAP7_75t_SL g978 ( 
.A(n_672),
.B(n_272),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_709),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_673),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_726),
.B(n_609),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_726),
.B(n_503),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_734),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_783),
.B(n_286),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_703),
.B(n_245),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_665),
.B(n_251),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_734),
.B(n_616),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_749),
.B(n_616),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_665),
.A2(n_608),
.B1(n_546),
.B2(n_296),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_749),
.B(n_616),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_757),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_864),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_854),
.B(n_665),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_952),
.B(n_765),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_840),
.B(n_757),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_864),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_868),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_850),
.B(n_819),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_840),
.B(n_761),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_761),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_SL g1001 ( 
.A(n_891),
.B(n_783),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_831),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_891),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_854),
.Y(n_1004)
);

AND2x6_ASAP7_75t_SL g1005 ( 
.A(n_862),
.B(n_775),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_847),
.B(n_778),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_863),
.B(n_775),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_827),
.B(n_769),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_826),
.B(n_714),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_840),
.B(n_769),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_868),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_904),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_842),
.B(n_857),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_904),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_926),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_905),
.Y(n_1016)
);

OR2x4_ASAP7_75t_L g1017 ( 
.A(n_940),
.B(n_986),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_827),
.B(n_829),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_831),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_829),
.B(n_772),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_879),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_905),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_822),
.B(n_772),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_852),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_926),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_891),
.Y(n_1026)
);

BUFx12f_ASAP7_75t_L g1027 ( 
.A(n_941),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_852),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_844),
.B(n_779),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_910),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_844),
.B(n_779),
.Y(n_1031)
);

INVx8_ASAP7_75t_L g1032 ( 
.A(n_964),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_831),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_869),
.B(n_729),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_945),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_967),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_R g1038 ( 
.A(n_888),
.B(n_770),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_858),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_967),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_952),
.B(n_770),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_863),
.B(n_787),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_941),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_970),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_891),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_970),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_858),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_848),
.B(n_787),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_916),
.B(n_790),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_945),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_820),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_820),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_975),
.B(n_260),
.C(n_253),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_848),
.B(n_790),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_841),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_841),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_984),
.B(n_788),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_913),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_879),
.B(n_791),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_950),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_941),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_949),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_851),
.B(n_788),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_949),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_858),
.B(n_731),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_856),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_909),
.B(n_760),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_899),
.B(n_780),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_882),
.B(n_675),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_899),
.B(n_736),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_888),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_911),
.B(n_736),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_932),
.A2(n_691),
.B1(n_762),
.B2(n_721),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_933),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_861),
.B(n_731),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_911),
.B(n_914),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_914),
.B(n_691),
.Y(n_1079)
);

AO22x1_ASAP7_75t_L g1080 ( 
.A1(n_884),
.A2(n_279),
.B1(n_283),
.B2(n_267),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_903),
.A2(n_915),
.B(n_908),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_860),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_852),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_984),
.B(n_887),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_845),
.B(n_965),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_916),
.B(n_731),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_860),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_918),
.B(n_730),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_861),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_838),
.A2(n_730),
.B1(n_293),
.B2(n_286),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_921),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_SL g1092 ( 
.A(n_985),
.B(n_303),
.C(n_284),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_921),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_972),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_925),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_925),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_861),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_824),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_929),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_923),
.B(n_310),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_909),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_933),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_943),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_943),
.B(n_721),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_966),
.Y(n_1106)
);

AND3x1_ASAP7_75t_SL g1107 ( 
.A(n_956),
.B(n_290),
.C(n_288),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_818),
.B(n_311),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_966),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_979),
.B(n_762),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_979),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_982),
.Y(n_1112)
);

CKINVDCx14_ASAP7_75t_R g1113 ( 
.A(n_918),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_870),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_824),
.B(n_731),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_972),
.B(n_794),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_964),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_969),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_980),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_983),
.B(n_991),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_821),
.B(n_762),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_982),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_870),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_870),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_922),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_825),
.B(n_663),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_881),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_922),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_881),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_980),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_881),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_934),
.Y(n_1132)
);

CKINVDCx11_ASAP7_75t_R g1133 ( 
.A(n_955),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_825),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_830),
.B(n_799),
.Y(n_1135)
);

OA22x2_ASAP7_75t_L g1136 ( 
.A1(n_895),
.A2(n_290),
.B1(n_292),
.B2(n_288),
.Y(n_1136)
);

AND2x6_ASAP7_75t_L g1137 ( 
.A(n_942),
.B(n_663),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_SL g1138 ( 
.A(n_876),
.B(n_313),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_934),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_837),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_969),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_839),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_SL g1143 ( 
.A1(n_933),
.A2(n_389),
.B1(n_318),
.B2(n_326),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_961),
.B(n_799),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_875),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_978),
.A2(n_813),
.B1(n_816),
.B2(n_801),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_976),
.Y(n_1147)
);

AND3x1_ASAP7_75t_SL g1148 ( 
.A(n_948),
.B(n_317),
.C(n_316),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_969),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_962),
.B(n_732),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_834),
.B(n_667),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_981),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_843),
.B(n_883),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_SL g1154 ( 
.A(n_853),
.B(n_327),
.C(n_315),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_933),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_846),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_902),
.B(n_667),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_SL g1158 ( 
.A1(n_893),
.A2(n_329),
.B1(n_333),
.B2(n_339),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_898),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_852),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_964),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_978),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_846),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_987),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_964),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_867),
.B(n_855),
.Y(n_1166)
);

OR2x2_ASAP7_75t_SL g1167 ( 
.A(n_948),
.B(n_316),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_971),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_897),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_865),
.B(n_799),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_920),
.B(n_680),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_897),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_896),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_832),
.B(n_680),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_907),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_866),
.B(n_687),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_885),
.B(n_687),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_886),
.B(n_695),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_988),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_859),
.A2(n_359),
.B(n_331),
.C(n_325),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_871),
.B(n_695),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_954),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_897),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_823),
.B(n_890),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_990),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1013),
.B(n_836),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_998),
.A2(n_1006),
.B1(n_1159),
.B2(n_1015),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1000),
.A2(n_897),
.B1(n_946),
.B2(n_937),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1015),
.Y(n_1189)
);

OA22x2_ASAP7_75t_L g1190 ( 
.A1(n_1025),
.A2(n_977),
.B1(n_989),
.B2(n_959),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1060),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1069),
.B(n_889),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1002),
.B(n_919),
.Y(n_1193)
);

AOI31xp67_ASAP7_75t_L g1194 ( 
.A1(n_1151),
.A2(n_944),
.A3(n_873),
.B(n_874),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1069),
.B(n_892),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1003),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1081),
.A2(n_928),
.B(n_927),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1004),
.B(n_894),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1004),
.B(n_849),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_SL g1200 ( 
.A1(n_1176),
.A2(n_1181),
.B(n_1074),
.Y(n_1200)
);

NAND2x1_ASAP7_75t_L g1201 ( 
.A(n_1024),
.B(n_973),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1153),
.A2(n_946),
.B(n_937),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_931),
.B(n_930),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1021),
.B(n_835),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1151),
.A2(n_936),
.B(n_954),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1073),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1093),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1023),
.A2(n_954),
.B(n_951),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1072),
.A2(n_1166),
.B(n_1079),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1021),
.B(n_872),
.Y(n_1210)
);

INVx3_ASAP7_75t_SL g1211 ( 
.A(n_1163),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1083),
.A2(n_946),
.B(n_937),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1083),
.A2(n_946),
.B(n_937),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1096),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1085),
.A2(n_877),
.B1(n_880),
.B2(n_828),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1083),
.A2(n_1169),
.B(n_1160),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1061),
.A2(n_878),
.B(n_906),
.C(n_963),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1071),
.A2(n_953),
.B(n_939),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1003),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1071),
.A2(n_958),
.B(n_912),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1173),
.B(n_935),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1071),
.A2(n_882),
.B(n_968),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1084),
.B(n_340),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1173),
.B(n_900),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_SL g1225 ( 
.A1(n_1176),
.A2(n_747),
.B(n_743),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1034),
.B(n_347),
.C(n_343),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1061),
.A2(n_917),
.B(n_938),
.C(n_924),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1003),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1083),
.B(n_947),
.Y(n_1229)
);

OAI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1159),
.A2(n_363),
.B1(n_353),
.B2(n_356),
.Y(n_1230)
);

AO32x2_ASAP7_75t_L g1231 ( 
.A1(n_1098),
.A2(n_957),
.A3(n_968),
.B1(n_704),
.B2(n_675),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1036),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1096),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1099),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1018),
.A2(n_974),
.B(n_947),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_995),
.A2(n_712),
.B(n_705),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1065),
.A2(n_974),
.B1(n_957),
.B2(n_785),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1078),
.A2(n_712),
.B(n_705),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1105),
.A2(n_1110),
.B(n_1103),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_724),
.B(n_713),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1083),
.A2(n_763),
.B(n_704),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1180),
.A2(n_805),
.A3(n_794),
.B(n_801),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1002),
.B(n_713),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_1017),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_995),
.A2(n_728),
.B(n_724),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1175),
.B(n_728),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1103),
.A2(n_1104),
.B(n_1010),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1101),
.B(n_737),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1160),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1036),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1115),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1160),
.B(n_704),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_L g1253 ( 
.A1(n_999),
.A2(n_1010),
.B(n_1008),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1122),
.A2(n_1112),
.B(n_1084),
.C(n_1095),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1160),
.A2(n_767),
.B(n_763),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1160),
.A2(n_767),
.B(n_763),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1169),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1122),
.B(n_737),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_999),
.A2(n_740),
.B(n_739),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1094),
.B(n_993),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1168),
.B(n_739),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1104),
.A2(n_1114),
.B(n_1177),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1090),
.B(n_362),
.C(n_360),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1114),
.A2(n_755),
.B(n_740),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1180),
.A2(n_805),
.A3(n_808),
.B(n_816),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1169),
.A2(n_795),
.B(n_767),
.Y(n_1266)
);

NAND2x1_ASAP7_75t_L g1267 ( 
.A(n_1024),
.B(n_755),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1179),
.B(n_784),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1114),
.A2(n_1178),
.B(n_1135),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1121),
.A2(n_785),
.B(n_784),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_992),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1169),
.A2(n_817),
.B(n_795),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1169),
.A2(n_817),
.B(n_795),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1009),
.B(n_371),
.C(n_366),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1116),
.A2(n_901),
.B(n_960),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1073),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1062),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1185),
.B(n_802),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1116),
.B(n_802),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1016),
.A2(n_807),
.B(n_806),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1170),
.A2(n_817),
.B(n_738),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1003),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1022),
.A2(n_807),
.B(n_806),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1009),
.B(n_504),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1044),
.A2(n_811),
.B(n_808),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1020),
.A2(n_811),
.B(n_815),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_993),
.B(n_382),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1125),
.B(n_385),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1029),
.A2(n_441),
.A3(n_320),
.B(n_322),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1044),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1128),
.B(n_387),
.Y(n_1291)
);

NOR4xp25_ASAP7_75t_L g1292 ( 
.A(n_1184),
.B(n_317),
.C(n_416),
.D(n_397),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1123),
.A2(n_505),
.B(n_504),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1132),
.B(n_398),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1101),
.B(n_401),
.Y(n_1295)
);

O2A1O1Ixp5_ASAP7_75t_L g1296 ( 
.A1(n_1108),
.A2(n_442),
.B(n_322),
.C(n_325),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1058),
.B(n_408),
.Y(n_1297)
);

OAI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1100),
.A2(n_417),
.B(n_443),
.Y(n_1298)
);

NOR2x1_ASAP7_75t_SL g1299 ( 
.A(n_1117),
.B(n_320),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1115),
.Y(n_1300)
);

INVx6_ASAP7_75t_SL g1301 ( 
.A(n_1007),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1129),
.A2(n_738),
.B(n_692),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_692),
.B(n_803),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1017),
.A2(n_803),
.B1(n_434),
.B2(n_433),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1139),
.B(n_409),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1051),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1058),
.B(n_1118),
.Y(n_1307)
);

NOR2x1_ASAP7_75t_SL g1308 ( 
.A(n_1117),
.B(n_331),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1050),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_L g1310 ( 
.A(n_1141),
.B(n_107),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1147),
.A2(n_803),
.B(n_633),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1066),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1152),
.A2(n_803),
.B(n_633),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1050),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1031),
.A2(n_442),
.A3(n_369),
.B(n_370),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1152),
.B(n_420),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1164),
.B(n_424),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1164),
.B(n_432),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1048),
.A2(n_441),
.A3(n_369),
.B(n_370),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1003),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1091),
.A2(n_1109),
.B1(n_1111),
.B2(n_1106),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1141),
.B(n_114),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1070),
.B(n_359),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1002),
.B(n_653),
.Y(n_1324)
);

NOR2x1_ASAP7_75t_SL g1325 ( 
.A(n_1117),
.B(n_373),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1131),
.A2(n_638),
.B(n_658),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1052),
.B(n_379),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1055),
.B(n_379),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1024),
.A2(n_644),
.B(n_636),
.Y(n_1329)
);

OAI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1138),
.A2(n_381),
.B(n_383),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1054),
.A2(n_633),
.B(n_635),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1066),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1026),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1049),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1075),
.A2(n_512),
.B(n_513),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_L g1336 ( 
.A1(n_1184),
.A2(n_381),
.B(n_383),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1123),
.A2(n_1127),
.B(n_1124),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1019),
.B(n_653),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1097),
.A2(n_386),
.B(n_391),
.Y(n_1339)
);

AOI211x1_ASAP7_75t_L g1340 ( 
.A1(n_1120),
.A2(n_386),
.B(n_391),
.C(n_396),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1146),
.A2(n_803),
.B(n_644),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1017),
.B(n_22),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1019),
.B(n_653),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1157),
.A2(n_638),
.B(n_658),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1157),
.A2(n_638),
.B(n_658),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1051),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1057),
.B(n_396),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1068),
.B(n_397),
.Y(n_1348)
);

OA22x2_ASAP7_75t_L g1349 ( 
.A1(n_1143),
.A2(n_416),
.B1(n_422),
.B2(n_423),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1124),
.A2(n_531),
.B(n_513),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1186),
.B(n_1064),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1192),
.B(n_1082),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1238),
.A2(n_997),
.B(n_996),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1186),
.A2(n_1215),
.B1(n_1334),
.B2(n_1162),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1336),
.A2(n_1162),
.B1(n_1149),
.B2(n_1102),
.Y(n_1355)
);

BUFx2_ASAP7_75t_SL g1356 ( 
.A(n_1277),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1244),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_SL g1358 ( 
.A1(n_1299),
.A2(n_1059),
.B(n_1140),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1200),
.A2(n_1012),
.B(n_1011),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1285),
.A2(n_1030),
.B(n_1014),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1195),
.B(n_1087),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1206),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1334),
.B(n_1059),
.Y(n_1363)
);

BUFx2_ASAP7_75t_R g1364 ( 
.A(n_1211),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1189),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1233),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1234),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1260),
.B(n_1251),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1204),
.A2(n_1098),
.B1(n_1042),
.B2(n_1150),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1342),
.A2(n_1154),
.B(n_1092),
.C(n_1119),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1297),
.A2(n_1113),
.B1(n_1007),
.B2(n_1001),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1207),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1238),
.A2(n_1037),
.B(n_1035),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1191),
.B(n_1064),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1270),
.A2(n_1174),
.B(n_1046),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1207),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1254),
.B(n_1140),
.Y(n_1377)
);

XNOR2xp5_ASAP7_75t_L g1378 ( 
.A(n_1206),
.B(n_1158),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1209),
.A2(n_1049),
.B(n_1040),
.Y(n_1379)
);

OAI222xp33_ASAP7_75t_L g1380 ( 
.A1(n_1349),
.A2(n_1136),
.B1(n_1102),
.B2(n_1076),
.C1(n_1155),
.C2(n_1142),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1323),
.B(n_1042),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1214),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1223),
.B(n_1042),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1214),
.B(n_1049),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1298),
.A2(n_1149),
.B1(n_1155),
.B2(n_1076),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1297),
.A2(n_1187),
.B1(n_1287),
.B2(n_1295),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1307),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1221),
.A2(n_1134),
.B1(n_1028),
.B2(n_1172),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1202),
.A2(n_1032),
.B(n_1001),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1270),
.A2(n_1127),
.B(n_1157),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1306),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1262),
.A2(n_1181),
.B(n_1176),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1306),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1262),
.A2(n_1181),
.B(n_1077),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1271),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1251),
.B(n_1134),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1263),
.A2(n_1163),
.B1(n_1156),
.B2(n_1063),
.Y(n_1397)
);

AOI21xp33_ASAP7_75t_L g1398 ( 
.A1(n_1226),
.A2(n_1145),
.B(n_1130),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1219),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1346),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1232),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1269),
.A2(n_1077),
.B(n_1067),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1330),
.A2(n_1190),
.B1(n_1342),
.B2(n_1244),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1285),
.A2(n_1033),
.B(n_1019),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1188),
.A2(n_1213),
.B(n_1212),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1271),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1296),
.A2(n_1067),
.B(n_1039),
.C(n_1047),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1254),
.B(n_1033),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1276),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1217),
.A2(n_1171),
.B(n_1097),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1249),
.B(n_1028),
.Y(n_1411)
);

INVx4_ASAP7_75t_SL g1412 ( 
.A(n_1219),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1240),
.A2(n_1039),
.B(n_1033),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1240),
.A2(n_1039),
.B(n_1047),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1216),
.A2(n_1032),
.B(n_1028),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1300),
.B(n_1007),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1280),
.A2(n_1047),
.B(n_1089),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1219),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1249),
.B(n_1172),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1286),
.A2(n_1171),
.B(n_1126),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1312),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1280),
.A2(n_1089),
.B(n_1136),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1219),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1232),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1283),
.A2(n_1089),
.B(n_522),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1290),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1276),
.A2(n_1167),
.B1(n_1113),
.B2(n_1043),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1190),
.A2(n_1171),
.B1(n_1137),
.B2(n_1126),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1321),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1250),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1269),
.A2(n_1239),
.B(n_1197),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1284),
.A2(n_1156),
.B1(n_1063),
.B2(n_1043),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1201),
.A2(n_1032),
.B(n_1172),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1293),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1249),
.A2(n_1032),
.B(n_1165),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1283),
.A2(n_525),
.B(n_533),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1331),
.A2(n_1126),
.B(n_635),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1246),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1228),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1332),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1239),
.A2(n_505),
.B(n_538),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1316),
.B(n_1144),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1199),
.B(n_1005),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1225),
.A2(n_525),
.B(n_533),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1301),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1264),
.A2(n_538),
.B(n_512),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1227),
.A2(n_422),
.B(n_423),
.C(n_444),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1327),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1228),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1317),
.B(n_1053),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1257),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1328),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1244),
.A2(n_1137),
.B1(n_1088),
.B2(n_1041),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_SL g1454 ( 
.A1(n_1227),
.A2(n_444),
.B(n_522),
.C(n_531),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1347),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1224),
.B(n_1167),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1348),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1248),
.B(n_1026),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1250),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1293),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1318),
.B(n_1210),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1258),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1350),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1261),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1279),
.B(n_1026),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1350),
.Y(n_1466)
);

AOI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1288),
.A2(n_1038),
.B(n_1182),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1268),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1278),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1289),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_SL g1471 ( 
.A1(n_1308),
.A2(n_1137),
.B(n_1107),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1337),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1309),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1332),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1248),
.B(n_1026),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1309),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1198),
.B(n_1117),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1289),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1248),
.B(n_1026),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1337),
.Y(n_1480)
);

INVx3_ASAP7_75t_SL g1481 ( 
.A(n_1211),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1264),
.A2(n_535),
.B(n_635),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1217),
.A2(n_1137),
.B(n_1086),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1289),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1292),
.B(n_1045),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1197),
.A2(n_535),
.B(n_1086),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1315),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1274),
.B(n_1080),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1247),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1315),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1314),
.Y(n_1491)
);

O2A1O1Ixp5_ASAP7_75t_SL g1492 ( 
.A1(n_1193),
.A2(n_658),
.B(n_1148),
.C(n_803),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1228),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1275),
.A2(n_1137),
.B(n_1086),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1314),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1282),
.B(n_1117),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1304),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1236),
.A2(n_1137),
.B(n_1183),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1245),
.A2(n_1183),
.B(n_1165),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1315),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1315),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1230),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1247),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1203),
.A2(n_1115),
.B(n_803),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1291),
.B(n_1045),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1301),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1294),
.B(n_1133),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1228),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1301),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1319),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1333),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1305),
.B(n_1133),
.C(n_1045),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1259),
.A2(n_1183),
.B(n_1165),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1282),
.B(n_1045),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1319),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1335),
.A2(n_994),
.B(n_1182),
.Y(n_1516)
);

BUFx2_ASAP7_75t_SL g1517 ( 
.A(n_1333),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1333),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1319),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1319),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1349),
.B(n_1045),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1282),
.B(n_1161),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1310),
.A2(n_1027),
.B1(n_1165),
.B2(n_1161),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1242),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1401),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1366),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_R g1528 ( 
.A(n_1362),
.B(n_1027),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1497),
.A2(n_1339),
.B1(n_1322),
.B2(n_1193),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1367),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1416),
.B(n_1196),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1356),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_L g1534 ( 
.A(n_1403),
.B(n_1340),
.C(n_1237),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1456),
.B(n_1324),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1497),
.A2(n_1335),
.B1(n_1343),
.B2(n_1338),
.Y(n_1536)
);

AO21x1_ASAP7_75t_L g1537 ( 
.A1(n_1369),
.A2(n_1253),
.B(n_1243),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1361),
.B(n_1320),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1351),
.B(n_1325),
.Y(n_1539)
);

AO31x2_ASAP7_75t_L g1540 ( 
.A1(n_1470),
.A2(n_1281),
.A3(n_1231),
.B(n_1302),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1456),
.B(n_1387),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1494),
.A2(n_1311),
.B(n_1313),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1355),
.A2(n_1333),
.B1(n_1056),
.B2(n_1196),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1416),
.B(n_1401),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1352),
.A2(n_1056),
.B1(n_1303),
.B2(n_1341),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1352),
.B(n_1242),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1354),
.A2(n_1343),
.B1(n_1338),
.B2(n_1324),
.C(n_1243),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1443),
.A2(n_1208),
.B1(n_1205),
.B2(n_1220),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1430),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1386),
.A2(n_1056),
.B1(n_1161),
.B2(n_1183),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1430),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1444),
.A2(n_1205),
.B(n_1218),
.Y(n_1552)
);

CKINVDCx16_ASAP7_75t_R g1553 ( 
.A(n_1427),
.Y(n_1553)
);

OAI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1502),
.A2(n_1345),
.B1(n_1344),
.B2(n_1329),
.C(n_1326),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1481),
.Y(n_1555)
);

NAND3x1_ASAP7_75t_L g1556 ( 
.A(n_1507),
.B(n_25),
.C(n_26),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1410),
.A2(n_1208),
.B(n_1194),
.Y(n_1557)
);

NAND2xp33_ASAP7_75t_R g1558 ( 
.A(n_1362),
.B(n_1235),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1476),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1426),
.Y(n_1560)
);

OAI21xp33_ASAP7_75t_L g1561 ( 
.A1(n_1461),
.A2(n_1220),
.B(n_1218),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1440),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1409),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1476),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1488),
.A2(n_1056),
.B1(n_1257),
.B2(n_1165),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1387),
.B(n_1242),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1368),
.B(n_1242),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1416),
.B(n_1056),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_R g1569 ( 
.A(n_1409),
.B(n_1161),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1365),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1475),
.Y(n_1571)
);

NAND2xp33_ASAP7_75t_R g1572 ( 
.A(n_1506),
.B(n_1235),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1442),
.B(n_115),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1364),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1450),
.A2(n_1257),
.B1(n_1161),
.B2(n_1183),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1370),
.A2(n_1267),
.B(n_1229),
.C(n_1272),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1448),
.A2(n_1222),
.B(n_1266),
.C(n_1256),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1491),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1452),
.A2(n_1222),
.B1(n_1229),
.B2(n_1255),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1357),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1506),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1455),
.B(n_1252),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1491),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1368),
.B(n_1265),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1399),
.Y(n_1585)
);

OAI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1371),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1363),
.B(n_1265),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1492),
.A2(n_1273),
.B(n_1241),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1453),
.A2(n_1252),
.B1(n_1231),
.B2(n_1265),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1372),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_1357),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1412),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1475),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1438),
.B(n_1265),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1363),
.B(n_31),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1428),
.A2(n_1483),
.B1(n_1457),
.B2(n_1381),
.Y(n_1596)
);

OR2x6_ASAP7_75t_L g1597 ( 
.A(n_1433),
.B(n_1231),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1368),
.B(n_1231),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1445),
.B(n_119),
.Y(n_1599)
);

AND2x6_ASAP7_75t_L g1600 ( 
.A(n_1485),
.B(n_122),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1383),
.B(n_31),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1385),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_1602)
);

INVx6_ASAP7_75t_L g1603 ( 
.A(n_1412),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1376),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1512),
.A2(n_608),
.B1(n_34),
.B2(n_37),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1464),
.B(n_32),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1468),
.B(n_38),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1395),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1374),
.B(n_41),
.Y(n_1609)
);

INVx5_ASAP7_75t_L g1610 ( 
.A(n_1399),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1485),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1447),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.C(n_52),
.Y(n_1612)
);

AND2x6_ASAP7_75t_L g1613 ( 
.A(n_1521),
.B(n_222),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1471),
.B(n_1377),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1471),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1377),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1469),
.B(n_55),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1429),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1405),
.A2(n_638),
.B(n_221),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1382),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_R g1621 ( 
.A(n_1445),
.B(n_220),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1474),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1521),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1444),
.A2(n_211),
.B(n_209),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1424),
.Y(n_1625)
);

BUFx8_ASAP7_75t_L g1626 ( 
.A(n_1509),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1475),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1391),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1478),
.A2(n_207),
.B(n_206),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1399),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1398),
.A2(n_1505),
.B1(n_1467),
.B2(n_1378),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1395),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1447),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.C(n_70),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1432),
.A2(n_638),
.B1(n_70),
.B2(n_73),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1406),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_SL g1636 ( 
.A1(n_1523),
.A2(n_65),
.B(n_74),
.C(n_76),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1479),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1436),
.A2(n_123),
.B(n_192),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1462),
.B(n_74),
.Y(n_1639)
);

AND2x2_ASAP7_75t_SL g1640 ( 
.A(n_1408),
.B(n_78),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1458),
.B(n_82),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1384),
.B(n_83),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1473),
.A2(n_84),
.B1(n_87),
.B2(n_90),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1397),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1505),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1378),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1458),
.B(n_97),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1481),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1393),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1421),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1509),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1384),
.B(n_99),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1408),
.A2(n_100),
.B1(n_135),
.B2(n_136),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1436),
.A2(n_144),
.B(n_145),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1459),
.A2(n_1493),
.B1(n_1501),
.B2(n_1520),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1459),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1479),
.B(n_146),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1465),
.B(n_196),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1400),
.B(n_159),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1465),
.B(n_189),
.Y(n_1660)
);

CKINVDCx6p67_ASAP7_75t_R g1661 ( 
.A(n_1517),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1379),
.A2(n_167),
.B(n_170),
.C(n_178),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1396),
.B(n_185),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1396),
.B(n_187),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1446),
.A2(n_188),
.B(n_1482),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1389),
.A2(n_1504),
.B(n_1454),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_R g1667 ( 
.A(n_1479),
.B(n_1518),
.Y(n_1667)
);

INVx8_ASAP7_75t_L g1668 ( 
.A(n_1514),
.Y(n_1668)
);

AOI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1420),
.A2(n_1437),
.B(n_1519),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1396),
.B(n_1388),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1454),
.B(n_1477),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1518),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1359),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1514),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1399),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1359),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_SL g1677 ( 
.A(n_1451),
.B(n_1435),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1484),
.B(n_1500),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1477),
.A2(n_1516),
.B1(n_1358),
.B2(n_1487),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1490),
.B(n_1510),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1514),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1380),
.A2(n_1515),
.B1(n_1358),
.B2(n_1524),
.C(n_1407),
.Y(n_1682)
);

BUFx12f_ASAP7_75t_L g1683 ( 
.A(n_1399),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1360),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1412),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1516),
.A2(n_1394),
.B1(n_1402),
.B2(n_1392),
.Y(n_1686)
);

OAI222xp33_ASAP7_75t_L g1687 ( 
.A1(n_1420),
.A2(n_1419),
.B1(n_1411),
.B2(n_1451),
.C1(n_1522),
.C2(n_1496),
.Y(n_1687)
);

INVx6_ASAP7_75t_L g1688 ( 
.A(n_1412),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1360),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1492),
.B(n_1522),
.C(n_1496),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1422),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1422),
.Y(n_1692)
);

NAND2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1418),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1516),
.B(n_1418),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1418),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1434),
.A2(n_1466),
.B1(n_1463),
.B2(n_1460),
.C(n_1353),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1418),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1423),
.B(n_1439),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1423),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1394),
.Y(n_1701)
);

AO31x2_ASAP7_75t_L g1702 ( 
.A1(n_1434),
.A2(n_1460),
.A3(n_1463),
.B(n_1466),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1394),
.B(n_1402),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1423),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1402),
.A2(n_1392),
.B1(n_1423),
.B2(n_1449),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1392),
.B(n_1439),
.Y(n_1706)
);

BUFx2_ASAP7_75t_SL g1707 ( 
.A(n_1439),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1646),
.A2(n_1489),
.B1(n_1503),
.B2(n_1431),
.C(n_1415),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1526),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1603),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1541),
.B(n_1439),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1640),
.A2(n_1489),
.B1(n_1503),
.B2(n_1353),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1602),
.A2(n_1480),
.B1(n_1472),
.B2(n_1375),
.C(n_1508),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1612),
.A2(n_1353),
.B1(n_1373),
.B2(n_1472),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1644),
.A2(n_1431),
.B1(n_1419),
.B2(n_1411),
.C(n_1486),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1631),
.A2(n_1411),
.B1(n_1419),
.B2(n_1508),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1564),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1612),
.A2(n_1373),
.B1(n_1480),
.B2(n_1486),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1641),
.B(n_1439),
.Y(n_1719)
);

AO21x2_ASAP7_75t_L g1720 ( 
.A1(n_1666),
.A2(n_1588),
.B(n_1557),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1535),
.B(n_1566),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1647),
.B(n_1449),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1633),
.A2(n_1373),
.B1(n_1486),
.B2(n_1375),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1602),
.A2(n_1375),
.B1(n_1511),
.B2(n_1508),
.C(n_1449),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1595),
.B(n_1441),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1530),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1555),
.Y(n_1727)
);

AOI222xp33_ASAP7_75t_L g1728 ( 
.A1(n_1633),
.A2(n_1511),
.B1(n_1449),
.B2(n_1508),
.C1(n_1404),
.C2(n_1498),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1618),
.A2(n_1441),
.B1(n_1390),
.B2(n_1431),
.Y(n_1729)
);

OR2x6_ASAP7_75t_L g1730 ( 
.A(n_1614),
.B(n_1498),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1666),
.A2(n_1425),
.B(n_1446),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1618),
.A2(n_1441),
.B1(n_1390),
.B2(n_1449),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1539),
.A2(n_1511),
.B1(n_1508),
.B2(n_1390),
.Y(n_1733)
);

OAI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1651),
.A2(n_1437),
.B(n_1482),
.C(n_1404),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1616),
.A2(n_1413),
.B1(n_1414),
.B2(n_1417),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1526),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1621),
.A2(n_1413),
.B1(n_1414),
.B2(n_1417),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1683),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1616),
.A2(n_1425),
.B1(n_1499),
.B2(n_1513),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1586),
.A2(n_1611),
.B1(n_1645),
.B2(n_1636),
.C(n_1534),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1529),
.A2(n_1499),
.B1(n_1513),
.B2(n_1556),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1586),
.B(n_1634),
.C(n_1643),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_SL g1743 ( 
.A1(n_1600),
.A2(n_1653),
.B1(n_1613),
.B2(n_1550),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1533),
.A2(n_1622),
.B1(n_1562),
.B2(n_1553),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1562),
.A2(n_1622),
.B1(n_1531),
.B2(n_1525),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1542),
.A2(n_1545),
.B(n_1619),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1600),
.A2(n_1653),
.B1(n_1613),
.B2(n_1550),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1531),
.A2(n_1536),
.B1(n_1625),
.B2(n_1685),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1544),
.B(n_1601),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1609),
.A2(n_1573),
.B(n_1662),
.C(n_1596),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1623),
.A2(n_1600),
.B1(n_1605),
.B2(n_1615),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1600),
.A2(n_1596),
.B1(n_1613),
.B2(n_1607),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1606),
.A2(n_1607),
.B1(n_1617),
.B2(n_1667),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1600),
.A2(n_1613),
.B1(n_1617),
.B2(n_1606),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1603),
.Y(n_1755)
);

AND2x4_ASAP7_75t_SL g1756 ( 
.A(n_1551),
.B(n_1583),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1563),
.Y(n_1757)
);

OAI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1554),
.A2(n_1639),
.B1(n_1619),
.B2(n_1652),
.C(n_1642),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1554),
.A2(n_1639),
.B1(n_1652),
.B2(n_1642),
.C(n_1650),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1544),
.B(n_1571),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1706),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1625),
.A2(n_1565),
.B1(n_1614),
.B2(n_1570),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1538),
.A2(n_1558),
.B1(n_1545),
.B2(n_1591),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1613),
.A2(n_1599),
.B1(n_1655),
.B2(n_1580),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1587),
.B(n_1546),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1706),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1599),
.A2(n_1648),
.B1(n_1542),
.B2(n_1560),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1687),
.A2(n_1577),
.B(n_1561),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1626),
.A2(n_1657),
.B1(n_1670),
.B2(n_1660),
.Y(n_1769)
);

OR2x2_ASAP7_75t_SL g1770 ( 
.A(n_1526),
.B(n_1559),
.Y(n_1770)
);

AO31x2_ASAP7_75t_L g1771 ( 
.A1(n_1537),
.A2(n_1589),
.A3(n_1676),
.B(n_1673),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1574),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1614),
.B(n_1695),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_1626),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1590),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1575),
.A2(n_1656),
.B1(n_1578),
.B2(n_1583),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1593),
.B(n_1627),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1548),
.A2(n_1658),
.B1(n_1660),
.B2(n_1582),
.C(n_1547),
.Y(n_1778)
);

AOI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1677),
.A2(n_1669),
.B(n_1671),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1546),
.B(n_1567),
.Y(n_1780)
);

NOR4xp25_ASAP7_75t_L g1781 ( 
.A(n_1589),
.B(n_1658),
.C(n_1594),
.D(n_1679),
.Y(n_1781)
);

AOI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1576),
.A2(n_1572),
.B(n_1594),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_SL g1783 ( 
.A(n_1549),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1687),
.A2(n_1557),
.B(n_1576),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1657),
.A2(n_1581),
.B1(n_1547),
.B2(n_1584),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1551),
.A2(n_1543),
.B1(n_1661),
.B2(n_1627),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1664),
.A2(n_1528),
.B1(n_1543),
.B2(n_1579),
.C(n_1659),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1637),
.A2(n_1559),
.B1(n_1688),
.B2(n_1603),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1637),
.B(n_1672),
.Y(n_1789)
);

AOI321xp33_ASAP7_75t_L g1790 ( 
.A1(n_1682),
.A2(n_1671),
.A3(n_1628),
.B1(n_1649),
.B2(n_1620),
.C(n_1604),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1682),
.A2(n_1686),
.B(n_1705),
.C(n_1629),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1663),
.A2(n_1559),
.B1(n_1629),
.B2(n_1532),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1688),
.A2(n_1681),
.B1(n_1674),
.B2(n_1675),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1697),
.A2(n_1690),
.B1(n_1678),
.B2(n_1680),
.C(n_1692),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1598),
.B(n_1635),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1592),
.A2(n_1638),
.B(n_1654),
.Y(n_1796)
);

BUFx6f_ASAP7_75t_L g1797 ( 
.A(n_1688),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1532),
.A2(n_1690),
.B(n_1568),
.Y(n_1798)
);

AO222x2_ASAP7_75t_L g1799 ( 
.A1(n_1568),
.A2(n_1699),
.B1(n_1569),
.B2(n_1668),
.C1(n_1608),
.C2(n_1632),
.Y(n_1799)
);

NAND2x1_ASAP7_75t_L g1800 ( 
.A(n_1592),
.B(n_1696),
.Y(n_1800)
);

AO31x2_ASAP7_75t_L g1801 ( 
.A1(n_1684),
.A2(n_1689),
.A3(n_1703),
.B(n_1701),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1697),
.A2(n_1691),
.B1(n_1588),
.B2(n_1703),
.C(n_1700),
.Y(n_1802)
);

BUFx4f_ASAP7_75t_SL g1803 ( 
.A(n_1585),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1693),
.A2(n_1668),
.B1(n_1610),
.B2(n_1630),
.Y(n_1804)
);

OAI211xp5_ASAP7_75t_L g1805 ( 
.A1(n_1704),
.A2(n_1668),
.B(n_1624),
.C(n_1698),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1585),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1597),
.A2(n_1624),
.B1(n_1585),
.B2(n_1694),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1693),
.A2(n_1630),
.B1(n_1610),
.B2(n_1694),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1694),
.B(n_1707),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_SL g1810 ( 
.A(n_1597),
.B(n_1610),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1610),
.A2(n_1630),
.B1(n_1540),
.B2(n_1597),
.C(n_1702),
.Y(n_1811)
);

OAI211xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1540),
.A2(n_1552),
.B(n_1702),
.C(n_1665),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1552),
.B(n_1641),
.Y(n_1813)
);

OAI211xp5_ASAP7_75t_L g1814 ( 
.A1(n_1646),
.A2(n_1013),
.B(n_850),
.C(n_998),
.Y(n_1814)
);

INVx2_ASAP7_75t_SL g1815 ( 
.A(n_1526),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1527),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1602),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.C(n_632),
.Y(n_1817)
);

OAI21xp33_ASAP7_75t_L g1818 ( 
.A1(n_1644),
.A2(n_1013),
.B(n_998),
.Y(n_1818)
);

INVx8_ASAP7_75t_L g1819 ( 
.A(n_1668),
.Y(n_1819)
);

OAI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1646),
.A2(n_1013),
.B(n_850),
.C(n_998),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1667),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1640),
.A2(n_838),
.B1(n_1013),
.B2(n_893),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1541),
.B(n_1438),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1562),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1526),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1644),
.A2(n_998),
.B1(n_1013),
.B2(n_838),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1526),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1646),
.A2(n_1013),
.B1(n_998),
.B2(n_1090),
.C(n_850),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1541),
.B(n_1438),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1541),
.B(n_1535),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1833)
);

OAI211xp5_ASAP7_75t_L g1834 ( 
.A1(n_1646),
.A2(n_1013),
.B(n_850),
.C(n_998),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1564),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1836)
);

OAI21xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1612),
.A2(n_1633),
.B(n_1640),
.Y(n_1837)
);

INVx4_ASAP7_75t_SL g1838 ( 
.A(n_1600),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1644),
.A2(n_998),
.B1(n_1013),
.B2(n_838),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1640),
.A2(n_838),
.B1(n_1013),
.B2(n_893),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1542),
.A2(n_998),
.B(n_1494),
.Y(n_1841)
);

OAI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1646),
.A2(n_1013),
.B(n_850),
.C(n_998),
.Y(n_1842)
);

CKINVDCx16_ASAP7_75t_R g1843 ( 
.A(n_1528),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1646),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.C(n_1090),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1641),
.B(n_1647),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1644),
.A2(n_998),
.B1(n_1013),
.B2(n_838),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1849)
);

NOR2xp67_ASAP7_75t_L g1850 ( 
.A(n_1533),
.B(n_1512),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1631),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1853)
);

OAI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1644),
.A2(n_998),
.B1(n_1013),
.B2(n_838),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1640),
.A2(n_838),
.B1(n_1013),
.B2(n_893),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1541),
.B(n_1438),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_SL g1857 ( 
.A1(n_1640),
.A2(n_838),
.B1(n_1013),
.B2(n_893),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1602),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.C(n_632),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1631),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1586),
.A2(n_1013),
.B(n_850),
.C(n_998),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_998),
.B2(n_850),
.Y(n_1862)
);

OA21x2_ASAP7_75t_L g1863 ( 
.A1(n_1666),
.A2(n_1557),
.B(n_1682),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1564),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1765),
.B(n_1761),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1773),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1863),
.B(n_1813),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1863),
.B(n_1720),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1761),
.B(n_1766),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1730),
.B(n_1810),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1730),
.B(n_1773),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1730),
.B(n_1773),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1863),
.B(n_1720),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1838),
.B(n_1801),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1771),
.B(n_1801),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1771),
.B(n_1801),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1775),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1780),
.B(n_1753),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1753),
.B(n_1805),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1771),
.B(n_1781),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1770),
.Y(n_1881)
);

AO31x2_ASAP7_75t_L g1882 ( 
.A1(n_1746),
.A2(n_1784),
.A3(n_1768),
.B(n_1841),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1721),
.B(n_1802),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1833),
.A2(n_1853),
.B1(n_1862),
.B2(n_1852),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1726),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1811),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1816),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1821),
.B(n_1832),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1795),
.B(n_1725),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1794),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1779),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1833),
.A2(n_1849),
.B1(n_1846),
.B2(n_1836),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1838),
.B(n_1807),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1712),
.B(n_1735),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1712),
.B(n_1735),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1731),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1762),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1824),
.B(n_1831),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1752),
.B(n_1782),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1711),
.B(n_1791),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1731),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1731),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1752),
.B(n_1729),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1708),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1851),
.A2(n_1860),
.B1(n_1817),
.B2(n_1858),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1729),
.B(n_1732),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1732),
.B(n_1743),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1799),
.B(n_1837),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1739),
.B(n_1728),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1733),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1812),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1737),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1713),
.B(n_1723),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1737),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1758),
.Y(n_1916)
);

OAI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1742),
.A2(n_1845),
.B1(n_1827),
.B2(n_1839),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1717),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1835),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1856),
.B(n_1763),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1759),
.B(n_1827),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1714),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1724),
.B(n_1718),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1790),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1718),
.B(n_1754),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1777),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1800),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1763),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1778),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1798),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1822),
.B(n_1836),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1715),
.Y(n_1932)
);

AND2x4_ASAP7_75t_SL g1933 ( 
.A(n_1767),
.B(n_1792),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1754),
.B(n_1838),
.Y(n_1934)
);

OAI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1846),
.A2(n_1853),
.B(n_1862),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1825),
.B(n_1864),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1719),
.B(n_1722),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1748),
.B(n_1741),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1776),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1829),
.B(n_1847),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1844),
.B(n_1785),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1796),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1839),
.B(n_1848),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1786),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1785),
.B(n_1792),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1808),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1849),
.B(n_1852),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1760),
.B(n_1749),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1767),
.B(n_1789),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1745),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1859),
.B(n_1861),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1888),
.B(n_1859),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1869),
.Y(n_1953)
);

OAI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1896),
.A2(n_1716),
.B(n_1769),
.Y(n_1954)
);

AOI33xp33_ASAP7_75t_L g1955 ( 
.A1(n_1905),
.A2(n_1857),
.A3(n_1855),
.B1(n_1823),
.B2(n_1840),
.B3(n_1854),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1888),
.B(n_1744),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1917),
.A2(n_1818),
.B(n_1848),
.Y(n_1957)
);

AOI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1917),
.A2(n_1830),
.B1(n_1854),
.B2(n_1834),
.C(n_1842),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1877),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1877),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1896),
.A2(n_1769),
.B(n_1804),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1869),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1867),
.B(n_1937),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1865),
.B(n_1815),
.Y(n_1964)
);

OAI211xp5_ASAP7_75t_L g1965 ( 
.A1(n_1905),
.A2(n_1820),
.B(n_1814),
.C(n_1740),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1936),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1874),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1867),
.B(n_1809),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1921),
.A2(n_1750),
.B1(n_1751),
.B2(n_1764),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1898),
.B(n_1850),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1887),
.Y(n_1971)
);

BUFx8_ASAP7_75t_L g1972 ( 
.A(n_1946),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1936),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1921),
.A2(n_1787),
.B(n_1793),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1887),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1867),
.B(n_1709),
.Y(n_1976)
);

NAND4xp25_ASAP7_75t_L g1977 ( 
.A(n_1951),
.B(n_1751),
.C(n_1828),
.D(n_1826),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1929),
.B(n_1843),
.Y(n_1978)
);

INVx4_ASAP7_75t_L g1979 ( 
.A(n_1927),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1943),
.A2(n_1783),
.B1(n_1727),
.B2(n_1774),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1898),
.B(n_1709),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1926),
.B(n_1828),
.Y(n_1982)
);

AOI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1884),
.A2(n_1783),
.B1(n_1788),
.B2(n_1734),
.C(n_1736),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_L g1984 ( 
.A(n_1943),
.B(n_1710),
.C(n_1755),
.Y(n_1984)
);

AOI33xp33_ASAP7_75t_L g1985 ( 
.A1(n_1924),
.A2(n_1756),
.A3(n_1736),
.B1(n_1757),
.B2(n_1772),
.B3(n_1803),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1909),
.A2(n_1819),
.B1(n_1738),
.B2(n_1755),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1926),
.B(n_1806),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1936),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1870),
.B(n_1819),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1909),
.A2(n_1738),
.B1(n_1710),
.B2(n_1755),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1879),
.A2(n_1756),
.B(n_1803),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1865),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1890),
.A2(n_1819),
.B1(n_1710),
.B2(n_1797),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1874),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1874),
.Y(n_1995)
);

OA21x2_ASAP7_75t_L g1996 ( 
.A1(n_1901),
.A2(n_1902),
.B(n_1942),
.Y(n_1996)
);

OAI33xp33_ASAP7_75t_L g1997 ( 
.A1(n_1884),
.A2(n_1797),
.A3(n_1892),
.B1(n_1924),
.B2(n_1951),
.B3(n_1929),
.Y(n_1997)
);

NAND3xp33_ASAP7_75t_L g1998 ( 
.A(n_1879),
.B(n_1797),
.C(n_1890),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1892),
.A2(n_1890),
.B1(n_1935),
.B2(n_1947),
.C(n_1932),
.Y(n_1999)
);

CKINVDCx16_ASAP7_75t_R g2000 ( 
.A(n_1881),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1935),
.B(n_1916),
.C(n_1932),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1947),
.A2(n_1938),
.B1(n_1946),
.B2(n_1916),
.Y(n_2002)
);

AO21x2_ASAP7_75t_L g2003 ( 
.A1(n_1901),
.A2(n_1902),
.B(n_1880),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1950),
.B(n_1919),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1918),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1919),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1874),
.Y(n_2007)
);

AO21x2_ASAP7_75t_L g2008 ( 
.A1(n_1901),
.A2(n_1902),
.B(n_1880),
.Y(n_2008)
);

O2A1O1Ixp5_ASAP7_75t_L g2009 ( 
.A1(n_1916),
.A2(n_1899),
.B(n_1910),
.C(n_1908),
.Y(n_2009)
);

AOI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1886),
.A2(n_1880),
.B1(n_1899),
.B2(n_1910),
.C(n_1950),
.Y(n_2010)
);

INVxp67_ASAP7_75t_SL g2011 ( 
.A(n_1891),
.Y(n_2011)
);

OR2x6_ASAP7_75t_L g2012 ( 
.A(n_1870),
.B(n_1871),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1914),
.A2(n_1923),
.B(n_1904),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1865),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1948),
.B(n_1931),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1891),
.Y(n_2016)
);

OAI221xp5_ASAP7_75t_L g2017 ( 
.A1(n_1886),
.A2(n_1920),
.B1(n_1938),
.B2(n_1899),
.C(n_1931),
.Y(n_2017)
);

INVx2_ASAP7_75t_SL g2018 ( 
.A(n_1918),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1926),
.B(n_1878),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1995),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1996),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1963),
.B(n_1967),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1998),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1958),
.A2(n_1908),
.B1(n_1907),
.B2(n_1910),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1996),
.Y(n_2025)
);

AND2x4_ASAP7_75t_SL g2026 ( 
.A(n_1989),
.B(n_1893),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1959),
.Y(n_2027)
);

OAI21xp5_ASAP7_75t_SL g2028 ( 
.A1(n_1965),
.A2(n_1908),
.B(n_1907),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1959),
.Y(n_2029)
);

NAND4xp25_ASAP7_75t_SL g2030 ( 
.A(n_2010),
.B(n_1907),
.C(n_1930),
.D(n_1878),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1992),
.B(n_1913),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1960),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1960),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_2003),
.B(n_1882),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1969),
.A2(n_1938),
.B1(n_1923),
.B2(n_1897),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_2014),
.B(n_1913),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1979),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1953),
.B(n_1886),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1971),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1967),
.B(n_1868),
.Y(n_2040)
);

OAI21x1_ASAP7_75t_L g2041 ( 
.A1(n_1961),
.A2(n_1996),
.B(n_1954),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1972),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_2003),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_2003),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1994),
.B(n_1868),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_2012),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2007),
.B(n_1873),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2008),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2007),
.B(n_1873),
.Y(n_2049)
);

NOR2x1_ASAP7_75t_L g2050 ( 
.A(n_1979),
.B(n_1912),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1972),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1962),
.B(n_2019),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2013),
.B(n_1920),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1970),
.B(n_1948),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2011),
.B(n_1912),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1966),
.B(n_1915),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2016),
.B(n_1885),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_2008),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2008),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1999),
.B(n_1930),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1995),
.B(n_1915),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1973),
.B(n_1885),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1995),
.B(n_1875),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_1988),
.B(n_1889),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_1957),
.A2(n_1914),
.B(n_1923),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1968),
.B(n_1875),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1968),
.B(n_1875),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1976),
.B(n_1876),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2015),
.B(n_1883),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1975),
.B(n_1883),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1976),
.B(n_1876),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1956),
.B(n_1948),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2073)
);

INVx2_ASAP7_75t_SL g2074 ( 
.A(n_2042),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2038),
.B(n_1964),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_2030),
.A2(n_2017),
.B1(n_1925),
.B2(n_2001),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2027),
.Y(n_2077)
);

BUFx2_ASAP7_75t_SL g2078 ( 
.A(n_2042),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2038),
.B(n_1964),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2023),
.B(n_2004),
.Y(n_2080)
);

OAI211xp5_ASAP7_75t_L g2081 ( 
.A1(n_2028),
.A2(n_1974),
.B(n_1977),
.C(n_1983),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2022),
.B(n_2012),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_2023),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2056),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2069),
.B(n_2006),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2027),
.Y(n_2087)
);

BUFx2_ASAP7_75t_SL g2088 ( 
.A(n_2042),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2029),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2029),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2032),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2021),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2032),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2070),
.B(n_1882),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_2051),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2069),
.B(n_1952),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2046),
.B(n_2000),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_2046),
.B(n_1870),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2052),
.B(n_1981),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2033),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2070),
.B(n_1882),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2066),
.B(n_1989),
.Y(n_2102)
);

AOI322xp5_ASAP7_75t_L g2103 ( 
.A1(n_2024),
.A2(n_2060),
.A3(n_2053),
.B1(n_2028),
.B2(n_1980),
.C1(n_1978),
.C2(n_1914),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2066),
.B(n_1989),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_2051),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2066),
.B(n_1989),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2052),
.B(n_1883),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_2050),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2056),
.B(n_2031),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_2055),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2021),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2067),
.B(n_1870),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2065),
.B(n_1897),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2033),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2031),
.B(n_1882),
.Y(n_2115)
);

AOI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2030),
.A2(n_1997),
.B1(n_1925),
.B2(n_2002),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2051),
.B(n_1972),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2064),
.Y(n_2118)
);

AOI33xp33_ASAP7_75t_L g2119 ( 
.A1(n_2061),
.A2(n_1903),
.A3(n_1925),
.B1(n_1895),
.B2(n_1894),
.B3(n_1940),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2039),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2021),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2067),
.B(n_1870),
.Y(n_2122)
);

OAI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2065),
.A2(n_1955),
.B(n_2035),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2072),
.B(n_2054),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2039),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2109),
.B(n_2055),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2121),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2117),
.B(n_2035),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_2109),
.B(n_2036),
.Y(n_2129)
);

INVxp67_ASAP7_75t_L g2130 ( 
.A(n_2078),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2123),
.A2(n_1903),
.B1(n_1945),
.B2(n_1934),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2077),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2077),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2102),
.B(n_2067),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_2103),
.B(n_2009),
.Y(n_2135)
);

NAND2xp33_ASAP7_75t_SL g2136 ( 
.A(n_2076),
.B(n_1985),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_2103),
.A2(n_1974),
.B(n_2050),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2102),
.B(n_2063),
.Y(n_2138)
);

NOR2x1p5_ASAP7_75t_L g2139 ( 
.A(n_2084),
.B(n_1881),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2104),
.B(n_2063),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2113),
.B(n_2062),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2104),
.B(n_2063),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2080),
.B(n_2062),
.Y(n_2143)
);

A2O1A1Ixp33_ASAP7_75t_L g2144 ( 
.A1(n_2123),
.A2(n_1991),
.B(n_1933),
.C(n_2041),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2096),
.B(n_2068),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2106),
.B(n_2068),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2119),
.B(n_2068),
.Y(n_2147)
);

A2O1A1Ixp33_ASAP7_75t_SL g2148 ( 
.A1(n_2081),
.A2(n_1928),
.B(n_1927),
.C(n_1986),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2110),
.B(n_2107),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2078),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2106),
.B(n_2071),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2098),
.B(n_2026),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2116),
.B(n_2071),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2116),
.B(n_2071),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2121),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2073),
.B(n_2040),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2118),
.B(n_2036),
.Y(n_2157)
);

NAND4xp25_ASAP7_75t_L g2158 ( 
.A(n_2094),
.B(n_2034),
.C(n_1928),
.D(n_1903),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2124),
.B(n_2057),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_SL g2160 ( 
.A(n_2086),
.B(n_1990),
.C(n_2005),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2121),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2087),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2099),
.B(n_2074),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2085),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2087),
.Y(n_2165)
);

NOR3xp33_ASAP7_75t_SL g2166 ( 
.A(n_2088),
.B(n_2005),
.C(n_1984),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2073),
.B(n_2082),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2115),
.B(n_2064),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2089),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2082),
.B(n_2040),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2089),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2083),
.B(n_2040),
.Y(n_2172)
);

INVx3_ASAP7_75t_SL g2173 ( 
.A(n_2074),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2115),
.B(n_2057),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2090),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2121),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2083),
.B(n_2045),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2108),
.Y(n_2178)
);

NAND2xp33_ASAP7_75t_SL g2179 ( 
.A(n_2097),
.B(n_1940),
.Y(n_2179)
);

OAI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2135),
.A2(n_2097),
.B(n_2108),
.Y(n_2180)
);

AOI222xp33_ASAP7_75t_L g2181 ( 
.A1(n_2136),
.A2(n_1895),
.B1(n_1894),
.B2(n_1906),
.C1(n_1945),
.C2(n_1941),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2131),
.B(n_2095),
.Y(n_2182)
);

AOI21xp33_ASAP7_75t_L g2183 ( 
.A1(n_2148),
.A2(n_2105),
.B(n_2095),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2126),
.B(n_2094),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2159),
.B(n_2105),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2139),
.B(n_2088),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2137),
.A2(n_2026),
.B1(n_1881),
.B2(n_1939),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2132),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_2137),
.A2(n_2144),
.B(n_2160),
.Y(n_2189)
);

AOI21xp33_ASAP7_75t_L g2190 ( 
.A1(n_2150),
.A2(n_2101),
.B(n_2034),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2143),
.B(n_2075),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2126),
.B(n_2101),
.Y(n_2192)
);

NOR3xp33_ASAP7_75t_L g2193 ( 
.A(n_2130),
.B(n_1961),
.C(n_2041),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2132),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2133),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2139),
.B(n_2098),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2179),
.A2(n_2098),
.B1(n_1871),
.B2(n_1872),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2133),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2162),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2128),
.A2(n_2041),
.B(n_1954),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2150),
.B(n_2075),
.Y(n_2201)
);

NAND4xp25_ASAP7_75t_L g2202 ( 
.A(n_2153),
.B(n_1993),
.C(n_1900),
.D(n_2034),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2129),
.B(n_2079),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2164),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2167),
.B(n_2146),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2162),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2167),
.B(n_2098),
.Y(n_2207)
);

OAI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2154),
.A2(n_1939),
.B1(n_1944),
.B2(n_2079),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2173),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2163),
.B(n_2061),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2127),
.Y(n_2211)
);

INVx1_ASAP7_75t_SL g2212 ( 
.A(n_2173),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2147),
.B(n_2061),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2166),
.A2(n_2026),
.B1(n_1944),
.B2(n_1871),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2141),
.A2(n_1933),
.B(n_1945),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_2173),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2152),
.A2(n_1871),
.B1(n_1872),
.B2(n_1893),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2158),
.A2(n_1933),
.B(n_1982),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2157),
.A2(n_2018),
.B(n_1900),
.Y(n_2219)
);

OAI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2180),
.A2(n_2158),
.B1(n_2178),
.B2(n_1900),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2209),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2181),
.B(n_2204),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2205),
.B(n_2146),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2212),
.B(n_2216),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2209),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2205),
.B(n_2151),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2182),
.B(n_2151),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2191),
.B(n_2149),
.Y(n_2228)
);

OAI21xp33_ASAP7_75t_L g2229 ( 
.A1(n_2189),
.A2(n_2174),
.B(n_2157),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2201),
.B(n_2134),
.Y(n_2230)
);

OAI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2202),
.A2(n_2178),
.B1(n_1904),
.B2(n_1911),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2206),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2201),
.B(n_2134),
.Y(n_2233)
);

AOI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2187),
.A2(n_2152),
.B1(n_2172),
.B2(n_2170),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2196),
.B(n_2152),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2206),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2185),
.B(n_2152),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2188),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2186),
.A2(n_2177),
.B1(n_2172),
.B2(n_2170),
.Y(n_2239)
);

NAND3xp33_ASAP7_75t_L g2240 ( 
.A(n_2183),
.B(n_2174),
.C(n_2169),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2186),
.Y(n_2241)
);

OAI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2200),
.A2(n_2129),
.B1(n_2168),
.B2(n_2175),
.C(n_2171),
.Y(n_2242)
);

OAI21xp33_ASAP7_75t_L g2243 ( 
.A1(n_2213),
.A2(n_2168),
.B(n_2156),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_SL g2244 ( 
.A1(n_2214),
.A2(n_2175),
.B(n_2171),
.Y(n_2244)
);

OAI21xp33_ASAP7_75t_L g2245 ( 
.A1(n_2203),
.A2(n_2177),
.B(n_2156),
.Y(n_2245)
);

XNOR2x1_ASAP7_75t_L g2246 ( 
.A(n_2208),
.B(n_1940),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_2215),
.A2(n_1895),
.B1(n_1894),
.B2(n_1904),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2218),
.B(n_2207),
.Y(n_2248)
);

AOI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2220),
.A2(n_2190),
.B1(n_2219),
.B2(n_2193),
.C(n_2198),
.Y(n_2249)
);

INVxp67_ASAP7_75t_L g2250 ( 
.A(n_2241),
.Y(n_2250)
);

XOR2xp5_ASAP7_75t_L g2251 ( 
.A(n_2224),
.B(n_2217),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2241),
.Y(n_2252)
);

NOR3xp33_ASAP7_75t_SL g2253 ( 
.A(n_2222),
.B(n_2194),
.C(n_2195),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2221),
.B(n_2207),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2221),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2235),
.B(n_2196),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2232),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2225),
.B(n_2203),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2236),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2238),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2230),
.B(n_2199),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2225),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2220),
.B(n_2197),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2233),
.Y(n_2264)
);

AOI21xp33_ASAP7_75t_L g2265 ( 
.A1(n_2240),
.A2(n_2184),
.B(n_2192),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2223),
.B(n_2226),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2228),
.Y(n_2267)
);

AOI31xp33_ASAP7_75t_L g2268 ( 
.A1(n_2247),
.A2(n_2192),
.A3(n_2184),
.B(n_2210),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_SL g2269 ( 
.A(n_2229),
.B(n_2145),
.C(n_2169),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_2248),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2239),
.B(n_2138),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2246),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2262),
.Y(n_2273)
);

AOI211xp5_ASAP7_75t_L g2274 ( 
.A1(n_2265),
.A2(n_2231),
.B(n_2244),
.C(n_2242),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_2255),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_2250),
.Y(n_2276)
);

NAND4xp25_ASAP7_75t_L g2277 ( 
.A(n_2264),
.B(n_2270),
.C(n_2267),
.D(n_2258),
.Y(n_2277)
);

NOR4xp25_ASAP7_75t_L g2278 ( 
.A(n_2270),
.B(n_2231),
.C(n_2245),
.D(n_2243),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2256),
.B(n_2237),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2262),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2269),
.A2(n_2247),
.B(n_2234),
.C(n_2237),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2255),
.Y(n_2282)
);

A2O1A1Ixp33_ASAP7_75t_L g2283 ( 
.A1(n_2253),
.A2(n_2227),
.B(n_2246),
.C(n_2165),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2272),
.A2(n_2142),
.B1(n_2138),
.B2(n_2140),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2252),
.B(n_2140),
.Y(n_2285)
);

NAND5xp2_ASAP7_75t_L g2286 ( 
.A(n_2267),
.B(n_1934),
.C(n_1941),
.D(n_2142),
.E(n_2165),
.Y(n_2286)
);

AOI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2274),
.A2(n_2251),
.B(n_2263),
.Y(n_2287)
);

AOI221xp5_ASAP7_75t_L g2288 ( 
.A1(n_2278),
.A2(n_2249),
.B1(n_2272),
.B2(n_2268),
.C(n_2251),
.Y(n_2288)
);

OAI211xp5_ASAP7_75t_SL g2289 ( 
.A1(n_2281),
.A2(n_2254),
.B(n_2261),
.C(n_2260),
.Y(n_2289)
);

OAI211xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2283),
.A2(n_2261),
.B(n_2260),
.C(n_2257),
.Y(n_2290)
);

AOI211xp5_ASAP7_75t_L g2291 ( 
.A1(n_2283),
.A2(n_2256),
.B(n_2271),
.C(n_2266),
.Y(n_2291)
);

AOI321xp33_ASAP7_75t_L g2292 ( 
.A1(n_2279),
.A2(n_2271),
.A3(n_2266),
.B1(n_2259),
.B2(n_2257),
.C(n_2211),
.Y(n_2292)
);

AOI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2277),
.A2(n_2259),
.B1(n_2211),
.B2(n_2176),
.C(n_2161),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2276),
.A2(n_2058),
.B1(n_2161),
.B2(n_2155),
.C1(n_2127),
.C2(n_2176),
.Y(n_2294)
);

OAI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2285),
.A2(n_2176),
.B1(n_2161),
.B2(n_2155),
.C(n_2127),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2286),
.A2(n_2155),
.B1(n_2058),
.B2(n_2111),
.C(n_2092),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_R g2297 ( 
.A(n_2275),
.B(n_1934),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_R g2298 ( 
.A(n_2297),
.B(n_2275),
.Y(n_2298)
);

INVx3_ASAP7_75t_SL g2299 ( 
.A(n_2292),
.Y(n_2299)
);

AOI21xp33_ASAP7_75t_SL g2300 ( 
.A1(n_2294),
.A2(n_2282),
.B(n_2280),
.Y(n_2300)
);

NOR2x1_ASAP7_75t_L g2301 ( 
.A(n_2290),
.B(n_2273),
.Y(n_2301)
);

NAND2xp33_ASAP7_75t_SL g2302 ( 
.A(n_2291),
.B(n_2282),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2288),
.A2(n_2284),
.B1(n_2020),
.B2(n_2037),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2287),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2289),
.A2(n_1941),
.B(n_1893),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2301),
.B(n_2092),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2298),
.Y(n_2307)
);

INVxp33_ASAP7_75t_L g2308 ( 
.A(n_2303),
.Y(n_2308)
);

NAND4xp75_ASAP7_75t_L g2309 ( 
.A(n_2299),
.B(n_2293),
.C(n_2296),
.D(n_2295),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2304),
.B(n_2112),
.Y(n_2310)
);

NOR3x1_ASAP7_75t_L g2311 ( 
.A(n_2305),
.B(n_2020),
.C(n_2018),
.Y(n_2311)
);

NOR3xp33_ASAP7_75t_L g2312 ( 
.A(n_2302),
.B(n_2037),
.C(n_2111),
.Y(n_2312)
);

NOR2xp67_ASAP7_75t_SL g2313 ( 
.A(n_2300),
.B(n_1918),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2313),
.B(n_2090),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2310),
.Y(n_2315)
);

NAND3xp33_ASAP7_75t_L g2316 ( 
.A(n_2312),
.B(n_2111),
.C(n_2037),
.Y(n_2316)
);

NAND5xp2_ASAP7_75t_L g2317 ( 
.A(n_2308),
.B(n_1949),
.C(n_2112),
.D(n_2122),
.E(n_2049),
.Y(n_2317)
);

NOR3xp33_ASAP7_75t_L g2318 ( 
.A(n_2307),
.B(n_2037),
.C(n_1987),
.Y(n_2318)
);

OAI321xp33_ASAP7_75t_L g2319 ( 
.A1(n_2309),
.A2(n_2020),
.A3(n_2122),
.B1(n_1866),
.B2(n_1942),
.C(n_1922),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2315),
.Y(n_2320)
);

OR2x6_ASAP7_75t_L g2321 ( 
.A(n_2314),
.B(n_2306),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2316),
.Y(n_2322)
);

OAI221xp5_ASAP7_75t_R g2323 ( 
.A1(n_2318),
.A2(n_2311),
.B1(n_2306),
.B2(n_2125),
.C(n_2120),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2321),
.B(n_2319),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2321),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2325),
.A2(n_2320),
.B1(n_2322),
.B2(n_2324),
.Y(n_2326)
);

AOI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2326),
.A2(n_2323),
.B1(n_2317),
.B2(n_2125),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2326),
.B(n_2120),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2328),
.B(n_2091),
.Y(n_2329)
);

OAI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2327),
.A2(n_2114),
.B1(n_2100),
.B2(n_2093),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2330),
.A2(n_2114),
.B1(n_2100),
.B2(n_2093),
.Y(n_2331)
);

AOI322xp5_ASAP7_75t_L g2332 ( 
.A1(n_2331),
.A2(n_2329),
.A3(n_2025),
.B1(n_2091),
.B2(n_2047),
.C1(n_2049),
.C2(n_2045),
.Y(n_2332)
);

OAI221xp5_ASAP7_75t_R g2333 ( 
.A1(n_2332),
.A2(n_2048),
.B1(n_2044),
.B2(n_2043),
.C(n_2059),
.Y(n_2333)
);

AOI211xp5_ASAP7_75t_L g2334 ( 
.A1(n_2333),
.A2(n_2043),
.B(n_2048),
.C(n_2044),
.Y(n_2334)
);


endmodule