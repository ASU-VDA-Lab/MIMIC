module fake_jpeg_9015_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_25),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_27),
.C(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_48),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_33),
.B1(n_32),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_64),
.B1(n_68),
.B2(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_59),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_33),
.B1(n_31),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_42),
.B1(n_32),
.B2(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_23),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_33),
.B1(n_32),
.B2(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_33),
.B1(n_42),
.B2(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_27),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_27),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_40),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_53),
.C(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_22),
.B1(n_30),
.B2(n_23),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_17),
.B(n_16),
.C(n_24),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_61),
.B(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_49),
.B1(n_47),
.B2(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_95),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_46),
.B1(n_56),
.B2(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_23),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_44),
.B1(n_47),
.B2(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_109),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_107),
.B1(n_103),
.B2(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_104),
.C(n_89),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_21),
.B(n_53),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_97),
.CI(n_92),
.CON(n_145),
.SN(n_145)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_87),
.C(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_22),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_1),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_120),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_97),
.B(n_75),
.Y(n_149)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_121),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_60),
.B1(n_57),
.B2(n_26),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_117),
.B1(n_123),
.B2(n_24),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_67),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_145),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_95),
.C(n_91),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_146),
.C(n_102),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_86),
.B1(n_122),
.B2(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_89),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_160),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_124),
.A3(n_110),
.B1(n_115),
.B2(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_165),
.B(n_168),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_108),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_177),
.C(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_175),
.B(n_180),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_93),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_152),
.B1(n_148),
.B2(n_137),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_116),
.A3(n_119),
.B1(n_106),
.B2(n_90),
.C1(n_93),
.C2(n_82),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_183),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_129),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_150),
.B(n_138),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_187),
.B(n_195),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_149),
.B1(n_131),
.B2(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_154),
.B1(n_168),
.B2(n_164),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_128),
.B1(n_137),
.B2(n_149),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_194),
.B1(n_196),
.B2(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_199),
.C(n_203),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_149),
.B1(n_126),
.B2(n_127),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_151),
.B(n_145),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_130),
.B(n_145),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_132),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_134),
.C(n_141),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_141),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_134),
.C(n_82),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_163),
.C(n_155),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_216),
.B(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_219),
.C(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_188),
.C(n_203),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_171),
.C(n_154),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_75),
.C(n_169),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_153),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_200),
.B1(n_191),
.B2(n_174),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_159),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_166),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_8),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_158),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_202),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_234),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_196),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_240),
.C(n_248),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_224),
.B(n_231),
.C(n_209),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_192),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_211),
.CI(n_223),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_192),
.B1(n_193),
.B2(n_187),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_249),
.B1(n_245),
.B2(n_254),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_252),
.B1(n_214),
.B2(n_227),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_16),
.C(n_17),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_169),
.B1(n_113),
.B2(n_90),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_222),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_262),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_268),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_212),
.B(n_215),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_16),
.B(n_28),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_220),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_242),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.C(n_272),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_235),
.C(n_240),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_88),
.B1(n_72),
.B2(n_74),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_74),
.B1(n_67),
.B2(n_46),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_21),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_251),
.C(n_248),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_281),
.C(n_285),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_234),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_9),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_233),
.C(n_241),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_14),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_286),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_276),
.B(n_269),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_264),
.B1(n_260),
.B2(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_74),
.C(n_56),
.Y(n_285)
);

OAI322xp33_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_17),
.A3(n_28),
.B1(n_24),
.B2(n_12),
.C1(n_5),
.C2(n_6),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_11),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_12),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_308)
);

AOI31xp67_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_8),
.A3(n_15),
.B(n_14),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_266),
.CI(n_261),
.CON(n_291),
.SN(n_291)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_300),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_278),
.B1(n_273),
.B2(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_297),
.C(n_298),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_267),
.B1(n_271),
.B2(n_28),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_11),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_11),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_9),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_274),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_8),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_293),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_56),
.A3(n_50),
.B1(n_62),
.B2(n_7),
.C1(n_6),
.C2(n_13),
.Y(n_309)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_310),
.B(n_7),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_50),
.A3(n_62),
.B1(n_7),
.B2(n_15),
.C1(n_3),
.C2(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_295),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_317),
.B(n_307),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_316),
.B(n_1),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_62),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_15),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_324)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_303),
.B(n_2),
.Y(n_321)
);

AOI321xp33_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_316),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_3),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_324),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_3),
.Y(n_328)
);


endmodule