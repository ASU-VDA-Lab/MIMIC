module real_jpeg_15037_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_275, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_275;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_48),
.B1(n_63),
.B2(n_66),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_48),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_3),
.A2(n_32),
.B1(n_34),
.B2(n_48),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_63),
.C(n_78),
.Y(n_144)
);

NAND2x1_ASAP7_75t_SL g148 ( 
.A(n_6),
.B(n_35),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_67),
.B(n_155),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_31),
.B(n_34),
.C(n_182),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_6),
.A2(n_32),
.B1(n_34),
.B2(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_46),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_32),
.B1(n_34),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_8),
.A2(n_43),
.B1(n_63),
.B2(n_66),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_101),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_63),
.B1(n_66),
.B2(n_101),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_32),
.B1(n_34),
.B2(n_101),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_32),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_12),
.A2(n_40),
.B1(n_63),
.B2(n_66),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_32),
.B1(n_34),
.B2(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_14),
.A2(n_57),
.B1(n_63),
.B2(n_66),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_63),
.B1(n_66),
.B2(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_15),
.A2(n_32),
.B1(n_34),
.B2(n_82),
.Y(n_113)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

XNOR2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.C(n_93),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_22),
.A2(n_23),
.B1(n_85),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_84),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_44),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_26),
.B(n_44),
.C(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_27),
.A2(n_41),
.B1(n_42),
.B2(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_27),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_27),
.A2(n_41),
.B1(n_201),
.B2(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_27),
.A2(n_188),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_104),
.Y(n_103)
);

NOR2x1_ASAP7_75t_R g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_30),
.A2(n_36),
.B(n_140),
.Y(n_182)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_32),
.B(n_51),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_34),
.A2(n_47),
.A3(n_52),
.B1(n_225),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_35),
.B(n_104),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_36),
.A2(n_37),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_37),
.B(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_39),
.A2(n_41),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_41),
.A2(n_103),
.B(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_54),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_49),
.B(n_140),
.C(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_50),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_50),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_50),
.A2(n_100),
.B(n_122),
.Y(n_249)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_55),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_59),
.A2(n_73),
.B1(n_74),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_68),
.B1(n_69),
.B2(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_66),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_66),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_67),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_67),
.A2(n_72),
.B1(n_184),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_67),
.A2(n_72),
.B1(n_208),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_69),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_68),
.A2(n_69),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_68),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_69),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_72),
.A2(n_161),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_72),
.B(n_140),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_72),
.A2(n_169),
.B(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_81),
.B2(n_83),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_76),
.B1(n_83),
.B2(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_81),
.B1(n_83),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_76),
.B(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_76),
.A2(n_83),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_91),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_80),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_80),
.B(n_140),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_80),
.A2(n_152),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_85),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_87),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_92),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_93),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_102),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_94),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_95),
.B(n_97),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_96),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_98),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_99),
.B(n_102),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_127),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_115),
.B2(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_114),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_112),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_110),
.A2(n_141),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_126),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_268),
.B(n_273),
.Y(n_129)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_242),
.A3(n_261),
.B1(n_266),
.B2(n_267),
.C(n_275),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_217),
.B(n_241),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_195),
.B(n_216),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_177),
.B(n_194),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_157),
.B(n_176),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_153),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_165),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_170),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_189),
.C(n_193),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_183),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_209),
.B2(n_210),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_212),
.C(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_203),
.C(n_207),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_232),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_233),
.C(n_234),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_231),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_227),
.C(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_254),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_254),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.C(n_253),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_245),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_251),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_253),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.C(n_260),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_272),
.Y(n_273)
);


endmodule