module real_aes_830_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_835, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_836, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_835;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_836;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g569 ( .A(n_0), .B(n_201), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_1), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g136 ( .A(n_2), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_3), .B(n_548), .Y(n_585) );
NAND2xp33_ASAP7_75t_SL g625 ( .A(n_4), .B(n_157), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_5), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g618 ( .A(n_6), .Y(n_618) );
INVx1_ASAP7_75t_L g168 ( .A(n_7), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_8), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_9), .Y(n_183) );
AND2x2_ASAP7_75t_L g583 ( .A(n_10), .B(n_160), .Y(n_583) );
INVx2_ASAP7_75t_L g128 ( .A(n_11), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_12), .Y(n_490) );
INVx1_ASAP7_75t_L g202 ( .A(n_13), .Y(n_202) );
AOI221x1_ASAP7_75t_L g621 ( .A1(n_14), .A2(n_125), .B1(n_550), .B2(n_622), .C(n_624), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_15), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g494 ( .A(n_16), .Y(n_494) );
INVx1_ASAP7_75t_L g199 ( .A(n_17), .Y(n_199) );
INVx1_ASAP7_75t_SL g253 ( .A(n_18), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_19), .B(n_151), .Y(n_215) );
AOI33xp33_ASAP7_75t_L g239 ( .A1(n_20), .A2(n_53), .A3(n_133), .B1(n_144), .B2(n_240), .B3(n_241), .Y(n_239) );
AOI221xp5_ASAP7_75t_SL g559 ( .A1(n_21), .A2(n_44), .B1(n_548), .B2(n_550), .C(n_560), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_22), .A2(n_550), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_23), .B(n_201), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_24), .A2(n_38), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_24), .Y(n_109) );
INVx1_ASAP7_75t_L g176 ( .A(n_25), .Y(n_176) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_26), .A2(n_91), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g161 ( .A(n_26), .B(n_91), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_27), .B(n_204), .Y(n_553) );
INVxp67_ASAP7_75t_L g620 ( .A(n_28), .Y(n_620) );
AND2x2_ASAP7_75t_L g607 ( .A(n_29), .B(n_159), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_30), .B(n_131), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_31), .A2(n_550), .B(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_32), .Y(n_498) );
OAI22x1_ASAP7_75t_R g111 ( .A1(n_33), .A2(n_37), .B1(n_112), .B2(n_113), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_33), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_33), .B(n_471), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_34), .B(n_204), .Y(n_561) );
AND2x2_ASAP7_75t_L g138 ( .A(n_35), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g143 ( .A(n_35), .Y(n_143) );
AND2x2_ASAP7_75t_L g157 ( .A(n_35), .B(n_136), .Y(n_157) );
OR2x6_ASAP7_75t_L g492 ( .A(n_36), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_37), .Y(n_112) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_38), .A2(n_104), .B1(n_502), .B2(n_507), .C(n_516), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_38), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_39), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_40), .B(n_131), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_41), .A2(n_126), .B1(n_193), .B2(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_42), .B(n_217), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_43), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_43), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_45), .B(n_151), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_46), .A2(n_83), .B1(n_141), .B2(n_550), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_47), .B(n_201), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_48), .B(n_165), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_49), .B(n_151), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_50), .Y(n_212) );
AND2x2_ASAP7_75t_L g572 ( .A(n_51), .B(n_159), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_52), .B(n_159), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_54), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g134 ( .A(n_55), .Y(n_134) );
INVx1_ASAP7_75t_L g153 ( .A(n_55), .Y(n_153) );
AND2x2_ASAP7_75t_L g158 ( .A(n_56), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_57), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g166 ( .A1(n_58), .A2(n_76), .B1(n_131), .B2(n_141), .C(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_59), .B(n_131), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_60), .B(n_548), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_61), .B(n_126), .Y(n_185) );
AOI21xp5_ASAP7_75t_SL g223 ( .A1(n_62), .A2(n_141), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g598 ( .A(n_63), .B(n_159), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_64), .B(n_204), .Y(n_570) );
INVx1_ASAP7_75t_L g196 ( .A(n_65), .Y(n_196) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_66), .B(n_160), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_67), .B(n_201), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_68), .A2(n_550), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g148 ( .A(n_69), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_70), .B(n_204), .Y(n_589) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_71), .B(n_165), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_72), .A2(n_141), .B(n_147), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g523 ( .A1(n_73), .A2(n_95), .B1(n_524), .B2(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_73), .Y(n_524) );
INVx1_ASAP7_75t_L g139 ( .A(n_74), .Y(n_139) );
INVx1_ASAP7_75t_L g155 ( .A(n_74), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_75), .B(n_131), .Y(n_242) );
AND2x2_ASAP7_75t_L g255 ( .A(n_77), .B(n_125), .Y(n_255) );
INVx1_ASAP7_75t_L g197 ( .A(n_78), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_79), .A2(n_141), .B(n_252), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_80), .A2(n_141), .B(n_214), .C(n_218), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_81), .A2(n_86), .B1(n_131), .B2(n_548), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_82), .B(n_548), .Y(n_597) );
INVx1_ASAP7_75t_L g495 ( .A(n_84), .Y(n_495) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_85), .B(n_125), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_87), .A2(n_141), .B1(n_237), .B2(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_88), .B(n_201), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_89), .B(n_201), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_90), .A2(n_550), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g225 ( .A(n_92), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_93), .B(n_204), .Y(n_595) );
AND2x2_ASAP7_75t_L g243 ( .A(n_94), .B(n_125), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_95), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_96), .A2(n_174), .B(n_175), .C(n_178), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_97), .B(n_548), .Y(n_571) );
INVxp67_ASAP7_75t_L g623 ( .A(n_98), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_99), .B(n_204), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_100), .A2(n_550), .B(n_551), .Y(n_549) );
BUFx2_ASAP7_75t_L g506 ( .A(n_101), .Y(n_506) );
BUFx2_ASAP7_75t_SL g513 ( .A(n_101), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_102), .B(n_151), .Y(n_226) );
OAI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_487), .B(n_496), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B1(n_485), .B2(n_486), .Y(n_106) );
INVx1_ASAP7_75t_L g486 ( .A(n_107), .Y(n_486) );
INVx2_ASAP7_75t_L g485 ( .A(n_110), .Y(n_485) );
XNOR2x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_113), .A2(n_358), .B(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_113), .A2(n_116), .B1(n_403), .B2(n_835), .Y(n_535) );
NAND4xp75_ASAP7_75t_L g114 ( .A(n_115), .B(n_357), .C(n_402), .D(n_471), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR4xp25_ASAP7_75t_L g530 ( .A(n_116), .B(n_358), .C(n_403), .D(n_531), .Y(n_530) );
NAND2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_317), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_273), .C(n_298), .Y(n_117) );
OAI222xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_187), .B1(n_228), .B2(n_244), .C1(n_260), .C2(n_267), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_162), .Y(n_120) );
AND2x2_ASAP7_75t_L g482 ( .A(n_121), .B(n_296), .Y(n_482) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_123), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_123), .B(n_171), .Y(n_272) );
INVx3_ASAP7_75t_L g287 ( .A(n_123), .Y(n_287) );
AND2x2_ASAP7_75t_L g420 ( .A(n_123), .B(n_421), .Y(n_420) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_129), .B(n_158), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_124), .A2(n_125), .B1(n_173), .B2(n_179), .Y(n_172) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_124), .A2(n_129), .B(n_158), .Y(n_305) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_126), .B(n_182), .Y(n_181) );
AOI21x1_ASAP7_75t_L g565 ( .A1(n_126), .A2(n_566), .B(n_572), .Y(n_565) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_128), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g193 ( .A(n_128), .B(n_161), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_140), .Y(n_129) );
INVx1_ASAP7_75t_L g186 ( .A(n_131), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_131), .A2(n_141), .B1(n_617), .B2(n_619), .Y(n_616) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
INVx1_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
OR2x6_ASAP7_75t_L g149 ( .A(n_133), .B(n_145), .Y(n_149) );
INVxp33_ASAP7_75t_L g240 ( .A(n_133), .Y(n_240) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g146 ( .A(n_134), .B(n_136), .Y(n_146) );
AND2x4_ASAP7_75t_L g204 ( .A(n_134), .B(n_154), .Y(n_204) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g550 ( .A(n_138), .B(n_146), .Y(n_550) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
AND2x6_ASAP7_75t_L g201 ( .A(n_139), .B(n_152), .Y(n_201) );
INVxp67_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NOR2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g241 ( .A(n_144), .Y(n_241) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_150), .C(n_156), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_149), .A2(n_156), .B(n_168), .C(n_169), .Y(n_167) );
INVxp67_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_177), .B1(n_196), .B2(n_197), .Y(n_195) );
INVx2_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_149), .A2(n_156), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_149), .A2(n_156), .B(n_253), .C(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
AND2x4_ASAP7_75t_L g548 ( .A(n_151), .B(n_157), .Y(n_548) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_156), .B(n_193), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_156), .A2(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g237 ( .A(n_156), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_156), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_156), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_156), .A2(n_569), .B(n_570), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_156), .A2(n_588), .B(n_589), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_156), .A2(n_595), .B(n_596), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_156), .A2(n_604), .B(n_605), .Y(n_603) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_159), .Y(n_248) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_159), .A2(n_559), .B(n_563), .Y(n_558) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g350 ( .A(n_162), .B(n_303), .Y(n_350) );
AND2x2_ASAP7_75t_L g352 ( .A(n_162), .B(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g387 ( .A(n_162), .Y(n_387) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_171), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVxp67_ASAP7_75t_L g270 ( .A(n_164), .Y(n_270) );
INVx1_ASAP7_75t_L g289 ( .A(n_164), .Y(n_289) );
AND2x4_ASAP7_75t_L g296 ( .A(n_164), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_164), .B(n_234), .Y(n_312) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_164), .Y(n_421) );
INVx1_ASAP7_75t_L g431 ( .A(n_164), .Y(n_431) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
INVx2_ASAP7_75t_SL g218 ( .A(n_165), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_165), .A2(n_547), .B(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
INVx2_ASAP7_75t_L g284 ( .A(n_171), .Y(n_284) );
INVx1_ASAP7_75t_L g365 ( .A(n_171), .Y(n_365) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_180), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_177), .B(n_193), .C(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_189), .B(n_219), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_189), .B(n_246), .Y(n_340) );
INVx2_ASAP7_75t_L g361 ( .A(n_189), .Y(n_361) );
AND2x2_ASAP7_75t_L g369 ( .A(n_189), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_206), .Y(n_189) );
AND2x4_ASAP7_75t_L g259 ( .A(n_190), .B(n_207), .Y(n_259) );
INVx1_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
AND2x2_ASAP7_75t_L g442 ( .A(n_190), .B(n_247), .Y(n_442) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g280 ( .A(n_191), .B(n_207), .Y(n_280) );
INVx2_ASAP7_75t_L g316 ( .A(n_191), .Y(n_316) );
AND2x2_ASAP7_75t_L g395 ( .A(n_191), .B(n_247), .Y(n_395) );
NOR2x1_ASAP7_75t_SL g438 ( .A(n_191), .B(n_220), .Y(n_438) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_194), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_193), .A2(n_223), .B(n_227), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_193), .A2(n_585), .B(n_586), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_193), .B(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_193), .B(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_193), .B(n_623), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_198), .B(n_205), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B1(n_202), .B2(n_203), .Y(n_198) );
INVxp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g278 ( .A(n_206), .Y(n_278) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g292 ( .A(n_207), .B(n_220), .Y(n_292) );
INVx1_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_207), .Y(n_416) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_213), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .C(n_212), .Y(n_209) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_218), .A2(n_235), .B(n_243), .Y(n_234) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_218), .A2(n_235), .B(n_243), .Y(n_285) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_218), .A2(n_577), .B(n_580), .Y(n_576) );
AND2x2_ASAP7_75t_L g279 ( .A(n_219), .B(n_280), .Y(n_279) );
OR2x6_ASAP7_75t_L g360 ( .A(n_219), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g398 ( .A(n_219), .B(n_395), .Y(n_398) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx4_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_220), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g327 ( .A(n_220), .Y(n_327) );
OR2x2_ASAP7_75t_L g333 ( .A(n_220), .B(n_247), .Y(n_333) );
AND2x4_ASAP7_75t_L g347 ( .A(n_220), .B(n_308), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_220), .B(n_316), .Y(n_348) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g392 ( .A(n_231), .B(n_311), .Y(n_392) );
BUFx2_ASAP7_75t_L g444 ( .A(n_231), .Y(n_444) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g475 ( .A(n_233), .B(n_387), .Y(n_475) );
INVx2_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_242), .Y(n_235) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_256), .Y(n_244) );
AND2x2_ASAP7_75t_L g291 ( .A(n_245), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x4_ASAP7_75t_SL g276 ( .A(n_246), .B(n_266), .Y(n_276) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g264 ( .A(n_247), .Y(n_264) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_247), .Y(n_370) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_247), .Y(n_437) );
INVx1_ASAP7_75t_L g477 ( .A(n_247), .Y(n_477) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_255), .Y(n_247) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_248), .A2(n_592), .B(n_598), .Y(n_591) );
AO21x2_ASAP7_75t_L g600 ( .A1(n_248), .A2(n_601), .B(n_607), .Y(n_600) );
AO21x2_ASAP7_75t_L g645 ( .A1(n_248), .A2(n_601), .B(n_607), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
BUFx2_ASAP7_75t_L g391 ( .A(n_256), .Y(n_391) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x4_ASAP7_75t_L g307 ( .A(n_257), .B(n_308), .Y(n_307) );
NOR2xp67_ASAP7_75t_SL g339 ( .A(n_257), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g412 ( .A(n_257), .B(n_395), .Y(n_412) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_257), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g464 ( .A(n_257), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g331 ( .A(n_258), .Y(n_331) );
INVx4_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g326 ( .A(n_259), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_259), .B(n_324), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_259), .B(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_259), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g409 ( .A(n_263), .B(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
AND2x2_ASAP7_75t_L g443 ( .A(n_268), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g451 ( .A(n_268), .B(n_380), .Y(n_451) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g320 ( .A(n_269), .B(n_305), .Y(n_320) );
AND2x4_ASAP7_75t_L g353 ( .A(n_269), .B(n_287), .Y(n_353) );
INVx1_ASAP7_75t_L g470 ( .A(n_269), .Y(n_470) );
AND2x2_ASAP7_75t_L g356 ( .A(n_271), .B(n_296), .Y(n_356) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g377 ( .A(n_272), .B(n_312), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_281), .B1(n_290), .B2(n_293), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_279), .Y(n_274) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_275), .A2(n_344), .B1(n_452), .B2(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_276), .B(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g345 ( .A(n_276), .B(n_277), .Y(n_345) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_276), .B(n_347), .Y(n_375) );
AOI211xp5_ASAP7_75t_SL g463 ( .A1(n_276), .A2(n_464), .B(n_466), .C(n_467), .Y(n_463) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_277), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_277), .B(n_323), .Y(n_449) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g354 ( .A(n_279), .Y(n_354) );
INVx2_ASAP7_75t_L g410 ( .A(n_280), .Y(n_410) );
AND2x2_ASAP7_75t_L g484 ( .A(n_280), .B(n_477), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_281), .A2(n_433), .B(n_439), .Y(n_432) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g419 ( .A(n_283), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g429 ( .A(n_283), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g336 ( .A(n_284), .B(n_289), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g338 ( .A(n_284), .B(n_305), .Y(n_338) );
AND2x2_ASAP7_75t_L g380 ( .A(n_284), .B(n_305), .Y(n_380) );
INVx2_ASAP7_75t_L g297 ( .A(n_285), .Y(n_297) );
AND2x4_ASAP7_75t_L g303 ( .A(n_285), .B(n_304), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx3_ASAP7_75t_L g295 ( .A(n_287), .Y(n_295) );
INVx3_ASAP7_75t_L g301 ( .A(n_288), .Y(n_301) );
BUFx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_292), .A2(n_398), .B(n_474), .Y(n_478) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_295), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_295), .B(n_370), .Y(n_385) );
OR2x2_ASAP7_75t_L g400 ( .A(n_295), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_295), .B(n_311), .Y(n_407) );
AND2x2_ASAP7_75t_L g363 ( .A(n_296), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_296), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g396 ( .A(n_296), .B(n_365), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_306), .B1(n_309), .B2(n_313), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp67_ASAP7_75t_L g373 ( .A(n_301), .B(n_302), .Y(n_373) );
NOR2xp67_ASAP7_75t_SL g411 ( .A(n_301), .B(n_319), .Y(n_411) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_305), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g314 ( .A(n_307), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g378 ( .A(n_307), .B(n_324), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_307), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g481 ( .A(n_315), .B(n_347), .Y(n_481) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_316), .B(n_427), .Y(n_426) );
NOR2xp67_ASAP7_75t_SL g317 ( .A(n_318), .B(n_341), .Y(n_317) );
OAI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_328), .C(n_337), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_319), .A2(n_372), .B(n_382), .C(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g461 ( .A(n_320), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g372 ( .A(n_324), .B(n_348), .Y(n_372) );
AND2x2_ASAP7_75t_L g459 ( .A(n_324), .B(n_438), .Y(n_459) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g427 ( .A(n_327), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_331), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g401 ( .A(n_336), .Y(n_401) );
NAND2xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_339), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_349), .B1(n_351), .B2(n_354), .C(n_355), .Y(n_341) );
NOR4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .C(n_346), .D(n_348), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g460 ( .A(n_347), .B(n_423), .Y(n_460) );
INVx2_ASAP7_75t_L g466 ( .A(n_347), .Y(n_466) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_350), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g453 ( .A(n_353), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND4xp75_ASAP7_75t_L g358 ( .A(n_359), .B(n_381), .C(n_388), .D(n_397), .Y(n_358) );
OA211x2_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_366), .C(n_374), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_360), .B(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g454 ( .A(n_364), .Y(n_454) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g462 ( .A(n_365), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_373), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_378), .B2(n_379), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_378), .A2(n_429), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g457 ( .A(n_379), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_380), .B(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVxp67_ASAP7_75t_L g455 ( .A(n_391), .Y(n_455) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_395), .B(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_396), .A2(n_459), .B1(n_481), .B2(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND3x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_445), .C(n_458), .Y(n_403) );
NOR3x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_417), .C(n_432), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_413), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_411), .B2(n_412), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_422), .B1(n_424), .B2(n_428), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g476 ( .A(n_426), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g465 ( .A(n_442), .Y(n_465) );
OAI21xp5_ASAP7_75t_SL g473 ( .A1(n_443), .A2(n_474), .B(n_476), .Y(n_473) );
NOR2x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_456), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_450), .B1(n_452), .B2(n_455), .Y(n_446) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_461), .C(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g534 ( .A(n_471), .Y(n_534) );
NOR2x1_ASAP7_75t_SL g471 ( .A(n_472), .B(n_479), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g501 ( .A(n_489), .Y(n_501) );
BUFx2_ASAP7_75t_L g515 ( .A(n_489), .Y(n_515) );
BUFx2_ASAP7_75t_L g833 ( .A(n_489), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x6_ASAP7_75t_SL g528 ( .A(n_490), .B(n_492), .Y(n_528) );
OR2x6_ASAP7_75t_SL g538 ( .A(n_490), .B(n_491), .Y(n_538) );
OR2x2_ASAP7_75t_L g827 ( .A(n_490), .B(n_492), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
CKINVDCx12_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
NOR2x1_ASAP7_75t_R g497 ( .A(n_498), .B(n_499), .Y(n_497) );
CKINVDCx11_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_SL g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_504), .A2(n_511), .B(n_514), .Y(n_510) );
INVx2_ASAP7_75t_L g832 ( .A(n_504), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g831 ( .A(n_506), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
CKINVDCx11_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx8_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_818), .B(n_828), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_526), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_520), .A2(n_820), .B(n_823), .Y(n_819) );
INVxp33_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B1(n_536), .B2(n_539), .Y(n_526) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_527), .A2(n_821), .B(n_822), .Y(n_820) );
CKINVDCx11_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g821 ( .A(n_529), .Y(n_821) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
NAND2x1_ASAP7_75t_SL g822 ( .A(n_537), .B(n_539), .Y(n_822) );
CKINVDCx11_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_710), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_638), .C(n_688), .Y(n_541) );
OAI211xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_573), .B(n_608), .C(n_627), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x2_ASAP7_75t_L g637 ( .A(n_544), .B(n_556), .Y(n_637) );
INVx1_ASAP7_75t_L g768 ( .A(n_544), .Y(n_768) );
NOR2x1p5_ASAP7_75t_L g800 ( .A(n_544), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g613 ( .A(n_545), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g659 ( .A(n_545), .Y(n_659) );
OR2x2_ASAP7_75t_L g663 ( .A(n_545), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_545), .B(n_558), .Y(n_675) );
OR2x2_ASAP7_75t_L g697 ( .A(n_545), .B(n_558), .Y(n_697) );
AND2x4_ASAP7_75t_L g703 ( .A(n_545), .B(n_667), .Y(n_703) );
OR2x2_ASAP7_75t_L g720 ( .A(n_545), .B(n_615), .Y(n_720) );
INVx1_ASAP7_75t_L g755 ( .A(n_545), .Y(n_755) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_545), .Y(n_777) );
OR2x2_ASAP7_75t_L g791 ( .A(n_545), .B(n_724), .Y(n_791) );
AND2x4_ASAP7_75t_SL g795 ( .A(n_545), .B(n_615), .Y(n_795) );
OR2x6_ASAP7_75t_L g545 ( .A(n_546), .B(n_554), .Y(n_545) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g747 ( .A(n_556), .B(n_703), .Y(n_747) );
AND2x2_ASAP7_75t_L g794 ( .A(n_556), .B(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_564), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g612 ( .A(n_558), .Y(n_612) );
AND2x2_ASAP7_75t_L g657 ( .A(n_558), .B(n_564), .Y(n_657) );
INVx2_ASAP7_75t_L g664 ( .A(n_558), .Y(n_664) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_558), .Y(n_785) );
BUFx3_ASAP7_75t_L g801 ( .A(n_558), .Y(n_801) );
INVx2_ASAP7_75t_L g626 ( .A(n_564), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_564), .B(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g724 ( .A(n_564), .B(n_664), .Y(n_724) );
INVx1_ASAP7_75t_L g742 ( .A(n_564), .Y(n_742) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_564), .Y(n_758) );
INVx1_ASAP7_75t_L g780 ( .A(n_564), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_564), .B(n_659), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_564), .B(n_615), .Y(n_817) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_581), .Y(n_574) );
AND2x4_ASAP7_75t_L g631 ( .A(n_575), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g642 ( .A(n_575), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_575), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g682 ( .A(n_575), .B(n_590), .Y(n_682) );
AND2x2_ASAP7_75t_L g692 ( .A(n_575), .B(n_591), .Y(n_692) );
OR2x2_ASAP7_75t_L g772 ( .A(n_575), .B(n_687), .Y(n_772) );
OAI322xp33_ASAP7_75t_L g802 ( .A1(n_575), .A2(n_715), .A3(n_754), .B1(n_787), .B2(n_803), .C1(n_804), .C2(n_805), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_575), .B(n_785), .Y(n_803) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_581), .A2(n_749), .B1(n_753), .B2(n_756), .Y(n_748) );
AOI211xp5_ASAP7_75t_L g808 ( .A1(n_581), .A2(n_809), .B(n_810), .C(n_813), .Y(n_808) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_582), .B(n_590), .Y(n_581) );
AND2x4_ASAP7_75t_L g630 ( .A(n_582), .B(n_600), .Y(n_630) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_582), .Y(n_634) );
INVx5_ASAP7_75t_L g646 ( .A(n_582), .Y(n_646) );
INVx2_ASAP7_75t_L g655 ( .A(n_582), .Y(n_655) );
AND2x2_ASAP7_75t_L g678 ( .A(n_582), .B(n_591), .Y(n_678) );
AND2x2_ASAP7_75t_L g707 ( .A(n_582), .B(n_599), .Y(n_707) );
OR2x2_ASAP7_75t_L g716 ( .A(n_582), .B(n_636), .Y(n_716) );
OR2x2_ASAP7_75t_L g731 ( .A(n_582), .B(n_645), .Y(n_731) );
OR2x6_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_590), .B(n_609), .Y(n_608) );
INVx3_ASAP7_75t_SL g715 ( .A(n_590), .Y(n_715) );
AND2x2_ASAP7_75t_L g738 ( .A(n_590), .B(n_646), .Y(n_738) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_599), .Y(n_590) );
INVx2_ASAP7_75t_L g632 ( .A(n_591), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_591), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g649 ( .A(n_591), .B(n_600), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_591), .B(n_600), .Y(n_687) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_591), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_591), .B(n_646), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_600), .Y(n_668) );
AND2x2_ASAP7_75t_L g752 ( .A(n_600), .B(n_636), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_606), .Y(n_601) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_610), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x6_ASAP7_75t_SL g816 ( .A(n_611), .B(n_817), .Y(n_816) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_612), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_612), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g764 ( .A(n_612), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_613), .A2(n_673), .B1(n_676), .B2(n_683), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_614), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g708 ( .A(n_614), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_614), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_SL g763 ( .A(n_614), .B(n_764), .Y(n_763) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_626), .Y(n_614) );
AND2x2_ASAP7_75t_L g658 ( .A(n_615), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g667 ( .A(n_615), .Y(n_667) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_615), .A2(n_674), .B1(n_726), .B2(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g733 ( .A(n_615), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_615), .B(n_727), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_615), .B(n_657), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_615), .B(n_664), .Y(n_806) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_621), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_633), .B(n_637), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND4xp25_ASAP7_75t_SL g676 ( .A(n_629), .B(n_677), .C(n_679), .D(n_681), .Y(n_676) );
INVx2_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_630), .B(n_737), .Y(n_766) );
AND2x2_ASAP7_75t_L g793 ( .A(n_630), .B(n_631), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_630), .B(n_653), .Y(n_804) );
INVx1_ASAP7_75t_L g669 ( .A(n_631), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_631), .A2(n_694), .B1(n_705), .B2(n_708), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_631), .B(n_644), .C(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_631), .B(n_646), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_631), .B(n_654), .Y(n_797) );
AND2x2_ASAP7_75t_L g729 ( .A(n_632), .B(n_636), .Y(n_729) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_632), .Y(n_790) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g685 ( .A(n_634), .Y(n_685) );
INVx1_ASAP7_75t_L g775 ( .A(n_635), .Y(n_775) );
AND2x2_ASAP7_75t_L g782 ( .A(n_635), .B(n_646), .Y(n_782) );
BUFx2_ASAP7_75t_L g737 ( .A(n_636), .Y(n_737) );
NAND3xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_660), .C(n_672), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_647), .A3(n_650), .B(n_656), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_640), .A2(n_694), .B1(n_698), .B2(n_699), .Y(n_693) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g679 ( .A(n_642), .B(n_680), .Y(n_679) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_642), .B(n_706), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g774 ( .A1(n_643), .A2(n_745), .B(n_775), .C(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_644), .B(n_790), .Y(n_789) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_645), .B(n_653), .Y(n_680) );
AND2x2_ASAP7_75t_L g698 ( .A(n_645), .B(n_678), .Y(n_698) );
AND2x2_ASAP7_75t_L g815 ( .A(n_648), .B(n_737), .Y(n_815) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g671 ( .A(n_649), .B(n_655), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_654), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g746 ( .A(n_654), .B(n_729), .Y(n_746) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_655), .B(n_729), .Y(n_735) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_L g727 ( .A(n_657), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_658), .B(n_758), .Y(n_757) );
AOI32xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_668), .A3(n_669), .B1(n_670), .B2(n_836), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_661), .A2(n_746), .B1(n_782), .B2(n_783), .C(n_786), .Y(n_781) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_664), .Y(n_709) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g674 ( .A(n_666), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g779 ( .A(n_667), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_668), .B(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_670), .A2(n_713), .B1(n_717), .B2(n_721), .C(n_725), .Y(n_712) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_675), .A2(n_689), .B(n_693), .C(n_704), .Y(n_688) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g786 ( .A1(n_681), .A2(n_691), .A3(n_740), .B1(n_787), .B2(n_788), .C1(n_789), .C2(n_791), .Y(n_786) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g813 ( .A1(n_684), .A2(n_814), .B(n_816), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g770 ( .A1(n_690), .A2(n_771), .B(n_773), .C(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g812 ( .A(n_697), .B(n_778), .Y(n_812) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_703), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g787 ( .A(n_703), .Y(n_787) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_707), .A2(n_744), .A3(n_746), .B(n_747), .Y(n_743) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_769), .Y(n_710) );
NAND5xp2_ASAP7_75t_L g711 ( .A(n_712), .B(n_732), .C(n_743), .D(n_748), .E(n_759), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g810 ( .A1(n_715), .A2(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g783 ( .A(n_719), .B(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_736), .C(n_739), .Y(n_732) );
INVxp33_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
OR2x2_ASAP7_75t_L g761 ( .A(n_737), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_740), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_SL g749 ( .A(n_750), .B(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g811 ( .A(n_752), .Y(n_811) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_763), .B(n_765), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_761), .A2(n_766), .B(n_767), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g769 ( .A(n_770), .B(n_781), .C(n_792), .D(n_808), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_779), .B(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g809 ( .A(n_791), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_796), .B2(n_798), .C(n_802), .Y(n_792) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OR2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
INVxp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
endmodule