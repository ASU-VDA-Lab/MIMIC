module fake_jpeg_32108_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_37),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_4),
.B(n_5),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_26),
.C(n_34),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_17),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_24),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_53),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_18),
.C(n_15),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.C(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_27),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_22),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_20),
.B(n_24),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_16),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_66),
.B1(n_54),
.B2(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_32),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_33),
.B1(n_16),
.B2(n_23),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_47),
.C(n_50),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_42),
.B1(n_65),
.B2(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_42),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_81),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_85),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_76),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_75),
.B(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_77),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_81),
.C(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_98),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_74),
.B(n_79),
.C(n_43),
.D(n_59),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_100),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_79),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_94),
.B(n_97),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_100),
.B(n_11),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_105),
.B1(n_9),
.B2(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_63),
.Y(n_108)
);


endmodule