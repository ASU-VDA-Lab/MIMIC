module fake_jpeg_8454_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_30),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_17),
.Y(n_37)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_10),
.C(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_30),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_14),
.B1(n_19),
.B2(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_38),
.B1(n_39),
.B2(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_10),
.A3(n_12),
.B1(n_16),
.B2(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_19),
.B1(n_15),
.B2(n_11),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_25),
.B(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_46),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_9),
.C(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_47),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_13),
.B1(n_22),
.B2(n_16),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_56),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_20),
.B1(n_18),
.B2(n_13),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_71),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_65),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_62),
.Y(n_86)
);

NOR4xp25_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_57),
.C(n_46),
.D(n_49),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_78),
.A3(n_75),
.B1(n_70),
.B2(n_64),
.C1(n_73),
.C2(n_81),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_52),
.B(n_43),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_67),
.B(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_67),
.B1(n_79),
.B2(n_75),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_61),
.B(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_63),
.B1(n_56),
.B2(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

AO221x1_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_59),
.B1(n_54),
.B2(n_64),
.C(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_24),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_85),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_102),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_93),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_105),
.B(n_43),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);

NOR2xp67_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_6),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_7),
.Y(n_110)
);


endmodule