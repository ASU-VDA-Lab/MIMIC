module fake_netlist_6_3182_n_2438 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2438);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2438;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_437;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_1207;
wire n_811;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_100),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_4),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_119),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_169),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_88),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_93),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_44),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_94),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_133),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_84),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_55),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_32),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_74),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_185),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_88),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_219),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_126),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_134),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_21),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_127),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_111),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_54),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_193),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_97),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_159),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_227),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_72),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_168),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_49),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_167),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_151),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_160),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_76),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_194),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_7),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_182),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_82),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_109),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_226),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_112),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_81),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_124),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_162),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_106),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_223),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_32),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_145),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_33),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_40),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_198),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_164),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_9),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_25),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_186),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_46),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_0),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_212),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_104),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_148),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_140),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_59),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_100),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_45),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_10),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_21),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_82),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_117),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_104),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_73),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_116),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_64),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_139),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_78),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_205),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_147),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_217),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_208),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_63),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_9),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_92),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_42),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_68),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_71),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_58),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_61),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_24),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_170),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_44),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_231),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_56),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_166),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_210),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_71),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_47),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_1),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_222),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_171),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_40),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_172),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_197),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_85),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_1),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_45),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_53),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_81),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_174),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_189),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_121),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_78),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_209),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_218),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_106),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_156),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_180),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_6),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_72),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_142),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_53),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_26),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_13),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_24),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_49),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_203),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_184),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_105),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_138),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_27),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_30),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_86),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_136),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_199),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_173),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_20),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_52),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_143),
.Y(n_401)
);

BUFx8_ASAP7_75t_SL g402 ( 
.A(n_18),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_213),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_16),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_202),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_153),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_19),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_94),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_74),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_211),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_230),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_86),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_176),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_61),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_77),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_90),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_187),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_137),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_177),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_3),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_149),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_36),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_113),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_70),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_95),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_110),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_105),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_47),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_56),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_155),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_235),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_181),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_69),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_115),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_4),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_38),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_112),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_50),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_17),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_114),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_34),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_228),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_51),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_34),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_220),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_0),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_120),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_109),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_3),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_67),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_233),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_75),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_196),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_95),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_107),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_43),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_63),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_123),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_135),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_20),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_101),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_15),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_64),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_96),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_303),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_303),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_402),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_303),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_344),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_239),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_303),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_402),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_250),
.B(n_5),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_321),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_237),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_247),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_303),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_303),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_252),
.B(n_5),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_271),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_336),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_274),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_246),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_274),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_371),
.B(n_8),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_274),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_240),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_244),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_252),
.B(n_321),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_271),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_358),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_251),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_255),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_357),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_358),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_364),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_358),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_371),
.B(n_8),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_256),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_357),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_265),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_357),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_337),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_247),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_418),
.B(n_252),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_409),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_371),
.B(n_10),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_266),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_269),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_260),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_397),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_246),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_418),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_260),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_258),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_258),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_270),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_270),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_284),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_361),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_272),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_284),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_302),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_275),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_324),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_278),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_292),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_361),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_292),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_302),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_293),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_L g544 ( 
.A(n_371),
.B(n_11),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_340),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_293),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_285),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_248),
.B(n_11),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_361),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_340),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_295),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_295),
.B(n_13),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_307),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_248),
.B(n_14),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_286),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_297),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_304),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_246),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_307),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_249),
.B(n_254),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_310),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_308),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_308),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_325),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_453),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_311),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_426),
.B(n_14),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_325),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_249),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_331),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_312),
.Y(n_572)
);

INVxp33_ASAP7_75t_SL g573 ( 
.A(n_238),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_453),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_254),
.B(n_15),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_331),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_324),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_316),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_397),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_319),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_329),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_432),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_432),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_342),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_289),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_342),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_399),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_289),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_345),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_345),
.Y(n_590)
);

INVxp33_ASAP7_75t_SL g591 ( 
.A(n_241),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_346),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_488),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_489),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_493),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_494),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_519),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_466),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_540),
.B(n_348),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_526),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_503),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_486),
.B(n_280),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_505),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_570),
.B(n_348),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_504),
.B(n_280),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_561),
.B(n_348),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_490),
.B(n_415),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_516),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_577),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_559),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_468),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_559),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_522),
.B(n_280),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_517),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_504),
.B(n_415),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_471),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_533),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_484),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_R g630 ( 
.A(n_521),
.B(n_330),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_536),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_480),
.B(n_294),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_522),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_478),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_479),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_479),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_587),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_558),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_538),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_547),
.B(n_333),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_555),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_527),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_558),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_579),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_484),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_527),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_528),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_528),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_506),
.B(n_267),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_529),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_556),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_557),
.Y(n_654)
);

AND2x2_ASAP7_75t_SL g655 ( 
.A(n_548),
.B(n_294),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_484),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_415),
.Y(n_658)
);

INVx6_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_507),
.B(n_338),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_531),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_583),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_535),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_534),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_562),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_484),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_567),
.Y(n_668)
);

CKINVDCx16_ASAP7_75t_R g669 ( 
.A(n_481),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_552),
.B(n_250),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_483),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_483),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_507),
.B(n_267),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_534),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_572),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_486),
.A2(n_288),
.B(n_276),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_510),
.B(n_276),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_501),
.B(n_399),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_542),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_539),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_485),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_513),
.B(n_408),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_487),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_545),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_578),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_510),
.B(n_512),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_R g690 ( 
.A(n_580),
.B(n_339),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_633),
.B(n_476),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_633),
.B(n_581),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_659),
.B(n_622),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_634),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_593),
.B(n_573),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_639),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_613),
.B(n_398),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_634),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_596),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_659),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_655),
.B(n_591),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_622),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_655),
.B(n_481),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_639),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_596),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_606),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_606),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_593),
.B(n_475),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_651),
.B(n_549),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_659),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_657),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_655),
.B(n_593),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_643),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_593),
.B(n_524),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_622),
.B(n_512),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_655),
.B(n_491),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_651),
.B(n_549),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_643),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_639),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_599),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_659),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_644),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_659),
.B(n_544),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_644),
.Y(n_724)
);

BUFx4f_ASAP7_75t_L g725 ( 
.A(n_607),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_644),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_659),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_657),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_599),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_607),
.B(n_398),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_601),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_638),
.B(n_491),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_635),
.Y(n_736)
);

AND2x6_ASAP7_75t_L g737 ( 
.A(n_607),
.B(n_398),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_593),
.B(n_537),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_603),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_603),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_618),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_618),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_613),
.B(n_398),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_607),
.B(n_408),
.Y(n_745)
);

INVx6_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_657),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_608),
.B(n_467),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_648),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_635),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_648),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_649),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_638),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_651),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_649),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_660),
.B(n_263),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_616),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_669),
.A2(n_354),
.B1(n_429),
.B2(n_391),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_677),
.B(n_263),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_660),
.B(n_537),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_SL g761 ( 
.A(n_680),
.B(n_552),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_673),
.B(n_514),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_635),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_673),
.B(n_514),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_657),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_624),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_641),
.B(n_472),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_620),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_604),
.B(n_351),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_673),
.B(n_515),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_614),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_657),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_604),
.B(n_351),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_641),
.B(n_585),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_620),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_679),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_616),
.B(n_508),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_679),
.B(n_398),
.Y(n_778)
);

AND2x2_ASAP7_75t_SL g779 ( 
.A(n_669),
.B(n_554),
.Y(n_779)
);

AO22x2_ASAP7_75t_L g780 ( 
.A1(n_680),
.A2(n_474),
.B1(n_454),
.B2(n_456),
.Y(n_780)
);

INVx6_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_667),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_667),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

BUFx4f_ASAP7_75t_L g785 ( 
.A(n_624),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_667),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_679),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_677),
.B(n_353),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_690),
.B(n_588),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_684),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_611),
.B(n_515),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_667),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_667),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_684),
.B(n_469),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_605),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_667),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_609),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_608),
.B(n_470),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_650),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_667),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_636),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_614),
.B(n_353),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_611),
.B(n_518),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_609),
.B(n_495),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_627),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_652),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_636),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_602),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_611),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_602),
.Y(n_814)
);

BUFx4f_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_594),
.B(n_473),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_677),
.B(n_518),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_602),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_631),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_631),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_396),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_637),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_637),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_670),
.B(n_495),
.Y(n_824)
);

NOR2x1p5_ASAP7_75t_L g825 ( 
.A(n_595),
.B(n_520),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_670),
.A2(n_575),
.B1(n_350),
.B2(n_359),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_520),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_602),
.Y(n_828)
);

OAI22xp33_ASAP7_75t_L g829 ( 
.A1(n_597),
.A2(n_454),
.B1(n_456),
.B2(n_264),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_656),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_602),
.B(n_396),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_671),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_598),
.A2(n_482),
.B1(n_497),
.B2(n_442),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_605),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_656),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_626),
.A2(n_288),
.B1(n_306),
.B2(n_291),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_617),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_661),
.B(n_523),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_617),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_615),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_617),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_617),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_625),
.A2(n_568),
.B1(n_426),
.B2(n_243),
.Y(n_843)
);

BUFx4f_ASAP7_75t_L g844 ( 
.A(n_624),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_661),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_SL g846 ( 
.A(n_626),
.B(n_354),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_628),
.B(n_523),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_664),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_690),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_664),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_665),
.B(n_525),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_761),
.A2(n_291),
.B1(n_322),
.B2(n_306),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_813),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_813),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_822),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_797),
.B(n_632),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_745),
.A2(n_566),
.B1(n_574),
.B2(n_550),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_849),
.B(n_640),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_822),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_830),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_702),
.B(n_754),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_725),
.B(n_322),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_725),
.B(n_642),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_753),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_SL g866 ( 
.A1(n_795),
.A2(n_474),
.B1(n_391),
.B2(n_429),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_797),
.B(n_653),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_754),
.B(n_654),
.Y(n_868)
);

O2A1O1Ixp5_ASAP7_75t_L g869 ( 
.A1(n_725),
.A2(n_658),
.B(n_689),
.C(n_341),
.Y(n_869)
);

BUFx5_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_790),
.A2(n_666),
.B1(n_676),
.B2(n_668),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_785),
.B(n_334),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_823),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_790),
.B(n_645),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_776),
.B(n_688),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_776),
.B(n_787),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_787),
.B(n_686),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_709),
.B(n_689),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_835),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_SL g881 ( 
.A1(n_795),
.A2(n_681),
.B1(n_687),
.B2(n_663),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_694),
.B(n_698),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_694),
.B(n_698),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_771),
.B(n_645),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_761),
.A2(n_341),
.B1(n_355),
.B2(n_334),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_756),
.B(n_686),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_760),
.A2(n_355),
.B1(n_383),
.B2(n_360),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_745),
.B(n_442),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_699),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_817),
.A2(n_383),
.B1(n_389),
.B2(n_360),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_823),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_817),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_699),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_821),
.B(n_629),
.Y(n_894)
);

NAND2x1_ASAP7_75t_L g895 ( 
.A(n_746),
.B(n_617),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_821),
.B(n_629),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_705),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_691),
.B(n_686),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_746),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_746),
.A2(n_413),
.B1(n_430),
.B2(n_389),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_821),
.B(n_708),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_746),
.B(n_686),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_705),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_714),
.B(n_645),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_791),
.B(n_686),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_777),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_759),
.B(n_629),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_791),
.B(n_629),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_701),
.A2(n_363),
.B1(n_370),
.B2(n_356),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_712),
.A2(n_374),
.B1(n_375),
.B2(n_372),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_703),
.A2(n_430),
.B(n_413),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_849),
.B(n_695),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_812),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_SL g914 ( 
.A(n_829),
.B(n_245),
.C(n_242),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_791),
.A2(n_806),
.B1(n_770),
.B2(n_762),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_806),
.B(n_646),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_716),
.A2(n_379),
.B1(n_380),
.B2(n_378),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_806),
.B(n_646),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_731),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_709),
.B(n_646),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_847),
.B(n_647),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_717),
.B(n_646),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_762),
.A2(n_434),
.B1(n_445),
.B2(n_431),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_835),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_794),
.A2(n_392),
.B1(n_403),
.B2(n_390),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_845),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_715),
.B(n_674),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_731),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_717),
.B(n_845),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_777),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_715),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_848),
.B(n_646),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_692),
.B(n_647),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_732),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_715),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_764),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_848),
.B(n_630),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_760),
.A2(n_826),
.B1(n_807),
.B2(n_769),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_816),
.B(n_647),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_779),
.A2(n_405),
.B1(n_410),
.B2(n_406),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_840),
.B(n_662),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_779),
.A2(n_411),
.B1(n_419),
.B2(n_417),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_807),
.B(n_662),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_852),
.B(n_630),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_764),
.B(n_658),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_852),
.B(n_610),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_827),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_759),
.B(n_421),
.Y(n_948)
);

AND2x6_ASAP7_75t_SL g949 ( 
.A(n_834),
.B(n_346),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_757),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_759),
.B(n_624),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_788),
.B(n_624),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_732),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_827),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_762),
.A2(n_459),
.B1(n_447),
.B2(n_431),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_773),
.B(n_757),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_713),
.B(n_610),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_788),
.B(n_434),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_718),
.B(n_610),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_711),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_733),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_733),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_734),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_749),
.B(n_751),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_805),
.A2(n_678),
.B(n_682),
.C(n_674),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_770),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_788),
.B(n_445),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_770),
.B(n_451),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_752),
.B(n_612),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_735),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_755),
.B(n_612),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_851),
.B(n_525),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_738),
.B(n_662),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_800),
.B(n_612),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_825),
.B(n_451),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_735),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_802),
.A2(n_458),
.B1(n_624),
.B2(n_359),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_809),
.B(n_619),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_834),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_850),
.B(n_619),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_740),
.B(n_619),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_785),
.B(n_458),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_734),
.B(n_663),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_838),
.Y(n_984)
);

OR2x6_ASAP7_75t_L g985 ( 
.A(n_774),
.B(n_350),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_740),
.B(n_623),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_L g987 ( 
.A(n_846),
.B(n_509),
.C(n_477),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_851),
.B(n_678),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_851),
.B(n_682),
.Y(n_989)
);

AND2x6_ASAP7_75t_SL g990 ( 
.A(n_758),
.B(n_365),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_824),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_730),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_693),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_741),
.B(n_623),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_838),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_741),
.B(n_685),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_SL g997 ( 
.A1(n_720),
.A2(n_687),
.B1(n_681),
.B2(n_395),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_742),
.B(n_623),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_824),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_785),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_697),
.A2(n_624),
.B1(n_366),
.B2(n_384),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_742),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_836),
.A2(n_685),
.B(n_530),
.C(n_365),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_743),
.B(n_624),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_711),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_831),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_697),
.A2(n_624),
.B1(n_384),
.B2(n_385),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_812),
.Y(n_1008)
);

BUFx8_ASAP7_75t_L g1009 ( 
.A(n_743),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_840),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_768),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_744),
.A2(n_385),
.B1(n_386),
.B2(n_366),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_815),
.B(n_301),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_729),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_843),
.B(n_264),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_812),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_846),
.A2(n_401),
.B1(n_301),
.B2(n_671),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_833),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_768),
.B(n_671),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_775),
.B(n_683),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_775),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_784),
.B(n_683),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_784),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_798),
.B(n_683),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_798),
.B(n_672),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_808),
.B(n_672),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_748),
.B(n_789),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_856),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_857),
.B(n_840),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_897),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_856),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_897),
.Y(n_1032)
);

AO22x1_ASAP7_75t_L g1033 ( 
.A1(n_1015),
.A2(n_778),
.B1(n_737),
.B2(n_730),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_938),
.A2(n_780),
.B1(n_744),
.B2(n_808),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_1000),
.B(n_815),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_1014),
.Y(n_1036)
);

INVx6_ASAP7_75t_L g1037 ( 
.A(n_870),
.Y(n_1037)
);

CKINVDCx6p67_ASAP7_75t_R g1038 ( 
.A(n_1010),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_865),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_1010),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_892),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_904),
.B(n_799),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_860),
.Y(n_1043)
);

CKINVDCx11_ASAP7_75t_R g1044 ( 
.A(n_979),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_963),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_860),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_966),
.B(n_767),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_903),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_1000),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_1027),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_867),
.B(n_706),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1006),
.A2(n_780),
.B1(n_819),
.B2(n_810),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_991),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_912),
.B(n_706),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1006),
.B(n_810),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_862),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_945),
.B(n_819),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_999),
.B(n_914),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_873),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_956),
.B(n_706),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_966),
.B(n_700),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_888),
.A2(n_885),
.B1(n_853),
.B2(n_945),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_979),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_879),
.B(n_820),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_873),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_891),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_892),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_903),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_879),
.B(n_936),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_892),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_SL g1071 ( 
.A(n_866),
.B(n_257),
.C(n_253),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_931),
.B(n_700),
.Y(n_1072)
);

AND2x4_ASAP7_75t_SL g1073 ( 
.A(n_874),
.B(n_707),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_SL g1074 ( 
.A1(n_941),
.A2(n_780),
.B1(n_707),
.B2(n_737),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_862),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_1000),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_1000),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_950),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_931),
.B(n_727),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_997),
.B(n_261),
.C(n_259),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_859),
.B(n_707),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_919),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_1000),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_898),
.B(n_820),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_936),
.B(n_841),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_891),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_906),
.B(n_818),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_919),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_913),
.B(n_815),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_999),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_934),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_934),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_953),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_930),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_874),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_939),
.B(n_837),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_953),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_961),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_874),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_882),
.B(n_837),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_961),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_947),
.B(n_780),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_888),
.A2(n_723),
.B(n_273),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_962),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_874),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_901),
.A2(n_844),
.B(n_842),
.C(n_837),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_862),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_983),
.B(n_277),
.C(n_262),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_962),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_SL g1110 ( 
.A(n_1009),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_883),
.B(n_877),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_881),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_954),
.B(n_832),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_921),
.B(n_818),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_927),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_976),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_899),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_889),
.B(n_842),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_901),
.A2(n_737),
.B1(n_730),
.B2(n_778),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_976),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_884),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_915),
.B(n_868),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_871),
.B(n_301),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_889),
.B(n_842),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_899),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1009),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_893),
.B(n_765),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_899),
.Y(n_1128)
);

OR2x4_ASAP7_75t_L g1129 ( 
.A(n_933),
.B(n_386),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1002),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_913),
.B(n_844),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_935),
.B(n_864),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1009),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1002),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_870),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_890),
.A2(n_721),
.B1(n_710),
.B2(n_727),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_985),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_893),
.B(n_765),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_928),
.B(n_765),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_992),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_985),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_895),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_SL g1143 ( 
.A(n_870),
.B(n_301),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_985),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1021),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1021),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_935),
.B(n_710),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_928),
.B(n_792),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_970),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_970),
.Y(n_1150)
);

BUFx8_ASAP7_75t_L g1151 ( 
.A(n_870),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1011),
.B(n_792),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_875),
.B(n_792),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_992),
.B(n_721),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1011),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_SL g1156 ( 
.A(n_943),
.B(n_281),
.C(n_279),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_984),
.B(n_832),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_927),
.B(n_796),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_985),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_858),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_927),
.B(n_796),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1018),
.B(n_818),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_929),
.B(n_796),
.Y(n_1163)
);

AND2x4_ASAP7_75t_SL g1164 ( 
.A(n_989),
.B(n_401),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_864),
.B(n_895),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_SL g1166 ( 
.A(n_973),
.B(n_283),
.C(n_282),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_880),
.B(n_828),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_989),
.B(n_988),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_988),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_870),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_924),
.B(n_828),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_996),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_937),
.B(n_828),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_913),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_854),
.Y(n_1175)
);

OR2x2_ASAP7_75t_SL g1176 ( 
.A(n_990),
.B(n_387),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_926),
.B(n_728),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1008),
.A2(n_844),
.B1(n_781),
.B2(n_728),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_996),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_905),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_887),
.B(n_290),
.C(n_287),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1023),
.B(n_728),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_855),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_995),
.B(n_541),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_972),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_992),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_870),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_870),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_R g1189 ( 
.A(n_944),
.B(n_296),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_SL g1190 ( 
.A(n_968),
.B(n_299),
.C(n_298),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_972),
.B(n_696),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_940),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_949),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1008),
.B(n_739),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_908),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_916),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_R g1197 ( 
.A(n_861),
.B(n_300),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1008),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_942),
.B(n_739),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_992),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_989),
.A2(n_730),
.B1(n_737),
.B2(n_401),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_876),
.B(n_920),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_975),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_922),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_918),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_946),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_964),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_886),
.B(n_696),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_968),
.B(n_704),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_R g1210 ( 
.A(n_951),
.B(n_952),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_975),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_965),
.A2(n_750),
.B(n_763),
.C(n_736),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_981),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1016),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_986),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1016),
.B(n_739),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1016),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_994),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_998),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_878),
.B(n_747),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1026),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1019),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1020),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1106),
.A2(n_907),
.B(n_958),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1114),
.B(n_993),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1089),
.A2(n_907),
.B(n_958),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1069),
.B(n_993),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1214),
.A2(n_1083),
.B(n_1135),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1089),
.A2(n_1131),
.B(n_1035),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1089),
.A2(n_967),
.B(n_863),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1052),
.A2(n_1017),
.B1(n_948),
.B2(n_967),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1212),
.A2(n_900),
.A3(n_1024),
.B(n_1022),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1214),
.A2(n_952),
.B(n_951),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1076),
.B(n_960),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1131),
.A2(n_863),
.B(n_869),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1076),
.B(n_960),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1042),
.A2(n_975),
.B1(n_948),
.B2(n_1013),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1069),
.B(n_923),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1214),
.B(n_1083),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1180),
.A2(n_896),
.B(n_894),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1121),
.B(n_987),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1062),
.A2(n_863),
.B1(n_872),
.B2(n_894),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1207),
.B(n_911),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1135),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1207),
.B(n_911),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1149),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1214),
.B(n_896),
.Y(n_1247)
);

AO21x1_ASAP7_75t_L g1248 ( 
.A1(n_1143),
.A2(n_982),
.B(n_872),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1083),
.A2(n_1005),
.B(n_960),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1169),
.B(n_925),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1135),
.A2(n_1170),
.B(n_1194),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1036),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1111),
.B(n_911),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1180),
.A2(n_982),
.B(n_902),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1135),
.B(n_932),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1149),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1169),
.B(n_975),
.Y(n_1257)
);

AOI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1084),
.A2(n_1220),
.B(n_1092),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1091),
.A2(n_1025),
.B(n_959),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1037),
.A2(n_872),
.B1(n_1013),
.B2(n_910),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1064),
.B(n_955),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1057),
.B(n_1172),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1170),
.A2(n_1005),
.B(n_992),
.Y(n_1263)
);

CKINVDCx9p33_ASAP7_75t_R g1264 ( 
.A(n_1036),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1155),
.A2(n_969),
.A3(n_971),
.B(n_957),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1131),
.A2(n_1004),
.B(n_978),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1045),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1155),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1172),
.B(n_909),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1150),
.A2(n_980),
.B(n_974),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1195),
.A2(n_1003),
.B(n_917),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1037),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1170),
.B(n_1005),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1076),
.B(n_1077),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1170),
.A2(n_783),
.B(n_747),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1150),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1195),
.A2(n_1007),
.B(n_1001),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1044),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1216),
.A2(n_783),
.B(n_747),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1179),
.B(n_1012),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1035),
.A2(n_750),
.B(n_736),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1185),
.B(n_1053),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_SL g1283 ( 
.A1(n_1055),
.A2(n_778),
.B(n_737),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1045),
.Y(n_1284)
);

AO32x2_ASAP7_75t_L g1285 ( 
.A1(n_1052),
.A2(n_803),
.A3(n_786),
.B1(n_783),
.B2(n_778),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1136),
.A2(n_803),
.A3(n_786),
.B1(n_778),
.B2(n_449),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1178),
.A2(n_803),
.B(n_786),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1040),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_801),
.A3(n_804),
.B(n_763),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1035),
.A2(n_804),
.B(n_801),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1174),
.A2(n_772),
.B(n_711),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1091),
.A2(n_811),
.A3(n_719),
.B(n_722),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1039),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1092),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1174),
.A2(n_811),
.B(n_719),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1196),
.A2(n_977),
.B(n_722),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1174),
.A2(n_772),
.B(n_711),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1179),
.B(n_704),
.Y(n_1298)
);

AOI21xp33_ASAP7_75t_L g1299 ( 
.A1(n_1160),
.A2(n_309),
.B(n_305),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1198),
.A2(n_726),
.B(n_724),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1049),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1151),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1030),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1196),
.A2(n_726),
.B(n_724),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1063),
.B(n_401),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1185),
.B(n_268),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1097),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1122),
.A2(n_778),
.B(n_737),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1191),
.B(n_543),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1210),
.B(n_711),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1078),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1123),
.A2(n_315),
.B(n_313),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1198),
.A2(n_492),
.B(n_487),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1049),
.B(n_772),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1191),
.B(n_1168),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1097),
.A2(n_675),
.B(n_672),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1198),
.A2(n_496),
.B(n_492),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1223),
.B(n_1202),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1104),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1073),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1217),
.A2(n_1077),
.B(n_1076),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1049),
.B(n_772),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1030),
.Y(n_1323)
);

AOI211x1_ASAP7_75t_L g1324 ( 
.A1(n_1102),
.A2(n_387),
.B(n_448),
.C(n_449),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1223),
.B(n_814),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1143),
.A2(n_407),
.B(n_388),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1217),
.A2(n_782),
.B(n_772),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1202),
.B(n_814),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1217),
.A2(n_793),
.B(n_782),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1077),
.A2(n_793),
.B(n_782),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1034),
.A2(n_498),
.B(n_496),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1104),
.Y(n_1332)
);

INVx3_ASAP7_75t_SL g1333 ( 
.A(n_1110),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_730),
.B(n_766),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1168),
.B(n_543),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1077),
.A2(n_793),
.B(n_782),
.Y(n_1336)
);

AND2x6_ASAP7_75t_SL g1337 ( 
.A(n_1102),
.B(n_388),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1127),
.A2(n_499),
.B(n_498),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1037),
.A2(n_781),
.B1(n_793),
.B2(n_782),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1138),
.A2(n_500),
.B(n_499),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1049),
.A2(n_793),
.B(n_814),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1053),
.B(n_317),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1100),
.A2(n_766),
.B(n_814),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1139),
.A2(n_502),
.B(n_500),
.Y(n_1344)
);

AO21x1_ASAP7_75t_L g1345 ( 
.A1(n_1034),
.A2(n_433),
.B(n_407),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1167),
.A2(n_766),
.B(n_814),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_502),
.B(n_675),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1109),
.Y(n_1348)
);

OA22x2_ASAP7_75t_L g1349 ( 
.A1(n_1160),
.A2(n_464),
.B1(n_440),
.B2(n_463),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1168),
.A2(n_730),
.B1(n_781),
.B2(n_839),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1171),
.A2(n_766),
.B(n_839),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1168),
.B(n_268),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1163),
.A2(n_766),
.B(n_839),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1205),
.A2(n_675),
.B(n_438),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1199),
.A2(n_438),
.B(n_433),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1049),
.B(n_839),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1037),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1109),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1162),
.B(n_839),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1221),
.B(n_781),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1187),
.A2(n_448),
.B(n_440),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1187),
.A2(n_462),
.B(n_452),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1152),
.A2(n_551),
.B(n_546),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1188),
.A2(n_1186),
.B(n_1140),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1221),
.B(n_318),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1130),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1209),
.A2(n_462),
.B(n_452),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1107),
.A2(n_425),
.B1(n_323),
.B2(n_326),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1074),
.A2(n_463),
.B1(n_464),
.B2(n_589),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1103),
.A2(n_1119),
.B(n_1130),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1188),
.A2(n_551),
.B(n_546),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1118),
.A2(n_560),
.B(n_553),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1222),
.B(n_320),
.Y(n_1373)
);

BUFx4_ASAP7_75t_SL g1374 ( 
.A(n_1126),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1124),
.A2(n_560),
.B(n_553),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1222),
.B(n_327),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1206),
.B(n_328),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1032),
.A2(n_564),
.B(n_563),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1145),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1209),
.A2(n_564),
.B(n_563),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1113),
.B(n_565),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1107),
.A2(n_423),
.B1(n_335),
.B2(n_343),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1206),
.B(n_332),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1145),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1151),
.B(n_347),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1032),
.A2(n_569),
.B(n_565),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1146),
.A2(n_592),
.A3(n_590),
.B(n_589),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1094),
.B(n_569),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1048),
.A2(n_576),
.B(n_571),
.Y(n_1389)
);

INVx5_ASAP7_75t_L g1390 ( 
.A(n_1140),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1056),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1048),
.A2(n_576),
.B(n_571),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1078),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_R g1394 ( 
.A(n_1278),
.B(n_1063),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1347),
.A2(n_1082),
.B(n_1068),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1315),
.B(n_1056),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1347),
.A2(n_1082),
.B(n_1068),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1229),
.A2(n_1093),
.B(n_1088),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1252),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1372),
.A2(n_1146),
.B(n_1093),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1229),
.A2(n_1098),
.B(n_1088),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1237),
.A2(n_1058),
.B(n_1123),
.C(n_1181),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1244),
.A2(n_1165),
.B(n_1132),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1276),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1318),
.B(n_1095),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1355),
.A2(n_1060),
.B(n_1051),
.C(n_1029),
.Y(n_1406)
);

NAND3x1_ASAP7_75t_L g1407 ( 
.A(n_1241),
.B(n_1080),
.C(n_1071),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1267),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1295),
.A2(n_1101),
.B(n_1098),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1228),
.A2(n_1075),
.B(n_1151),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1261),
.A2(n_1075),
.B1(n_1192),
.B2(n_1115),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1299),
.A2(n_1141),
.B(n_1144),
.C(n_1054),
.Y(n_1412)
);

AO21x1_ASAP7_75t_L g1413 ( 
.A1(n_1242),
.A2(n_1208),
.B(n_1031),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1295),
.A2(n_1300),
.B(n_1290),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1278),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1227),
.B(n_1095),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1225),
.A2(n_1115),
.B1(n_1159),
.B2(n_1137),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1282),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1300),
.A2(n_1116),
.B(n_1101),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1281),
.A2(n_1120),
.B(n_1116),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1246),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1281),
.A2(n_1134),
.B(n_1120),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1293),
.B(n_1081),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1345),
.A2(n_1134),
.B(n_1213),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1290),
.A2(n_1031),
.B(n_1028),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1305),
.B(n_1166),
.C(n_1156),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1250),
.A2(n_1159),
.B1(n_1137),
.B2(n_1132),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1313),
.A2(n_1043),
.B(n_1028),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1252),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1244),
.A2(n_1251),
.B(n_1273),
.Y(n_1431)
);

NOR2x1_ASAP7_75t_L g1432 ( 
.A(n_1288),
.B(n_1040),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1246),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1315),
.B(n_1113),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1313),
.A2(n_1046),
.B(n_1043),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1243),
.A2(n_1182),
.B(n_1177),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1248),
.A2(n_1119),
.B(n_1153),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1309),
.B(n_1050),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1317),
.A2(n_1059),
.B(n_1046),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1333),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1317),
.A2(n_1065),
.B(n_1059),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1333),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1235),
.A2(n_1066),
.B(n_1065),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1357),
.Y(n_1444)
);

NOR2x1_ASAP7_75t_R g1445 ( 
.A(n_1288),
.B(n_1126),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1256),
.Y(n_1446)
);

AOI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1258),
.A2(n_1259),
.B(n_1231),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1235),
.A2(n_1316),
.B(n_1226),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1250),
.A2(n_1132),
.B1(n_1090),
.B2(n_1087),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1226),
.A2(n_1086),
.B(n_1066),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1230),
.A2(n_1086),
.B(n_1208),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1230),
.A2(n_1215),
.B(n_1213),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1262),
.B(n_1105),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1224),
.A2(n_1218),
.B(n_1215),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1268),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1312),
.A2(n_1105),
.B1(n_1099),
.B2(n_1183),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1374),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1294),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1231),
.A2(n_1219),
.A3(n_1218),
.B(n_1085),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1244),
.B(n_1041),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1224),
.A2(n_1219),
.B(n_1067),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1311),
.A2(n_1081),
.B1(n_1129),
.B2(n_1203),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1264),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1309),
.B(n_1157),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1264),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1393),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1245),
.A2(n_1157),
.B(n_1204),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1244),
.B(n_1357),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1335),
.B(n_1158),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1271),
.A2(n_1204),
.B(n_1132),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1367),
.A2(n_1190),
.B(n_1108),
.C(n_1164),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1303),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1257),
.A2(n_1175),
.B1(n_1183),
.B2(n_1050),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1357),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1338),
.A2(n_1067),
.B(n_1041),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1269),
.A2(n_1164),
.B(n_1073),
.C(n_1175),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1338),
.A2(n_1067),
.B(n_1041),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1357),
.A2(n_1244),
.B1(n_1238),
.B2(n_1391),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1381),
.B(n_1050),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1381),
.B(n_1050),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1357),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1307),
.Y(n_1482)
);

AO21x1_ASAP7_75t_L g1483 ( 
.A1(n_1253),
.A2(n_1147),
.B(n_1184),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1282),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1273),
.A2(n_1165),
.B(n_1132),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1303),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1340),
.A2(n_1070),
.B(n_1117),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1363),
.A2(n_1096),
.B(n_1189),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1340),
.A2(n_1070),
.B(n_1117),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1344),
.A2(n_1070),
.B(n_1117),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1260),
.A2(n_1033),
.B(n_1184),
.C(n_1125),
.Y(n_1491)
);

AOI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1372),
.A2(n_1375),
.B(n_1363),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1293),
.B(n_1090),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1240),
.A2(n_1165),
.B(n_1151),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1335),
.B(n_1158),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1391),
.B(n_1272),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1323),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1342),
.A2(n_1112),
.B1(n_1133),
.B2(n_1203),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1342),
.B(n_1129),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1323),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1272),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1391),
.A2(n_1047),
.B1(n_1165),
.B2(n_1129),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1301),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1378),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1377),
.B(n_1211),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1344),
.A2(n_1128),
.B(n_1125),
.Y(n_1506)
);

BUFx2_ASAP7_75t_R g1507 ( 
.A(n_1385),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1375),
.A2(n_1128),
.B(n_1125),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1319),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1380),
.B(n_1158),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1383),
.B(n_1211),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1301),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1378),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1332),
.Y(n_1514)
);

CKINVDCx9p33_ASAP7_75t_R g1515 ( 
.A(n_1365),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_SL g1516 ( 
.A1(n_1239),
.A2(n_1165),
.B(n_1079),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1348),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_1337),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1386),
.A2(n_586),
.B(n_584),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1388),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1233),
.A2(n_1128),
.B(n_1142),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1354),
.A2(n_1158),
.B(n_1161),
.C(n_1201),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1386),
.A2(n_586),
.B(n_584),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1280),
.A2(n_1047),
.B1(n_1061),
.B2(n_1161),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1389),
.A2(n_1392),
.B(n_1254),
.Y(n_1525)
);

AO31x2_ASAP7_75t_L g1526 ( 
.A1(n_1326),
.A2(n_1287),
.A3(n_1359),
.B(n_1361),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1389),
.Y(n_1527)
);

AO31x2_ASAP7_75t_L g1528 ( 
.A1(n_1362),
.A2(n_1358),
.A3(n_1379),
.B(n_1366),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1266),
.A2(n_1142),
.B(n_1154),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1306),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1301),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1320),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1247),
.A2(n_1186),
.B(n_1140),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1392),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1369),
.B(n_1161),
.Y(n_1535)
);

INVx8_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1247),
.A2(n_1186),
.B(n_1140),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1352),
.A2(n_1047),
.B1(n_1197),
.B2(n_1161),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1369),
.B(n_1047),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1266),
.A2(n_1142),
.B(n_1154),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1272),
.B(n_1047),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1249),
.A2(n_1186),
.B(n_1140),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1239),
.B(n_1186),
.Y(n_1543)
);

AO32x2_ASAP7_75t_L g1544 ( 
.A1(n_1285),
.A2(n_1176),
.A3(n_1033),
.B1(n_1038),
.B2(n_268),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1302),
.B(n_1061),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1301),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1384),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_1373),
.B(n_1133),
.Y(n_1548)
);

INVx4_ASAP7_75t_SL g1549 ( 
.A(n_1292),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1387),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1369),
.B(n_1147),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1321),
.A2(n_592),
.B(n_590),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1376),
.A2(n_1061),
.B1(n_1079),
.B2(n_1072),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_L g1554 ( 
.A(n_1368),
.B(n_1382),
.C(n_1324),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1385),
.A2(n_1061),
.B1(n_1147),
.B2(n_1072),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1304),
.A2(n_1147),
.B(n_1079),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1279),
.A2(n_1275),
.B(n_1364),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1298),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1283),
.A2(n_1200),
.B(n_1079),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1308),
.A2(n_1072),
.B(n_352),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1277),
.A2(n_1072),
.B(n_362),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1292),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1328),
.B(n_1038),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1255),
.A2(n_1263),
.B(n_1353),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1296),
.A2(n_420),
.B(n_367),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1331),
.B(n_268),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1331),
.A2(n_1200),
.B(n_1176),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1390),
.B(n_1200),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1390),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1349),
.A2(n_1193),
.B1(n_416),
.B2(n_461),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1349),
.A2(n_1193),
.B1(n_314),
.B2(n_460),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1255),
.A2(n_1200),
.B(n_232),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1370),
.B(n_1232),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1371),
.A2(n_414),
.B(n_457),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1291),
.A2(n_1200),
.B(n_224),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1387),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1320),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1341),
.B(n_118),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1520),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1499),
.A2(n_1370),
.B1(n_314),
.B2(n_1320),
.Y(n_1580)
);

CKINVDCx6p67_ASAP7_75t_R g1581 ( 
.A(n_1415),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1463),
.A2(n_314),
.B1(n_1274),
.B2(n_444),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1434),
.B(n_1387),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_SL g1584 ( 
.A(n_1415),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1428),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1404),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1408),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1530),
.A2(n_1325),
.B1(n_373),
.B2(n_376),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1458),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1418),
.A2(n_1310),
.B1(n_1274),
.B2(n_1236),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1482),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1421),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1449),
.B(n_1479),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1536),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1484),
.A2(n_1310),
.B1(n_1234),
.B2(n_1236),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1509),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1464),
.B(n_1360),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1514),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1554),
.A2(n_314),
.B1(n_1270),
.B2(n_381),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1571),
.A2(n_349),
.B1(n_368),
.B2(n_400),
.C(n_404),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1468),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_R g1603 ( 
.A(n_1465),
.B(n_1270),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1405),
.B(n_1387),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1402),
.A2(n_435),
.B1(n_428),
.B2(n_427),
.C(n_424),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1413),
.A2(n_1334),
.B(n_1314),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1570),
.A2(n_369),
.B1(n_455),
.B2(n_446),
.C(n_443),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1410),
.B(n_1234),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1448),
.A2(n_1327),
.B(n_1297),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1517),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1464),
.B(n_377),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1426),
.A2(n_1270),
.B1(n_439),
.B2(n_436),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1492),
.A2(n_1314),
.B(n_1322),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1505),
.A2(n_382),
.B1(n_393),
.B2(n_394),
.C(n_412),
.Y(n_1614)
);

INVx6_ASAP7_75t_L g1615 ( 
.A(n_1481),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1468),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1547),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1407),
.A2(n_437),
.B1(n_1350),
.B2(n_1322),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_SL g1620 ( 
.A1(n_1471),
.A2(n_1356),
.B(n_1285),
.C(n_1286),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1481),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1481),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1493),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1473),
.A2(n_1390),
.B1(n_1356),
.B2(n_1339),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1405),
.B(n_1265),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1446),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1541),
.B(n_1390),
.Y(n_1627)
);

NOR2x1p5_ASAP7_75t_L g1628 ( 
.A(n_1511),
.B(n_1285),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1438),
.A2(n_1330),
.B1(n_1336),
.B2(n_1329),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1480),
.A2(n_1343),
.B1(n_1346),
.B2(n_1351),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1446),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1427),
.A2(n_1286),
.B1(n_1232),
.B2(n_1265),
.Y(n_1632)
);

OAI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1411),
.A2(n_1286),
.B1(n_1232),
.B2(n_18),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1541),
.B(n_1292),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1472),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1481),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1408),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1453),
.B(n_1265),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1472),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1453),
.B(n_1265),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1535),
.B(n_1551),
.Y(n_1641)
);

NAND2xp33_ASAP7_75t_R g1642 ( 
.A(n_1465),
.B(n_1556),
.Y(n_1642)
);

CKINVDCx11_ASAP7_75t_R g1643 ( 
.A(n_1518),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1539),
.A2(n_1286),
.B1(n_1232),
.B2(n_1292),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1412),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1416),
.B(n_1289),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1462),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1539),
.A2(n_1289),
.B1(n_23),
.B2(n_29),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1456),
.A2(n_1289),
.B1(n_30),
.B2(n_31),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1566),
.A2(n_1289),
.B1(n_31),
.B2(n_33),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1566),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1455),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1416),
.B(n_35),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1466),
.B(n_37),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1469),
.B(n_37),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1536),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1466),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1469),
.B(n_1495),
.Y(n_1658)
);

AND2x2_ASAP7_75t_SL g1659 ( 
.A(n_1556),
.B(n_38),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1396),
.B(n_39),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1563),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_1661)
);

CKINVDCx8_ASAP7_75t_R g1662 ( 
.A(n_1440),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1448),
.A2(n_221),
.B(n_216),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1463),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1396),
.B(n_48),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1440),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1498),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1535),
.B(n_215),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1538),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1568),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1495),
.A2(n_57),
.B1(n_60),
.B2(n_62),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1430),
.B(n_60),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1431),
.A2(n_214),
.B(n_201),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1548),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.C(n_67),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1394),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1396),
.B(n_69),
.Y(n_1676)
);

AOI222xp33_ASAP7_75t_L g1677 ( 
.A1(n_1518),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.C1(n_77),
.C2(n_79),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1406),
.B(n_79),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1495),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1518),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1536),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1423),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1510),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_1683)
);

BUFx8_ASAP7_75t_L g1684 ( 
.A(n_1503),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1497),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1497),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1510),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1541),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1502),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_1689)
);

AOI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1561),
.A2(n_1470),
.B(n_1524),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1558),
.B(n_99),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1551),
.B(n_144),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1433),
.B(n_1558),
.Y(n_1693)
);

BUFx2_ASAP7_75t_SL g1694 ( 
.A(n_1399),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1486),
.B(n_200),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1442),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1496),
.B(n_141),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1476),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.C(n_108),
.Y(n_1698)
);

AOI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1492),
.A2(n_152),
.B(n_191),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1568),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1399),
.B(n_102),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1417),
.B(n_103),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1407),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1500),
.B(n_192),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1545),
.B(n_113),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1562),
.Y(n_1706)
);

OR2x6_ASAP7_75t_L g1707 ( 
.A(n_1410),
.B(n_158),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1536),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1568),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1503),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_R g1711 ( 
.A(n_1556),
.B(n_161),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1545),
.A2(n_1567),
.B1(n_1553),
.B2(n_1565),
.Y(n_1712)
);

BUFx12f_ASAP7_75t_L g1713 ( 
.A(n_1457),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1545),
.A2(n_1567),
.B1(n_1565),
.B2(n_1483),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_L g1715 ( 
.A(n_1522),
.B(n_1403),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1555),
.A2(n_114),
.B1(n_122),
.B2(n_129),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1467),
.A2(n_1413),
.B1(n_1485),
.B2(n_1436),
.C(n_1491),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1432),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1528),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_R g1720 ( 
.A(n_1578),
.B(n_130),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1496),
.B(n_131),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1516),
.A2(n_132),
.B(n_154),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1507),
.A2(n_165),
.B1(n_175),
.B2(n_178),
.Y(n_1723)
);

O2A1O1Ixp5_ASAP7_75t_SL g1724 ( 
.A1(n_1550),
.A2(n_1576),
.B(n_1527),
.C(n_1478),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1461),
.A2(n_179),
.B(n_183),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1567),
.A2(n_1565),
.B1(n_1483),
.B2(n_1494),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1442),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1496),
.B(n_1501),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1577),
.B(n_1532),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1494),
.A2(n_1424),
.B1(n_1578),
.B2(n_1574),
.Y(n_1730)
);

NAND3x1_ASAP7_75t_L g1731 ( 
.A(n_1515),
.B(n_188),
.C(n_1447),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1578),
.A2(n_1532),
.B1(n_1574),
.B2(n_1560),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1457),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1544),
.B(n_1528),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1516),
.A2(n_1578),
.B1(n_1543),
.B2(n_1573),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1424),
.A2(n_1574),
.B1(n_1560),
.B2(n_1501),
.Y(n_1736)
);

OR2x6_ASAP7_75t_L g1737 ( 
.A(n_1572),
.B(n_1543),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1542),
.A2(n_1557),
.B(n_1537),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1560),
.A2(n_1501),
.B1(n_1437),
.B2(n_1573),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1528),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1460),
.A2(n_1474),
.B1(n_1444),
.B2(n_1546),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1437),
.A2(n_1488),
.B1(n_1546),
.B2(n_1512),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1460),
.A2(n_1474),
.B1(n_1444),
.B2(n_1569),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1528),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1531),
.Y(n_1745)
);

CKINVDCx8_ASAP7_75t_R g1746 ( 
.A(n_1531),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1488),
.A2(n_1549),
.B1(n_1572),
.B2(n_1552),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1460),
.A2(n_1569),
.B1(n_1533),
.B2(n_1447),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1451),
.A2(n_1552),
.B(n_1452),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1531),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_L g1751 ( 
.A(n_1531),
.B(n_1569),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1564),
.B(n_1575),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1544),
.B(n_1528),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1531),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1544),
.B(n_1459),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1454),
.A2(n_1575),
.B(n_1451),
.C(n_1452),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1459),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1544),
.B(n_1459),
.Y(n_1758)
);

AO31x2_ASAP7_75t_L g1759 ( 
.A1(n_1527),
.A2(n_1504),
.A3(n_1534),
.B(n_1513),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_L g1760 ( 
.A(n_1400),
.B(n_1525),
.C(n_1504),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1445),
.B(n_1488),
.Y(n_1761)
);

INVx4_ASAP7_75t_SL g1762 ( 
.A(n_1459),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1450),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1459),
.B(n_1526),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1557),
.A2(n_1564),
.B(n_1540),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1544),
.A2(n_1521),
.B1(n_1559),
.B2(n_1540),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1549),
.A2(n_1559),
.B1(n_1534),
.B2(n_1513),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1400),
.A2(n_1525),
.B1(n_1519),
.B2(n_1523),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1549),
.A2(n_1521),
.B1(n_1400),
.B2(n_1525),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1450),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1398),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1519),
.A2(n_1523),
.B1(n_1526),
.B2(n_1549),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1398),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1529),
.A2(n_1508),
.B1(n_1477),
.B2(n_1475),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1678),
.A2(n_1475),
.B(n_1477),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1698),
.A2(n_1659),
.B1(n_1667),
.B2(n_1669),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1715),
.A2(n_1529),
.B(n_1461),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1623),
.B(n_1526),
.Y(n_1779)
);

INVx5_ASAP7_75t_SL g1780 ( 
.A(n_1581),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1717),
.A2(n_1443),
.B(n_1414),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1647),
.A2(n_1526),
.B1(n_1397),
.B2(n_1395),
.C(n_1443),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1401),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1677),
.A2(n_1523),
.B1(n_1519),
.B2(n_1395),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1607),
.A2(n_1508),
.B1(n_1490),
.B2(n_1489),
.C(n_1487),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1659),
.A2(n_1490),
.B1(n_1489),
.B2(n_1487),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1582),
.A2(n_1441),
.B1(n_1439),
.B2(n_1435),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_1584),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1601),
.A2(n_1506),
.B1(n_1397),
.B2(n_1401),
.C(n_1425),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1615),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1590),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1675),
.A2(n_1661),
.B1(n_1645),
.B2(n_1674),
.C(n_1664),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1720),
.A2(n_1441),
.B1(n_1439),
.B2(n_1435),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1612),
.A2(n_1429),
.B1(n_1425),
.B2(n_1420),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1680),
.A2(n_1429),
.B1(n_1419),
.B2(n_1409),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1682),
.A2(n_1409),
.B1(n_1419),
.B2(n_1422),
.C(n_1703),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1592),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_SL g1799 ( 
.A1(n_1715),
.A2(n_1702),
.B1(n_1716),
.B2(n_1649),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1678),
.A2(n_1605),
.B1(n_1651),
.B2(n_1687),
.C(n_1683),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1722),
.A2(n_1690),
.B(n_1600),
.C(n_1689),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1597),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1618),
.A2(n_1614),
.B1(n_1662),
.B2(n_1729),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1580),
.A2(n_1594),
.B(n_1761),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1723),
.A2(n_1718),
.B1(n_1761),
.B2(n_1666),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1733),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1599),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1608),
.A2(n_1751),
.B(n_1630),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1641),
.B(n_1655),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1587),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1688),
.A2(n_1679),
.B1(n_1671),
.B2(n_1633),
.C(n_1648),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1701),
.B(n_1660),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1611),
.A2(n_1720),
.B1(n_1653),
.B2(n_1650),
.C(n_1732),
.Y(n_1814)
);

OAI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1711),
.A2(n_1642),
.B1(n_1603),
.B2(n_1691),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1684),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1610),
.Y(n_1817)
);

AOI222xp33_ASAP7_75t_L g1818 ( 
.A1(n_1594),
.A2(n_1579),
.B1(n_1598),
.B2(n_1588),
.C1(n_1583),
.C2(n_1637),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1652),
.Y(n_1819)
);

OAI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1707),
.A2(n_1705),
.B1(n_1604),
.B2(n_1665),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1591),
.B(n_1596),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1711),
.A2(n_1730),
.B1(n_1676),
.B2(n_1672),
.C(n_1707),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1707),
.A2(n_1583),
.B1(n_1581),
.B2(n_1585),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1662),
.A2(n_1718),
.B1(n_1746),
.B2(n_1731),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1736),
.A2(n_1642),
.B(n_1646),
.Y(n_1825)
);

OAI211xp5_ASAP7_75t_L g1826 ( 
.A1(n_1654),
.A2(n_1657),
.B(n_1726),
.C(n_1643),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1746),
.A2(n_1731),
.B1(n_1696),
.B2(n_1727),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1668),
.A2(n_1692),
.B1(n_1707),
.B2(n_1735),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_SL g1829 ( 
.A1(n_1668),
.A2(n_1692),
.B1(n_1697),
.B2(n_1721),
.Y(n_1829)
);

BUFx12f_ASAP7_75t_L g1830 ( 
.A(n_1733),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1608),
.A2(n_1751),
.B(n_1629),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1643),
.A2(n_1666),
.B1(n_1697),
.B2(n_1721),
.Y(n_1832)
);

OAI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1603),
.A2(n_1638),
.B1(n_1640),
.B2(n_1625),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1620),
.A2(n_1632),
.B1(n_1673),
.B2(n_1714),
.C(n_1712),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1697),
.A2(n_1721),
.B1(n_1694),
.B2(n_1684),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1628),
.A2(n_1663),
.B(n_1704),
.C(n_1695),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1706),
.Y(n_1837)
);

OAI211xp5_ASAP7_75t_L g1838 ( 
.A1(n_1742),
.A2(n_1739),
.B(n_1620),
.C(n_1710),
.Y(n_1838)
);

A2O1A1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1663),
.A2(n_1704),
.B(n_1695),
.C(n_1624),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1634),
.A2(n_1693),
.B1(n_1713),
.B2(n_1728),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1670),
.B(n_1700),
.Y(n_1841)
);

OAI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1644),
.A2(n_1747),
.B(n_1693),
.C(n_1744),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1627),
.A2(n_1699),
.B(n_1753),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1634),
.A2(n_1713),
.B1(n_1627),
.B2(n_1709),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1719),
.A2(n_1740),
.B1(n_1773),
.B2(n_1634),
.C(n_1748),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1706),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1724),
.B(n_1684),
.C(n_1741),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1608),
.A2(n_1709),
.B1(n_1700),
.B2(n_1670),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1627),
.A2(n_1709),
.B1(n_1685),
.B2(n_1593),
.Y(n_1849)
);

OAI21xp33_ASAP7_75t_L g1850 ( 
.A1(n_1764),
.A2(n_1769),
.B(n_1757),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1734),
.A2(n_1753),
.B(n_1745),
.C(n_1766),
.Y(n_1851)
);

OAI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1608),
.A2(n_1615),
.B1(n_1621),
.B2(n_1636),
.Y(n_1852)
);

OAI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1621),
.A2(n_1636),
.B1(n_1622),
.B2(n_1595),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1622),
.A2(n_1752),
.B1(n_1749),
.B2(n_1767),
.C(n_1775),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1743),
.A2(n_1589),
.B1(n_1616),
.B2(n_1602),
.Y(n_1855)
);

BUFx12f_ASAP7_75t_L g1856 ( 
.A(n_1595),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1750),
.B(n_1754),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1595),
.A2(n_1708),
.B1(n_1656),
.B2(n_1681),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1737),
.A2(n_1656),
.B1(n_1681),
.B2(n_1708),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1756),
.A2(n_1760),
.B(n_1770),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1737),
.A2(n_1589),
.B1(n_1616),
.B2(n_1602),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1589),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1602),
.Y(n_1863)
);

BUFx12f_ASAP7_75t_L g1864 ( 
.A(n_1752),
.Y(n_1864)
);

AO31x2_ASAP7_75t_L g1865 ( 
.A1(n_1756),
.A2(n_1768),
.A3(n_1771),
.B(n_1763),
.Y(n_1865)
);

OAI221xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1752),
.A2(n_1758),
.B1(n_1734),
.B2(n_1755),
.C(n_1616),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1626),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1626),
.B(n_1685),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1631),
.A2(n_1686),
.B1(n_1639),
.B2(n_1635),
.Y(n_1869)
);

AOI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1635),
.A2(n_1774),
.B(n_1772),
.C(n_1619),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1619),
.B(n_1762),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1759),
.Y(n_1872)
);

AOI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1772),
.A2(n_1613),
.B1(n_1762),
.B2(n_1606),
.C(n_1725),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1606),
.A2(n_1725),
.B1(n_1762),
.B2(n_1609),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1606),
.A2(n_1042),
.B1(n_1192),
.B2(n_691),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1725),
.A2(n_1677),
.B1(n_1042),
.B2(n_655),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1698),
.A2(n_1042),
.B1(n_1123),
.B2(n_1305),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1623),
.B(n_1042),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1715),
.A2(n_1228),
.B(n_1244),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1880)
);

AOI33xp33_ASAP7_75t_L g1881 ( 
.A1(n_1680),
.A2(n_826),
.A3(n_829),
.B1(n_1571),
.B2(n_1675),
.B3(n_1651),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1706),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1677),
.A2(n_1042),
.B1(n_655),
.B2(n_1664),
.Y(n_1883)
);

NAND2x1p5_ASAP7_75t_L g1884 ( 
.A(n_1589),
.B(n_1602),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1677),
.B(n_1042),
.C(n_691),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1615),
.Y(n_1887)
);

OAI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1607),
.A2(n_691),
.B1(n_1042),
.B2(n_1305),
.C(n_794),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1698),
.A2(n_1042),
.B1(n_1123),
.B2(n_1305),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1698),
.A2(n_1042),
.B1(n_1123),
.B2(n_1305),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1623),
.B(n_1418),
.Y(n_1891)
);

AOI222xp33_ASAP7_75t_L g1892 ( 
.A1(n_1664),
.A2(n_655),
.B1(n_794),
.B2(n_1042),
.C1(n_670),
.C2(n_761),
.Y(n_1892)
);

OAI222xp33_ASAP7_75t_L g1893 ( 
.A1(n_1698),
.A2(n_1667),
.B1(n_1674),
.B2(n_1664),
.C1(n_1680),
.C2(n_1703),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1720),
.A2(n_1698),
.B1(n_1674),
.B2(n_1123),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1607),
.A2(n_691),
.B1(n_1042),
.B2(n_1305),
.C(n_794),
.Y(n_1895)
);

OAI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1720),
.A2(n_1698),
.B1(n_1674),
.B2(n_1123),
.Y(n_1896)
);

OAI211xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1677),
.A2(n_1080),
.B(n_1299),
.C(n_1607),
.Y(n_1897)
);

OAI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1607),
.A2(n_691),
.B1(n_1042),
.B2(n_1305),
.C(n_794),
.Y(n_1898)
);

OAI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1607),
.A2(n_691),
.B1(n_1042),
.B2(n_1305),
.C(n_794),
.Y(n_1899)
);

NAND3xp33_ASAP7_75t_L g1900 ( 
.A(n_1677),
.B(n_1042),
.C(n_691),
.Y(n_1900)
);

OAI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1720),
.A2(n_1698),
.B1(n_1674),
.B2(n_1123),
.Y(n_1901)
);

OAI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1678),
.A2(n_691),
.B(n_1042),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1623),
.B(n_1418),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1659),
.B(n_1042),
.Y(n_1904)
);

AOI21xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1677),
.A2(n_939),
.B(n_1042),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1615),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1584),
.Y(n_1907)
);

INVx5_ASAP7_75t_SL g1908 ( 
.A(n_1581),
.Y(n_1908)
);

OAI22xp33_ASAP7_75t_SL g1909 ( 
.A1(n_1698),
.A2(n_1123),
.B1(n_1678),
.B2(n_1305),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1720),
.A2(n_1042),
.B1(n_1192),
.B2(n_691),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1684),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1623),
.B(n_1418),
.Y(n_1912)
);

OR2x6_ASAP7_75t_L g1913 ( 
.A(n_1608),
.B(n_1410),
.Y(n_1913)
);

AOI222xp33_ASAP7_75t_L g1914 ( 
.A1(n_1664),
.A2(n_655),
.B1(n_794),
.B2(n_1042),
.C1(n_670),
.C2(n_761),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1587),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1733),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1647),
.A2(n_1042),
.B1(n_691),
.B2(n_1015),
.C(n_829),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1677),
.A2(n_1042),
.B1(n_655),
.B2(n_1664),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1715),
.A2(n_1228),
.B(n_1244),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1677),
.A2(n_1042),
.B1(n_655),
.B2(n_1664),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1677),
.A2(n_1042),
.B1(n_655),
.B2(n_1664),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1677),
.A2(n_691),
.B(n_1042),
.C(n_826),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_L g1923 ( 
.A(n_1677),
.B(n_1042),
.C(n_691),
.Y(n_1923)
);

NAND2x1_ASAP7_75t_L g1924 ( 
.A(n_1707),
.B(n_1410),
.Y(n_1924)
);

OA21x2_ASAP7_75t_L g1925 ( 
.A1(n_1717),
.A2(n_1749),
.B(n_1756),
.Y(n_1925)
);

AOI222xp33_ASAP7_75t_L g1926 ( 
.A1(n_1664),
.A2(n_655),
.B1(n_794),
.B2(n_1042),
.C1(n_670),
.C2(n_761),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1759),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1677),
.A2(n_1042),
.B1(n_655),
.B2(n_1664),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1698),
.A2(n_1042),
.B1(n_1123),
.B2(n_1305),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1586),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1586),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1647),
.A2(n_1042),
.B1(n_691),
.B2(n_1015),
.C(n_829),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1617),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1733),
.Y(n_1934)
);

AO21x2_ASAP7_75t_L g1935 ( 
.A1(n_1738),
.A2(n_1765),
.B(n_1749),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1586),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1698),
.A2(n_1042),
.B1(n_1123),
.B2(n_1305),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1938)
);

OAI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1607),
.A2(n_691),
.B1(n_1042),
.B2(n_1305),
.C(n_794),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1779),
.B(n_1866),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1872),
.B(n_1925),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1871),
.B(n_1851),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1851),
.B(n_1810),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1802),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1885),
.A2(n_1900),
.B1(n_1923),
.B2(n_1883),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1927),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1837),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1883),
.A2(n_1918),
.B1(n_1921),
.B2(n_1920),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1837),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1913),
.B(n_1783),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1864),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1882),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1882),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1930),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1865),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1918),
.A2(n_1920),
.B1(n_1921),
.B2(n_1928),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1931),
.B(n_1936),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1798),
.B(n_1803),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1808),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1862),
.Y(n_1960)
);

OAI321xp33_ASAP7_75t_L g1961 ( 
.A1(n_1928),
.A2(n_1896),
.A3(n_1901),
.B1(n_1894),
.B2(n_1922),
.C(n_1902),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1876),
.A2(n_1910),
.B1(n_1889),
.B2(n_1937),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1817),
.B(n_1792),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1783),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1913),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1897),
.A2(n_1939),
.B1(n_1895),
.B2(n_1899),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1846),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1925),
.B(n_1850),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1861),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1880),
.B(n_1886),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1938),
.B(n_1925),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1913),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1855),
.Y(n_1974)
);

INVxp67_ASAP7_75t_SL g1975 ( 
.A(n_1821),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1809),
.B(n_1831),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1888),
.A2(n_1898),
.B1(n_1932),
.B2(n_1917),
.C(n_1929),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1833),
.B(n_1854),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1860),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1833),
.B(n_1891),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1841),
.B(n_1867),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1863),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1903),
.B(n_1912),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1933),
.B(n_1813),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1840),
.B(n_1860),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1840),
.B(n_1860),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1781),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1868),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1836),
.B(n_1776),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1849),
.B(n_1844),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1821),
.B(n_1843),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1924),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1849),
.B(n_1844),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1878),
.B(n_1815),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1884),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1781),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1869),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1811),
.B(n_1915),
.Y(n_1999)
);

OR2x6_ASAP7_75t_L g2000 ( 
.A(n_1879),
.B(n_1919),
.Y(n_2000)
);

AO31x2_ASAP7_75t_L g2001 ( 
.A1(n_1795),
.A2(n_1787),
.A3(n_1778),
.B(n_1836),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1857),
.B(n_1870),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1848),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1848),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1781),
.Y(n_2005)
);

AOI222xp33_ASAP7_75t_L g2006 ( 
.A1(n_1800),
.A2(n_1812),
.B1(n_1893),
.B2(n_1793),
.C1(n_1894),
.C2(n_1896),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1935),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1852),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1878),
.B(n_1815),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1794),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1852),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1875),
.B(n_1805),
.Y(n_2012)
);

OAI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1905),
.A2(n_1901),
.B1(n_1814),
.B2(n_1822),
.Y(n_2013)
);

INVxp67_ASAP7_75t_R g2014 ( 
.A(n_1859),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1842),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1820),
.B(n_1818),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1935),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1873),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1904),
.B(n_1838),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1853),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_1847),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1823),
.B(n_1874),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1856),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1790),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1785),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1853),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1823),
.B(n_1828),
.Y(n_2027)
);

AO21x2_ASAP7_75t_L g2028 ( 
.A1(n_1839),
.A2(n_1904),
.B(n_1801),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1816),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1782),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1786),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1874),
.B(n_1816),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1826),
.B(n_1908),
.Y(n_2033)
);

AND2x4_ASAP7_75t_SL g2034 ( 
.A(n_1832),
.B(n_1906),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1834),
.B(n_1876),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1967),
.A2(n_1978),
.B1(n_1962),
.B2(n_2013),
.C(n_1945),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1960),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1950),
.B(n_1911),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1954),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1996),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1978),
.A2(n_1926),
.B1(n_1914),
.B2(n_1892),
.Y(n_2041)
);

AOI33xp33_ASAP7_75t_L g2042 ( 
.A1(n_2013),
.A2(n_1877),
.A3(n_1890),
.B1(n_1777),
.B2(n_1799),
.B3(n_1784),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1948),
.A2(n_1909),
.B1(n_1804),
.B2(n_1829),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1954),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1956),
.A2(n_1832),
.B1(n_1806),
.B2(n_1835),
.Y(n_2045)
);

OA21x2_ASAP7_75t_L g2046 ( 
.A1(n_1997),
.A2(n_2005),
.B(n_2017),
.Y(n_2046)
);

OAI211xp5_ASAP7_75t_L g2047 ( 
.A1(n_2006),
.A2(n_1784),
.B(n_1827),
.C(n_1881),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1984),
.B(n_1999),
.Y(n_2048)
);

INVx5_ASAP7_75t_SL g2049 ( 
.A(n_1977),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1984),
.B(n_1780),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1981),
.B(n_1995),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_L g2052 ( 
.A1(n_2006),
.A2(n_1881),
.B(n_1796),
.C(n_1824),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_1961),
.B(n_1906),
.C(n_1791),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_1999),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1962),
.A2(n_1780),
.B1(n_1908),
.B2(n_1791),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_2021),
.A2(n_1887),
.B1(n_1797),
.B2(n_1796),
.C(n_1858),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_2012),
.A2(n_1780),
.B1(n_1908),
.B2(n_1887),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1972),
.B(n_1807),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_2010),
.B(n_1858),
.Y(n_2059)
);

AOI211xp5_ASAP7_75t_SL g2060 ( 
.A1(n_1961),
.A2(n_1789),
.B(n_1907),
.C(n_1830),
.Y(n_2060)
);

OAI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2012),
.A2(n_1916),
.B1(n_1934),
.B2(n_2016),
.C(n_2035),
.Y(n_2061)
);

OAI21xp33_ASAP7_75t_L g2062 ( 
.A1(n_2016),
.A2(n_2030),
.B(n_2035),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1947),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1985),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1972),
.B(n_1964),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1947),
.Y(n_2066)
);

NOR2x1_ASAP7_75t_SL g2067 ( 
.A(n_1977),
.B(n_2028),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1949),
.Y(n_2068)
);

AOI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2021),
.A2(n_2030),
.B1(n_1976),
.B2(n_2019),
.C(n_2018),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1976),
.A2(n_2028),
.B1(n_2019),
.B2(n_2009),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_L g2071 ( 
.A(n_2018),
.B(n_1995),
.C(n_2009),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1944),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1964),
.B(n_1986),
.Y(n_2073)
);

INVx5_ASAP7_75t_SL g2074 ( 
.A(n_1977),
.Y(n_2074)
);

OAI221xp5_ASAP7_75t_L g2075 ( 
.A1(n_1979),
.A2(n_1975),
.B1(n_1992),
.B2(n_2015),
.C(n_1977),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_SL g2076 ( 
.A(n_1960),
.B(n_1983),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1960),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1949),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1983),
.B(n_2029),
.Y(n_2079)
);

CKINVDCx20_ASAP7_75t_R g2080 ( 
.A(n_1983),
.Y(n_2080)
);

NOR2x1_ASAP7_75t_SL g2081 ( 
.A(n_1977),
.B(n_2028),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_SL g2082 ( 
.A(n_2028),
.B(n_1992),
.Y(n_2082)
);

BUFx3_ASAP7_75t_L g2083 ( 
.A(n_2029),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1986),
.B(n_1987),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1979),
.A2(n_2015),
.B1(n_2033),
.B2(n_2014),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1987),
.B(n_2010),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1985),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2027),
.A2(n_1974),
.B1(n_1975),
.B2(n_1994),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1952),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1989),
.B(n_1982),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1952),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_2029),
.B(n_1951),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1989),
.B(n_1982),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1953),
.Y(n_2094)
);

OAI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_1981),
.A2(n_2025),
.B1(n_2024),
.B2(n_2033),
.C(n_2031),
.Y(n_2095)
);

AOI33xp33_ASAP7_75t_L g2096 ( 
.A1(n_2031),
.A2(n_2025),
.A3(n_2024),
.B1(n_1990),
.B2(n_1943),
.B3(n_2027),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_2025),
.B(n_2024),
.C(n_2011),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1996),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2000),
.A2(n_1990),
.B(n_1974),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1953),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1968),
.Y(n_2101)
);

OAI211xp5_ASAP7_75t_L g2102 ( 
.A1(n_2020),
.A2(n_2026),
.B(n_1969),
.C(n_1980),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2008),
.A2(n_1991),
.B1(n_1994),
.B2(n_2034),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2000),
.A2(n_1993),
.B(n_1990),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1946),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_1969),
.B(n_1941),
.Y(n_2106)
);

AOI31xp33_ASAP7_75t_L g2107 ( 
.A1(n_1943),
.A2(n_1942),
.A3(n_2002),
.B(n_1940),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_1966),
.Y(n_2108)
);

OAI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_1951),
.A2(n_2008),
.B1(n_2022),
.B2(n_2026),
.C(n_2020),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_1950),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_2023),
.Y(n_2111)
);

NAND4xp25_ASAP7_75t_L g2112 ( 
.A(n_1940),
.B(n_2011),
.C(n_1998),
.D(n_1958),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2000),
.A2(n_1990),
.B(n_1980),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2101),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_2106),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2106),
.B(n_1941),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2046),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2084),
.B(n_1988),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2084),
.B(n_1988),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2065),
.B(n_2001),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_2067),
.B(n_1993),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2051),
.B(n_1959),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2046),
.Y(n_2123)
);

INVx4_ASAP7_75t_L g2124 ( 
.A(n_2037),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2039),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2065),
.B(n_2001),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2070),
.B(n_1959),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2070),
.B(n_1963),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2046),
.Y(n_2129)
);

NOR2xp67_ASAP7_75t_L g2130 ( 
.A(n_2102),
.B(n_2007),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2086),
.B(n_1963),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2086),
.B(n_2073),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2067),
.B(n_2081),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2046),
.B(n_1955),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2073),
.B(n_2001),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2048),
.B(n_2063),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2090),
.B(n_2093),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2072),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2090),
.B(n_2001),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2063),
.B(n_1957),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2093),
.B(n_2001),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2039),
.Y(n_2142)
);

NOR2x1_ASAP7_75t_L g2143 ( 
.A(n_2104),
.B(n_1993),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2082),
.B(n_2001),
.Y(n_2144)
);

AND2x4_ASAP7_75t_SL g2145 ( 
.A(n_2080),
.B(n_2032),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2044),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2082),
.B(n_1997),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2081),
.B(n_1997),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2105),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2044),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2066),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2066),
.Y(n_2152)
);

AND4x1_ASAP7_75t_L g2153 ( 
.A(n_2036),
.B(n_2014),
.C(n_1942),
.D(n_2002),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2058),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2068),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_2040),
.Y(n_2156)
);

NAND4xp25_ASAP7_75t_L g2157 ( 
.A(n_2069),
.B(n_2041),
.C(n_2042),
.D(n_2047),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2068),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2078),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2127),
.B(n_2108),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2159),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2122),
.B(n_2088),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2132),
.B(n_2110),
.Y(n_2163)
);

INVxp67_ASAP7_75t_L g2164 ( 
.A(n_2122),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2127),
.B(n_2054),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2132),
.B(n_2110),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2118),
.B(n_2078),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2117),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2159),
.Y(n_2169)
);

INVx1_ASAP7_75t_SL g2170 ( 
.A(n_2154),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_2157),
.B(n_2061),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2136),
.B(n_2088),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_2133),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2136),
.B(n_2062),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2132),
.B(n_2058),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2120),
.B(n_2049),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2118),
.B(n_2089),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2159),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2158),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2118),
.B(n_2089),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2120),
.B(n_2049),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2120),
.B(n_2049),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_2157),
.B(n_2107),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2128),
.B(n_2071),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2128),
.B(n_2064),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2117),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2116),
.B(n_2091),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2156),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2158),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2158),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2158),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2125),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2125),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2131),
.B(n_2087),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2131),
.B(n_2096),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2116),
.B(n_2091),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2116),
.B(n_2094),
.Y(n_2197)
);

AOI32xp33_ASAP7_75t_L g2198 ( 
.A1(n_2135),
.A2(n_2060),
.A3(n_2045),
.B1(n_2043),
.B2(n_2109),
.Y(n_2198)
);

BUFx2_ASAP7_75t_L g2199 ( 
.A(n_2143),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2142),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2126),
.B(n_2139),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2126),
.B(n_2049),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2115),
.B(n_2094),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2117),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2117),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2134),
.Y(n_2206)
);

OAI33xp33_ASAP7_75t_L g2207 ( 
.A1(n_2151),
.A2(n_2112),
.A3(n_2085),
.B1(n_2097),
.B2(n_2100),
.B3(n_2050),
.Y(n_2207)
);

OAI21xp33_ASAP7_75t_SL g2208 ( 
.A1(n_2130),
.A2(n_2143),
.B(n_2154),
.Y(n_2208)
);

INVxp67_ASAP7_75t_L g2209 ( 
.A(n_2140),
.Y(n_2209)
);

NAND2x1_ASAP7_75t_SL g2210 ( 
.A(n_2130),
.B(n_2040),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2142),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2115),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2146),
.Y(n_2213)
);

INVxp67_ASAP7_75t_SL g2214 ( 
.A(n_2140),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2126),
.B(n_2139),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2139),
.B(n_2074),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2176),
.B(n_2135),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2161),
.Y(n_2218)
);

NAND4xp25_ASAP7_75t_L g2219 ( 
.A(n_2183),
.B(n_2171),
.C(n_2198),
.D(n_2055),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2176),
.B(n_2135),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2181),
.B(n_2141),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2169),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2169),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2178),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2174),
.B(n_2141),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2195),
.B(n_2141),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2207),
.B(n_2124),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2206),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2181),
.B(n_2119),
.Y(n_2229)
);

AOI21xp33_ASAP7_75t_L g2230 ( 
.A1(n_2208),
.A2(n_2095),
.B(n_2075),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2184),
.B(n_2119),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2182),
.B(n_2119),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2182),
.B(n_2137),
.Y(n_2233)
);

AOI32xp33_ASAP7_75t_L g2234 ( 
.A1(n_2208),
.A2(n_2144),
.A3(n_2145),
.B1(n_2076),
.B2(n_2153),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2172),
.B(n_2162),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2178),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2192),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2164),
.B(n_2124),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2198),
.B(n_2153),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2206),
.Y(n_2240)
);

NOR3xp33_ASAP7_75t_L g2241 ( 
.A(n_2199),
.B(n_2052),
.C(n_2124),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2192),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2202),
.B(n_2201),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2165),
.B(n_2137),
.Y(n_2244)
);

INVx2_ASAP7_75t_SL g2245 ( 
.A(n_2210),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2193),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2179),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2202),
.B(n_2137),
.Y(n_2248)
);

OAI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2210),
.A2(n_2099),
.B(n_2113),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2193),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2200),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2200),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2201),
.B(n_2144),
.Y(n_2253)
);

INVx5_ASAP7_75t_L g2254 ( 
.A(n_2199),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2165),
.B(n_2124),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2211),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2179),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2211),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2209),
.B(n_2124),
.Y(n_2259)
);

INVxp67_ASAP7_75t_SL g2260 ( 
.A(n_2212),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_SL g2261 ( 
.A(n_2175),
.B(n_2080),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2185),
.B(n_2037),
.Y(n_2262)
);

OR2x6_ASAP7_75t_L g2263 ( 
.A(n_2188),
.B(n_2104),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2213),
.Y(n_2264)
);

NAND3xp33_ASAP7_75t_L g2265 ( 
.A(n_2160),
.B(n_2056),
.C(n_2144),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2215),
.B(n_2121),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2194),
.B(n_2077),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2214),
.B(n_1971),
.Y(n_2268)
);

CKINVDCx16_ASAP7_75t_R g2269 ( 
.A(n_2170),
.Y(n_2269)
);

NAND4xp25_ASAP7_75t_SL g2270 ( 
.A(n_2216),
.B(n_2103),
.C(n_2057),
.D(n_2053),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2215),
.B(n_2121),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2243),
.B(n_2216),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2237),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2237),
.Y(n_2274)
);

NOR4xp25_ASAP7_75t_L g2275 ( 
.A(n_2239),
.B(n_2188),
.C(n_2160),
.D(n_2173),
.Y(n_2275)
);

AOI222xp33_ASAP7_75t_L g2276 ( 
.A1(n_2227),
.A2(n_2145),
.B1(n_2003),
.B2(n_2004),
.C1(n_2175),
.C2(n_1970),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2269),
.A2(n_2145),
.B1(n_2074),
.B2(n_2059),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2235),
.B(n_2163),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_SL g2279 ( 
.A1(n_2269),
.A2(n_2074),
.B1(n_2145),
.B2(n_2003),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2241),
.B(n_2163),
.Y(n_2280)
);

AOI21xp33_ASAP7_75t_SL g2281 ( 
.A1(n_2230),
.A2(n_2079),
.B(n_2092),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2243),
.B(n_2166),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2254),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2222),
.Y(n_2284)
);

AOI221xp5_ASAP7_75t_L g2285 ( 
.A1(n_2219),
.A2(n_2133),
.B1(n_2147),
.B2(n_2213),
.C(n_2173),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2242),
.Y(n_2286)
);

AOI221x1_ASAP7_75t_L g2287 ( 
.A1(n_2261),
.A2(n_2173),
.B1(n_2151),
.B2(n_2152),
.C(n_2155),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2242),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2270),
.A2(n_2133),
.B(n_2121),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2254),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2217),
.B(n_2166),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2246),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2262),
.B(n_2038),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2246),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2244),
.B(n_2187),
.Y(n_2295)
);

AOI222xp33_ASAP7_75t_L g2296 ( 
.A1(n_2265),
.A2(n_2004),
.B1(n_1970),
.B2(n_2133),
.C1(n_1991),
.C2(n_2074),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2217),
.B(n_2220),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2222),
.Y(n_2298)
);

OAI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_2234),
.A2(n_2133),
.B(n_2059),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_2255),
.Y(n_2300)
);

AOI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2249),
.A2(n_2133),
.B(n_2121),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2220),
.B(n_2173),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2260),
.B(n_2203),
.Y(n_2303)
);

O2A1O1Ixp33_ASAP7_75t_L g2304 ( 
.A1(n_2245),
.A2(n_2000),
.B(n_2022),
.C(n_2147),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2250),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2221),
.B(n_2121),
.Y(n_2306)
);

AOI31xp33_ASAP7_75t_L g2307 ( 
.A1(n_2245),
.A2(n_2238),
.A3(n_2259),
.B(n_2226),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2250),
.Y(n_2308)
);

AOI32xp33_ASAP7_75t_L g2309 ( 
.A1(n_2233),
.A2(n_2121),
.A3(n_2148),
.B1(n_2147),
.B2(n_2038),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2231),
.B(n_2187),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2223),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2223),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2224),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2276),
.B(n_2233),
.Y(n_2314)
);

OAI32xp33_ASAP7_75t_L g2315 ( 
.A1(n_2280),
.A2(n_2225),
.A3(n_2218),
.B1(n_2266),
.B2(n_2271),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2275),
.B(n_2248),
.Y(n_2316)
);

AOI32xp33_ASAP7_75t_L g2317 ( 
.A1(n_2299),
.A2(n_2248),
.A3(n_2221),
.B1(n_2229),
.B2(n_2232),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2284),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_SL g2319 ( 
.A1(n_2307),
.A2(n_2267),
.B(n_1951),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2300),
.B(n_2229),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2281),
.B(n_2254),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2284),
.Y(n_2322)
);

NAND3x2_ASAP7_75t_L g2323 ( 
.A(n_2272),
.B(n_2271),
.C(n_2266),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2298),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2279),
.A2(n_2263),
.B1(n_2232),
.B2(n_2254),
.Y(n_2325)
);

OAI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2287),
.A2(n_2254),
.B1(n_2263),
.B2(n_2000),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2298),
.Y(n_2327)
);

INVxp67_ASAP7_75t_SL g2328 ( 
.A(n_2283),
.Y(n_2328)
);

OAI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2287),
.A2(n_2254),
.B1(n_2263),
.B2(n_2000),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2278),
.B(n_2268),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2282),
.B(n_2218),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2272),
.B(n_2263),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2302),
.Y(n_2333)
);

OAI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2296),
.A2(n_2264),
.B(n_2258),
.Y(n_2334)
);

OAI21xp5_ASAP7_75t_L g2335 ( 
.A1(n_2289),
.A2(n_2264),
.B(n_2258),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2303),
.B(n_2228),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2277),
.A2(n_2256),
.B(n_2252),
.Y(n_2337)
);

OAI221xp5_ASAP7_75t_L g2338 ( 
.A1(n_2285),
.A2(n_2240),
.B1(n_2228),
.B2(n_2252),
.C(n_2251),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2311),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2295),
.B(n_2240),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2311),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2302),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2282),
.B(n_2253),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_2283),
.B(n_2111),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2316),
.B(n_2297),
.Y(n_2345)
);

NOR4xp25_ASAP7_75t_SL g2346 ( 
.A(n_2319),
.B(n_2273),
.C(n_2274),
.D(n_2286),
.Y(n_2346)
);

CKINVDCx20_ASAP7_75t_L g2347 ( 
.A(n_2321),
.Y(n_2347)
);

XOR2x2_ASAP7_75t_L g2348 ( 
.A(n_2321),
.B(n_2314),
.Y(n_2348)
);

OAI322xp33_ASAP7_75t_L g2349 ( 
.A1(n_2326),
.A2(n_2329),
.A3(n_2338),
.B1(n_2331),
.B2(n_2336),
.C1(n_2322),
.C2(n_2339),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2318),
.Y(n_2350)
);

XNOR2x2_ASAP7_75t_L g2351 ( 
.A(n_2334),
.B(n_2290),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2324),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2328),
.B(n_2290),
.Y(n_2353)
);

NAND4xp25_ASAP7_75t_SL g2354 ( 
.A(n_2317),
.B(n_2309),
.C(n_2301),
.D(n_2304),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2333),
.B(n_2297),
.Y(n_2355)
);

INVx1_ASAP7_75t_SL g2356 ( 
.A(n_2320),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2327),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_SL g2358 ( 
.A(n_2315),
.B(n_2293),
.C(n_2292),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2341),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2333),
.B(n_2291),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2342),
.B(n_2291),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2342),
.B(n_2288),
.Y(n_2362)
);

BUFx2_ASAP7_75t_L g2363 ( 
.A(n_2344),
.Y(n_2363)
);

AO22x1_ASAP7_75t_L g2364 ( 
.A1(n_2335),
.A2(n_2308),
.B1(n_2294),
.B2(n_2305),
.Y(n_2364)
);

INVx3_ASAP7_75t_SL g2365 ( 
.A(n_2336),
.Y(n_2365)
);

OAI32xp33_ASAP7_75t_L g2366 ( 
.A1(n_2344),
.A2(n_2310),
.A3(n_2295),
.B1(n_2313),
.B2(n_2312),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2330),
.B(n_2310),
.Y(n_2367)
);

XNOR2xp5_ASAP7_75t_L g2368 ( 
.A(n_2323),
.B(n_2038),
.Y(n_2368)
);

INVxp67_ASAP7_75t_L g2369 ( 
.A(n_2363),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2365),
.B(n_2343),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2355),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2358),
.A2(n_2325),
.B1(n_2332),
.B2(n_2326),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2355),
.Y(n_2373)
);

BUFx2_ASAP7_75t_SL g2374 ( 
.A(n_2353),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2353),
.Y(n_2375)
);

NOR4xp25_ASAP7_75t_L g2376 ( 
.A(n_2349),
.B(n_2329),
.C(n_2340),
.D(n_2312),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_L g2377 ( 
.A(n_2365),
.B(n_2332),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2353),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2346),
.A2(n_2337),
.B(n_2313),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2356),
.B(n_2343),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_2360),
.Y(n_2381)
);

NAND4xp75_ASAP7_75t_SL g2382 ( 
.A(n_2351),
.B(n_2306),
.C(n_2253),
.D(n_2148),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2348),
.B(n_2345),
.Y(n_2383)
);

OAI221xp5_ASAP7_75t_L g2384 ( 
.A1(n_2376),
.A2(n_2358),
.B1(n_2348),
.B2(n_2351),
.C(n_2361),
.Y(n_2384)
);

AOI221xp5_ASAP7_75t_SL g2385 ( 
.A1(n_2379),
.A2(n_2366),
.B1(n_2362),
.B2(n_2352),
.C(n_2357),
.Y(n_2385)
);

NOR2x1_ASAP7_75t_L g2386 ( 
.A(n_2374),
.B(n_2350),
.Y(n_2386)
);

NAND5xp2_ASAP7_75t_L g2387 ( 
.A(n_2372),
.B(n_2347),
.C(n_2359),
.D(n_2354),
.E(n_2364),
.Y(n_2387)
);

AOI222xp33_ASAP7_75t_L g2388 ( 
.A1(n_2383),
.A2(n_2368),
.B1(n_2367),
.B2(n_2306),
.C1(n_2251),
.C2(n_2256),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_2375),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_SL g2390 ( 
.A1(n_2377),
.A2(n_1951),
.B1(n_2111),
.B2(n_2023),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2369),
.B(n_2224),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2370),
.A2(n_2236),
.B1(n_2247),
.B2(n_2257),
.Y(n_2392)
);

A2O1A1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2382),
.A2(n_2236),
.B(n_2148),
.C(n_2257),
.Y(n_2393)
);

AOI211xp5_ASAP7_75t_L g2394 ( 
.A1(n_2371),
.A2(n_2023),
.B(n_2247),
.C(n_2203),
.Y(n_2394)
);

AOI222xp33_ASAP7_75t_L g2395 ( 
.A1(n_2381),
.A2(n_2205),
.B1(n_2204),
.B2(n_2168),
.C1(n_2186),
.C2(n_2034),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2380),
.B(n_2023),
.Y(n_2396)
);

AOI322xp5_ASAP7_75t_L g2397 ( 
.A1(n_2373),
.A2(n_2168),
.A3(n_2204),
.B1(n_2186),
.B2(n_2205),
.C1(n_2123),
.C2(n_2129),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2387),
.B(n_2378),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2389),
.B(n_2196),
.Y(n_2399)
);

AOI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2384),
.A2(n_2382),
.B1(n_2032),
.B2(n_1965),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2386),
.B(n_2189),
.Y(n_2401)
);

NAND4xp25_ASAP7_75t_L g2402 ( 
.A(n_2385),
.B(n_2032),
.C(n_2083),
.D(n_2156),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2389),
.B(n_2189),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2389),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_2391),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2396),
.Y(n_2406)
);

NOR2xp67_ASAP7_75t_L g2407 ( 
.A(n_2404),
.B(n_2392),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2399),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_R g2409 ( 
.A(n_2405),
.B(n_2023),
.Y(n_2409)
);

XNOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2406),
.B(n_2388),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2402),
.A2(n_2390),
.B(n_2394),
.Y(n_2411)
);

OA22x2_ASAP7_75t_L g2412 ( 
.A1(n_2403),
.A2(n_2395),
.B1(n_2393),
.B2(n_2397),
.Y(n_2412)
);

OAI21xp33_ASAP7_75t_L g2413 ( 
.A1(n_2398),
.A2(n_2205),
.B(n_2204),
.Y(n_2413)
);

AND3x4_ASAP7_75t_L g2414 ( 
.A(n_2401),
.B(n_2083),
.C(n_2032),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2408),
.B(n_2410),
.Y(n_2415)
);

NAND4xp25_ASAP7_75t_L g2416 ( 
.A(n_2411),
.B(n_2400),
.C(n_2403),
.D(n_2156),
.Y(n_2416)
);

NAND3xp33_ASAP7_75t_SL g2417 ( 
.A(n_2409),
.B(n_2168),
.C(n_2186),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2412),
.A2(n_2023),
.B1(n_1973),
.B2(n_1965),
.Y(n_2418)
);

NOR3xp33_ASAP7_75t_L g2419 ( 
.A(n_2407),
.B(n_2040),
.C(n_2098),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2414),
.A2(n_2413),
.B1(n_2167),
.B2(n_2177),
.Y(n_2420)
);

NOR4xp25_ASAP7_75t_L g2421 ( 
.A(n_2408),
.B(n_2191),
.C(n_2190),
.D(n_2197),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2418),
.A2(n_2197),
.B1(n_2196),
.B2(n_2180),
.Y(n_2422)
);

BUFx2_ASAP7_75t_L g2423 ( 
.A(n_2415),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2416),
.A2(n_2156),
.B1(n_2190),
.B2(n_2191),
.Y(n_2424)
);

A2O1A1Ixp33_ASAP7_75t_L g2425 ( 
.A1(n_2419),
.A2(n_2180),
.B(n_2177),
.C(n_2167),
.Y(n_2425)
);

CKINVDCx16_ASAP7_75t_R g2426 ( 
.A(n_2417),
.Y(n_2426)
);

NAND3xp33_ASAP7_75t_L g2427 ( 
.A(n_2423),
.B(n_2420),
.C(n_2421),
.Y(n_2427)
);

CKINVDCx20_ASAP7_75t_R g2428 ( 
.A(n_2426),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2428),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2429),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2429),
.B(n_2427),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2430),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2431),
.A2(n_2424),
.B(n_2422),
.Y(n_2433)
);

AOI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2433),
.A2(n_2425),
.B(n_2129),
.Y(n_2434)
);

OAI222xp33_ASAP7_75t_L g2435 ( 
.A1(n_2432),
.A2(n_2123),
.B1(n_2129),
.B2(n_2149),
.C1(n_2152),
.C2(n_2155),
.Y(n_2435)
);

NAND3xp33_ASAP7_75t_L g2436 ( 
.A(n_2434),
.B(n_2129),
.C(n_2123),
.Y(n_2436)
);

OAI221xp5_ASAP7_75t_R g2437 ( 
.A1(n_2436),
.A2(n_2435),
.B1(n_2149),
.B2(n_2123),
.C(n_2138),
.Y(n_2437)
);

AOI211xp5_ASAP7_75t_L g2438 ( 
.A1(n_2437),
.A2(n_2146),
.B(n_2150),
.C(n_2114),
.Y(n_2438)
);


endmodule