module fake_jpeg_7958_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_26),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_25),
.B1(n_10),
.B2(n_13),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_44),
.B(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_35),
.B1(n_33),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_23),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_17),
.B1(n_19),
.B2(n_1),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_19),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_32),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_30),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_38),
.C(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_35),
.B1(n_16),
.B2(n_30),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_39),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_61),
.C(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_51),
.C(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_69),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_58),
.B(n_53),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_63),
.C(n_66),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_44),
.B(n_36),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_8),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_17),
.Y(n_76)
);


endmodule