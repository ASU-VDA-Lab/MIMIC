module real_jpeg_20710_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_0),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_95),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_95),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_64),
.Y(n_275)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_85),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_85),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_85),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_5),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_91),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_252)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

BUFx3_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_9),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_97),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_97),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_236)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_11),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_12),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_12),
.B(n_29),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_16),
.B(n_45),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_100),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_12),
.A2(n_79),
.B1(n_80),
.B2(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_56),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_31),
.B(n_190),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_13),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_102),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_102),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_102),
.Y(n_159)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_31),
.A3(n_42),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_16),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_17),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_17),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_326),
.B(n_329),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_69),
.B(n_325),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_35),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_21),
.B(n_35),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_21),
.B(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_21),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_27),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_24),
.B(n_100),
.CON(n_99),
.SN(n_99)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_26),
.A2(n_29),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_26),
.A2(n_29),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_26),
.A2(n_29),
.B(n_33),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_31),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_28),
.A2(n_30),
.B1(n_99),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_30),
.B(n_100),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_65),
.C(n_67),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_36),
.A2(n_37),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.C(n_57),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_38),
.A2(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_38),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_38),
.A2(n_48),
.B1(n_295),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B(n_47),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_39),
.A2(n_44),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_39),
.A2(n_44),
.B1(n_84),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_39),
.A2(n_44),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_39),
.A2(n_44),
.B1(n_155),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_39),
.A2(n_44),
.B1(n_175),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_39),
.A2(n_44),
.B1(n_90),
.B2(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_39),
.A2(n_44),
.B1(n_86),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_39),
.A2(n_44),
.B1(n_229),
.B2(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_41),
.B(n_52),
.Y(n_185)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_42),
.A2(n_43),
.B(n_100),
.C(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_44),
.B(n_100),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_46),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_49),
.A2(n_50),
.B1(n_56),
.B2(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_55),
.B(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_50),
.A2(n_56),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_50),
.A2(n_56),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_54),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_54),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_51),
.A2(n_54),
.B1(n_129),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_51),
.A2(n_54),
.B1(n_110),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_51),
.A2(n_54),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_57),
.A2(n_58),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_62),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_59),
.A2(n_62),
.B1(n_108),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_59),
.A2(n_62),
.B1(n_236),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_322),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_67),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_318),
.B(n_324),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_287),
.A3(n_310),
.B1(n_316),
.B2(n_317),
.C(n_333),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_266),
.B(n_286),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_242),
.B(n_265),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_135),
.B(n_218),
.C(n_241),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_120),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_75),
.B(n_120),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_103),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_77),
.B(n_87),
.C(n_103),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_78),
.B(n_83),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_81),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_116),
.B1(n_119),
.B2(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_79),
.A2(n_80),
.B1(n_145),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_79),
.A2(n_80),
.B1(n_147),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_79),
.A2(n_80),
.B1(n_134),
.B2(n_177),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_79),
.A2(n_82),
.B1(n_119),
.B2(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_79),
.A2(n_117),
.B(n_227),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_80),
.B(n_100),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_98),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_105),
.B(n_111),
.C(n_112),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_142)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_132),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_131),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_217),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_212),
.B(n_216),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_198),
.B(n_211),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_179),
.B(n_197),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_167),
.B(n_178),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_156),
.B(n_166),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_148),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_161),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.C(n_176),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_187),
.B1(n_195),
.B2(n_196),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_194),
.C(n_195),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_199),
.B(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_208),
.C(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_240),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_230),
.B2(n_231),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_231),
.C(n_240),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_234),
.C(n_239),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_244),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_264),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_257),
.B2(n_258),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_258),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_252),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_256),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_260),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_278),
.B(n_281),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_268),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_284),
.B2(n_285),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_277),
.C(n_285),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B(n_276),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_289),
.C(n_300),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_289),
.B1(n_290),
.B2(n_315),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_276),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_302),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_296),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_304),
.C(n_309),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_301),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule