module fake_jpeg_12819_n_348 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_45),
.B(n_56),
.Y(n_103)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_10),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g87 ( 
.A(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_27),
.B(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_80),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_20),
.B1(n_40),
.B2(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_73),
.A2(n_75),
.B1(n_42),
.B2(n_39),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_81),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_40),
.B1(n_29),
.B2(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_41),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_21),
.B1(n_40),
.B2(n_43),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_109),
.B1(n_33),
.B2(n_23),
.Y(n_119)
);

INVx2_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_97),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_30),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_42),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_24),
.C(n_39),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_30),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_21),
.B1(n_43),
.B2(n_42),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_31),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_113),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_52),
.A2(n_21),
.B1(n_33),
.B2(n_26),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_46),
.A2(n_21),
.B1(n_38),
.B2(n_26),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_39),
.B1(n_23),
.B2(n_24),
.Y(n_125)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_0),
.B(n_2),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_37),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_43),
.B1(n_22),
.B2(n_31),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_136),
.B1(n_139),
.B2(n_99),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_124),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_125),
.A2(n_151),
.B1(n_113),
.B2(n_77),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_22),
.B1(n_42),
.B2(n_36),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_78),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_138),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_25),
.B1(n_36),
.B2(n_42),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_25),
.B1(n_37),
.B2(n_34),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_25),
.B1(n_37),
.B2(n_34),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_78),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_142),
.B(n_77),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_92),
.B1(n_70),
.B2(n_69),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_76),
.B(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_159),
.B(n_184),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_79),
.B1(n_98),
.B2(n_71),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_167),
.B1(n_178),
.B2(n_118),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_168),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_79),
.B1(n_98),
.B2(n_71),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_74),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_117),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_91),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_118),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_108),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_94),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_94),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_118),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_198),
.B1(n_219),
.B2(n_202),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_167),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_115),
.B(n_143),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_201),
.B(n_140),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_139),
.B1(n_119),
.B2(n_122),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_151),
.B1(n_130),
.B2(n_142),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_209),
.B1(n_214),
.B2(n_220),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_143),
.B(n_125),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_138),
.B1(n_125),
.B2(n_92),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_217),
.B(n_154),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_132),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_140),
.B1(n_174),
.B2(n_112),
.Y(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_126),
.B1(n_116),
.B2(n_123),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_116),
.B1(n_131),
.B2(n_123),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_121),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_216),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_118),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_150),
.B1(n_149),
.B2(n_135),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_179),
.A2(n_134),
.B1(n_100),
.B2(n_145),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_172),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_87),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_173),
.C(n_181),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_229),
.C(n_230),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_182),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_238),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_158),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_157),
.C(n_185),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_165),
.C(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_236),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_196),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_210),
.C(n_217),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_203),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_200),
.B1(n_209),
.B2(n_211),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_140),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_248),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_156),
.B1(n_189),
.B2(n_175),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_224),
.B1(n_231),
.B2(n_239),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_156),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_189),
.B(n_175),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_204),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_208),
.B(n_212),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_210),
.B(n_195),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_269),
.B1(n_271),
.B2(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_261),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_264),
.B1(n_237),
.B2(n_229),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_191),
.B1(n_198),
.B2(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_215),
.C(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_273),
.C(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_243),
.B(n_213),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_242),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_230),
.B(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_220),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_282),
.B1(n_288),
.B2(n_268),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_259),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_287),
.C(n_290),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_232),
.B1(n_235),
.B2(n_197),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_281),
.B(n_289),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_232),
.B1(n_238),
.B2(n_226),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_251),
.B1(n_233),
.B2(n_219),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_273),
.B1(n_255),
.B2(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_218),
.B1(n_207),
.B2(n_205),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g289 ( 
.A1(n_253),
.A2(n_250),
.B(n_207),
.C(n_174),
.D(n_87),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_197),
.C(n_161),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_247),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_291),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_276),
.B1(n_275),
.B2(n_281),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_297),
.B1(n_298),
.B2(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_274),
.B1(n_291),
.B2(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_258),
.B1(n_260),
.B2(n_255),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_252),
.C(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_265),
.C(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_254),
.C(n_267),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_263),
.B1(n_267),
.B2(n_245),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_311),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_282),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_289),
.B(n_285),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_284),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_169),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_163),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_299),
.C(n_298),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_304),
.B1(n_297),
.B2(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_263),
.B1(n_177),
.B2(n_161),
.Y(n_318)
);

A2O1A1O1Ixp25_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_307),
.B(n_315),
.C(n_317),
.D(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_327),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_110),
.Y(n_333)
);

OAI221xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_300),
.B1(n_295),
.B2(n_303),
.C(n_305),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_87),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_100),
.B1(n_70),
.B2(n_93),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_311),
.C(n_318),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_309),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_324),
.C(n_92),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_110),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_101),
.B1(n_7),
.B2(n_11),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_335),
.B(n_321),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_323),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_337),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_331),
.Y(n_343)
);

NAND2x1_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_340),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_344),
.Y(n_345)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_344),
.A3(n_341),
.B1(n_342),
.B2(n_328),
.C1(n_333),
.C2(n_334),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_14),
.B(n_15),
.Y(n_348)
);


endmodule