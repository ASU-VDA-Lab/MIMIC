module fake_jpeg_7493_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_45),
.Y(n_47)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_46),
.B(n_33),
.C(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_31),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_23),
.C(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_73),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_64),
.Y(n_105)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_67),
.B1(n_38),
.B2(n_68),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_9),
.C(n_16),
.Y(n_93)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_28),
.B1(n_17),
.B2(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_34),
.B1(n_33),
.B2(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_20),
.B1(n_18),
.B2(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_34),
.B1(n_33),
.B2(n_22),
.Y(n_74)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_46),
.B(n_42),
.C(n_38),
.D(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_12),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_78),
.B(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_90),
.B1(n_103),
.B2(n_107),
.Y(n_112)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_18),
.B(n_15),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_45),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_97),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_1),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_101),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_20),
.A3(n_9),
.B1(n_10),
.B2(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_104),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_15),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_61),
.B1(n_53),
.B2(n_49),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_1),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_59),
.A2(n_72),
.B1(n_58),
.B2(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_14),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_50),
.B(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_71),
.B1(n_51),
.B2(n_58),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_119),
.B1(n_131),
.B2(n_77),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_109),
.B1(n_102),
.B2(n_95),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_122),
.B1(n_137),
.B2(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_61),
.B1(n_53),
.B2(n_12),
.Y(n_122)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_3),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_80),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_93),
.B(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_141),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_86),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_146),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_76),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_92),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_92),
.C(n_105),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_170),
.Y(n_176)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_100),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_148),
.A2(n_158),
.B(n_161),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_154),
.B1(n_156),
.B2(n_168),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_138),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_155),
.B(n_173),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_77),
.B(n_97),
.C(n_94),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_82),
.B1(n_98),
.B2(n_96),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_106),
.B(n_75),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_4),
.B(n_5),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_114),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_114),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_96),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_111),
.B1(n_89),
.B2(n_87),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_111),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_91),
.C(n_106),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_5),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_5),
.B(n_6),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_6),
.B(n_7),
.Y(n_199)
);

NAND2x1p5_ASAP7_75t_R g173 ( 
.A(n_131),
.B(n_5),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_178),
.B(n_186),
.Y(n_223)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_140),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_182),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_116),
.B1(n_117),
.B2(n_122),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_185),
.B(n_194),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_117),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_133),
.B(n_132),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_116),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_143),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_114),
.B1(n_115),
.B2(n_129),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_164),
.B1(n_145),
.B2(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_153),
.B1(n_161),
.B2(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_6),
.B(n_8),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_146),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_141),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_113),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_135),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_158),
.B(n_153),
.C(n_155),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_213),
.B(n_216),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_142),
.B1(n_151),
.B2(n_168),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_179),
.B1(n_201),
.B2(n_192),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_195),
.B1(n_202),
.B2(n_188),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_155),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_113),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_155),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_186),
.B(n_200),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_166),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_226),
.A2(n_228),
.B1(n_180),
.B2(n_181),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_200),
.B1(n_174),
.B2(n_178),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_157),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_176),
.C(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_6),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_210),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_176),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_190),
.B1(n_194),
.B2(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_180),
.C(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_248),
.C(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_206),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_249),
.A2(n_207),
.B1(n_217),
.B2(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_215),
.A2(n_181),
.B1(n_182),
.B2(n_179),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_199),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_203),
.B1(n_124),
.B2(n_130),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_203),
.C(n_124),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.C(n_233),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_106),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_268),
.B1(n_208),
.B2(n_247),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_252),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_269),
.C(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_223),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_216),
.B1(n_224),
.B2(n_208),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_233),
.C(n_220),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_245),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_274),
.B(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_212),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_241),
.A2(n_216),
.B(n_208),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_279),
.C(n_284),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_287),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_237),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_222),
.B1(n_243),
.B2(n_232),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_250),
.A3(n_283),
.B1(n_265),
.B2(n_243),
.C1(n_239),
.C2(n_262),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_248),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_244),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_286),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_254),
.C(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_260),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_297),
.Y(n_310)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_257),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_272),
.B1(n_271),
.B2(n_274),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_265),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_208),
.B(n_231),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_264),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_250),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_293),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_299),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_287),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_311),
.B(n_299),
.Y(n_312)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_290),
.A3(n_286),
.B(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_268),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_312),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_317),
.A3(n_306),
.B1(n_304),
.B2(n_314),
.C1(n_292),
.C2(n_275),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_316),
.B(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_293),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_285),
.A3(n_263),
.B1(n_284),
.B2(n_259),
.C1(n_279),
.C2(n_255),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_10),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

AOI321xp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_323),
.A3(n_319),
.B1(n_322),
.B2(n_11),
.C(n_8),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_8),
.Y(n_327)
);


endmodule