module real_jpeg_24612_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_288;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_215;
wire n_286;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_30),
.B1(n_56),
.B2(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_30),
.B1(n_51),
.B2(n_109),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_2),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_27),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_27),
.B1(n_56),
.B2(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_59),
.B(n_65),
.C(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_55),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_4),
.A2(n_60),
.B(n_74),
.C(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_26),
.C(n_37),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_4),
.B(n_130),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_11),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_4),
.B(n_35),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_41),
.B1(n_56),
.B2(n_60),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_278),
.B1(n_291),
.B2(n_292),
.Y(n_13)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_14),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_134),
.B(n_277),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_111),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_16),
.B(n_111),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_91),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_17),
.B(n_82),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_18),
.B(n_47),
.C(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_19),
.B(n_33),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_20),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx3_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_31),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_24),
.B(n_31),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_26),
.B(n_233),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_27),
.A2(n_39),
.B(n_75),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_28),
.A2(n_95),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_28),
.B(n_225),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_29),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_31),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_31),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B(n_42),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_34),
.B(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_34),
.A2(n_88),
.B(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_35),
.B(n_195),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_38),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_40),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_40),
.B(n_208),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_42),
.B(n_205),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_43),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_43),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_69),
.B2(n_70),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_61),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_50),
.B(n_66),
.Y(n_144)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_62),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_55),
.B(n_108),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_71),
.B(n_156),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_71),
.A2(n_78),
.B(n_129),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_72),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_79),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_104),
.Y(n_158)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_77),
.B(n_149),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_79),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_90),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_83),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_83),
.A2(n_90),
.B1(n_190),
.B2(n_249),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_83),
.A2(n_115),
.B(n_117),
.Y(n_288)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_89),
.B(n_194),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_91),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_103),
.C(n_105),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_92),
.A2(n_93),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_100),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_97),
.B(n_218),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_101),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_103),
.A2(n_105),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_103),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_105),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_133),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_122),
.B2(n_123),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_113),
.B(n_123),
.C(n_133),
.Y(n_289)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_128),
.B(n_132),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_148),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_132),
.B(n_281),
.CI(n_288),
.CON(n_280),
.SN(n_280)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_272),
.B(n_276),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_183),
.B(n_258),
.C(n_271),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_171),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_137),
.B(n_171),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_153),
.B2(n_170),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_151),
.B2(n_152),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_140),
.B(n_152),
.C(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_143),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_144),
.B(n_160),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_145),
.A2(n_146),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_155),
.B(n_162),
.C(n_163),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.C(n_178),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_173),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_181),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_257),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_199),
.B(n_256),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_186),
.B(n_196),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_192),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_187),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_189),
.B(n_192),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_190),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_251),
.B(n_255),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_242),
.B(n_250),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_222),
.B(n_241),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_221),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_212),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_215),
.C(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_230),
.B(n_240),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_236),
.B(n_239),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_247),
.C(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_270),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_268),
.B2(n_269),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_269),
.C(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_290),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_289),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_280),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);


endmodule