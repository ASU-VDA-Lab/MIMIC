module fake_netlist_6_3054_n_2293 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_192, n_57, n_169, n_51, n_649, n_283, n_2293);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2293;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_907;
wire n_1446;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_687;
wire n_697;
wire n_890;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_682;
wire n_851;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_2292;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2016;
wire n_1905;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_1270;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g674 ( 
.A(n_17),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_30),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_588),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_311),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_642),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_96),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_604),
.Y(n_681)
);

BUFx5_ASAP7_75t_L g682 ( 
.A(n_483),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_143),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_146),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_653),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_606),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_548),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_338),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_191),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_154),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_647),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_498),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_641),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_636),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_449),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_398),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_89),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_522),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_165),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_651),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_232),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_31),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_459),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_471),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_328),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_7),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_625),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_509),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_19),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_38),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_393),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_193),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_646),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_639),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_621),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_174),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_623),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_635),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_628),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_121),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_350),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_73),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_466),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_74),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_279),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_118),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_644),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_45),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_649),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_63),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_345),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_301),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_319),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_574),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_187),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_631),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_103),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_476),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_633),
.Y(n_740)
);

BUFx2_ASAP7_75t_SL g741 ( 
.A(n_376),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_440),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_114),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_400),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_74),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_374),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_45),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_67),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_531),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_559),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_629),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_47),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_139),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_176),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_637),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_2),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_230),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_668),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_6),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_643),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_76),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_267),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_26),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_632),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_542),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_467),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_92),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_304),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_461),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_663),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_655),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_0),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_61),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_364),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_381),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_75),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_60),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_190),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_252),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_640),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_638),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_101),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_526),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_2),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_173),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_275),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_626),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_624),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_652),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_545),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_455),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_474),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_383),
.Y(n_793)
);

BUFx8_ASAP7_75t_SL g794 ( 
.A(n_520),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_204),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_657),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_645),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_427),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_243),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_418),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_654),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_235),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_593),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_318),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_55),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_310),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_656),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_505),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_525),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_339),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_295),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_445),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_341),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_630),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_506),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_549),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_514),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_650),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_323),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_15),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_305),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_86),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_300),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_297),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_0),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_48),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_565),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_205),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_291),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_524),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_124),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_290),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_44),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_127),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_616),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_550),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_622),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_124),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_453),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_113),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_239),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_77),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_268),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_206),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_214),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_362),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_166),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_479),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_627),
.Y(n_849)
);

INVxp33_ASAP7_75t_L g850 ( 
.A(n_674),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_831),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_831),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_831),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_690),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_675),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_683),
.Y(n_856)
);

CKINVDCx14_ASAP7_75t_R g857 ( 
.A(n_840),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_794),
.Y(n_858)
);

CKINVDCx16_ASAP7_75t_R g859 ( 
.A(n_824),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_682),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_710),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_711),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_721),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_761),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_723),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_682),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_707),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_729),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_698),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_738),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_743),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_763),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_767),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_776),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_677),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_682),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_784),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_680),
.Y(n_879)
);

INVxp33_ASAP7_75t_L g880 ( 
.A(n_805),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_728),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_820),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_750),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_833),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_679),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_834),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_687),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_682),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_678),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_693),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_696),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_689),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_695),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_712),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_719),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_681),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_720),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_726),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_736),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_756),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_739),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_740),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_685),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_755),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_700),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_757),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_697),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_686),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_705),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_691),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_682),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_699),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_751),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_762),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_764),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_765),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_779),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_730),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_733),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_780),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_701),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_783),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_751),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_786),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_688),
.B(n_1),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_793),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_803),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_808),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_749),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_819),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_823),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_702),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_792),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_760),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_837),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_839),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_845),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_798),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_692),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_676),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_725),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_703),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_694),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_718),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_706),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_802),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_727),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_813),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_827),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_835),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_870),
.A2(n_881),
.B1(n_859),
.B2(n_865),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_851),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_889),
.B(n_942),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_852),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_853),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_913),
.B(n_847),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_855),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_896),
.B(n_903),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_856),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_923),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_883),
.B(n_704),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_941),
.B(n_770),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_862),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_863),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_908),
.B(n_843),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_887),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_865),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_890),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_864),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_891),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_894),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_879),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_933),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_857),
.B(n_766),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_866),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_869),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_871),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_854),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_938),
.B(n_766),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_907),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_872),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_910),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_873),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_858),
.B(n_737),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_874),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_875),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_878),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_882),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_912),
.B(n_787),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_868),
.A2(n_782),
.B1(n_745),
.B2(n_747),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_884),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_932),
.B(n_832),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_886),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_925),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_861),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_921),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_941),
.B(n_811),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_895),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_897),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_945),
.B(n_828),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_898),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_899),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_925),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_940),
.B(n_829),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_901),
.B(n_830),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_902),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_904),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_947),
.B(n_708),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_906),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_914),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_915),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_916),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_850),
.B(n_709),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_917),
.B(n_836),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_905),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_939),
.Y(n_1016)
);

OA21x2_ASAP7_75t_L g1017 ( 
.A1(n_920),
.A2(n_924),
.B(n_922),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_867),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_926),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_927),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_943),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_944),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_R g1023 ( 
.A1(n_876),
.A2(n_773),
.B1(n_838),
.B2(n_753),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_877),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_928),
.B(n_841),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_930),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_931),
.B(n_713),
.Y(n_1027)
);

CKINVDCx11_ASAP7_75t_R g1028 ( 
.A(n_868),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_888),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_935),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_936),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_937),
.B(n_849),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_911),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_918),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_946),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_948),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_1015),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_994),
.B(n_949),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_989),
.B(n_934),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1018),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_994),
.B(n_950),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_967),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1018),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1029),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_1013),
.Y(n_1045)
);

INVx8_ASAP7_75t_L g1046 ( 
.A(n_1034),
.Y(n_1046)
);

BUFx10_ASAP7_75t_L g1047 ( 
.A(n_953),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_1029),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1033),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1003),
.B(n_715),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_973),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_1008),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_966),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_1033),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_1003),
.B(n_716),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_952),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_968),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_952),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_970),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_955),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_971),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_998),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1016),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_975),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1021),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_965),
.B(n_880),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_999),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1022),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_960),
.B(n_717),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1000),
.B(n_885),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1035),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_957),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_L g1073 ( 
.A(n_1005),
.B(n_676),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_960),
.B(n_722),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_982),
.B(n_909),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_959),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_960),
.B(n_724),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_979),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1014),
.B(n_714),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1001),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_975),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1002),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_963),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1006),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_964),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_976),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_983),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_SL g1088 ( 
.A(n_990),
.B(n_731),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1009),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_L g1090 ( 
.A(n_1032),
.B(n_676),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1010),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_958),
.B(n_1004),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_961),
.B(n_732),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_977),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_980),
.B(n_892),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_978),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_996),
.B(n_893),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_985),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1017),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_951),
.B(n_919),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1025),
.B(n_778),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1012),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_993),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_995),
.A2(n_741),
.B(n_900),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1036),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1019),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1020),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_995),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1024),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1024),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_962),
.B(n_742),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_983),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_997),
.B(n_734),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_986),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_SL g1115 ( 
.A(n_974),
.B(n_748),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_986),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_988),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_SL g1118 ( 
.A(n_956),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_988),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1026),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_992),
.B(n_746),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_SL g1122 ( 
.A(n_1027),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_972),
.B(n_900),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_954),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1011),
.B(n_860),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_954),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1017),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1031),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_1023),
.A2(n_860),
.B1(n_10),
.B2(n_18),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1030),
.Y(n_1130)
);

XNOR2xp5_ASAP7_75t_L g1131 ( 
.A(n_1037),
.B(n_929),
.Y(n_1131)
);

INVxp33_ASAP7_75t_L g1132 ( 
.A(n_1042),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1099),
.A2(n_984),
.B(n_981),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1053),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1057),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1059),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1061),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1108),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1062),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1109),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1066),
.B(n_1007),
.Y(n_1141)
);

INVxp33_ASAP7_75t_L g1142 ( 
.A(n_1042),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1067),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1092),
.B(n_969),
.Y(n_1144)
);

XOR2xp5_ASAP7_75t_L g1145 ( 
.A(n_1045),
.B(n_1028),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1080),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1082),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1081),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1048),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1123),
.B(n_969),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1048),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1084),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1089),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1091),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1102),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1106),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1107),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1038),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_SL g1159 ( 
.A(n_1039),
.B(n_735),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1041),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1130),
.Y(n_1161)
);

NOR2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1125),
.B(n_752),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1076),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1083),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1099),
.A2(n_981),
.B(n_987),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1078),
.B(n_991),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1045),
.B(n_759),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1127),
.B(n_744),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1085),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1127),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1128),
.B(n_772),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1052),
.B(n_777),
.Y(n_1173)
);

INVxp33_ASAP7_75t_L g1174 ( 
.A(n_1095),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1086),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1110),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1094),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1098),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1079),
.A2(n_758),
.B(n_754),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1070),
.B(n_822),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1103),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1048),
.Y(n_1182)
);

XNOR2xp5_ASAP7_75t_L g1183 ( 
.A(n_1101),
.B(n_768),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1124),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_1046),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1126),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1120),
.B(n_825),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1063),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1096),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1050),
.B(n_826),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1065),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_1046),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1068),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1055),
.B(n_842),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1047),
.B(n_769),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_1075),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1113),
.B(n_1),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1071),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1051),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1105),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1060),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1040),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1047),
.B(n_771),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1043),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1117),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1044),
.Y(n_1206)
);

XOR2xp5_ASAP7_75t_L g1207 ( 
.A(n_1121),
.B(n_774),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1049),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1127),
.B(n_775),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1112),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1114),
.B(n_781),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1119),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1100),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1056),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1058),
.Y(n_1215)
);

INVxp33_ASAP7_75t_SL g1216 ( 
.A(n_1097),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1104),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1093),
.B(n_785),
.Y(n_1220)
);

XNOR2xp5_ASAP7_75t_L g1221 ( 
.A(n_1129),
.B(n_788),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1064),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1064),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1064),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1087),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1087),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1087),
.Y(n_1227)
);

XNOR2x2_ASAP7_75t_L g1228 ( 
.A(n_1129),
.B(n_3),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1116),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1188),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1189),
.Y(n_1231)
);

NOR3x1_ASAP7_75t_L g1232 ( 
.A(n_1228),
.B(n_1150),
.C(n_1197),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_SL g1233 ( 
.A(n_1205),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1144),
.B(n_1111),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1211),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1158),
.B(n_1116),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1160),
.B(n_1171),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1180),
.B(n_1134),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1213),
.B(n_1174),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1132),
.B(n_1115),
.Y(n_1240)
);

BUFx4_ASAP7_75t_L g1241 ( 
.A(n_1185),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1172),
.Y(n_1242)
);

AND2x2_ASAP7_75t_SL g1243 ( 
.A(n_1196),
.B(n_1073),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1192),
.B(n_1088),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_1090),
.B1(n_848),
.B2(n_1122),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1186),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1136),
.B(n_1116),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1190),
.A2(n_1074),
.B(n_1077),
.C(n_1069),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1138),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1142),
.B(n_789),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1137),
.B(n_790),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1139),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1159),
.B(n_1173),
.C(n_1168),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1133),
.B(n_791),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1143),
.B(n_795),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1146),
.B(n_796),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1216),
.A2(n_1118),
.B1(n_848),
.B2(n_799),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1141),
.A2(n_800),
.B1(n_801),
.B2(n_797),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1217),
.B(n_1149),
.Y(n_1259)
);

AND3x1_ASAP7_75t_L g1260 ( 
.A(n_1187),
.B(n_3),
.C(n_4),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1147),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1149),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1195),
.B(n_804),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1203),
.B(n_806),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1152),
.B(n_807),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1153),
.A2(n_848),
.B1(n_810),
.B2(n_812),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1194),
.A2(n_814),
.B1(n_815),
.B2(n_809),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1154),
.B(n_816),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1155),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1156),
.B(n_817),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1140),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1157),
.A2(n_821),
.B1(n_844),
.B2(n_818),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1184),
.A2(n_846),
.B1(n_156),
.B2(n_157),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1169),
.B(n_4),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1163),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1167),
.B(n_155),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1162),
.B(n_5),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1183),
.B(n_5),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1149),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1209),
.B(n_6),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1220),
.B(n_158),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1207),
.B(n_7),
.C(n_8),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1166),
.B(n_8),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1148),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1179),
.B(n_159),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1210),
.B(n_9),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1199),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1151),
.B(n_160),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1164),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1161),
.B(n_9),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1218),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1176),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1151),
.B(n_161),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1165),
.B(n_11),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1151),
.B(n_162),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1200),
.A2(n_164),
.B1(n_167),
.B2(n_163),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1212),
.B(n_12),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1170),
.A2(n_169),
.B1(n_170),
.B2(n_168),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1175),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_L g1300 ( 
.A(n_1182),
.B(n_171),
.Y(n_1300)
);

NOR2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1214),
.B(n_1215),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1177),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1219),
.A2(n_1181),
.B1(n_1191),
.B2(n_1178),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1193),
.B(n_13),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1198),
.B(n_13),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1201),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1202),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1206),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1182),
.B(n_14),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1231),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1238),
.B(n_1182),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1259),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1252),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1261),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1259),
.B(n_1204),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_SL g1316 ( 
.A(n_1263),
.B(n_1145),
.C(n_1208),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1253),
.B(n_1131),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1234),
.B(n_1222),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1244),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1262),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1262),
.B(n_1227),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1235),
.B(n_1229),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1262),
.Y(n_1323)
);

INVx5_ASAP7_75t_L g1324 ( 
.A(n_1279),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1269),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1239),
.B(n_1221),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1284),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1233),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1277),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1309),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1240),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1242),
.B(n_1223),
.Y(n_1332)
);

NAND3xp33_ASAP7_75t_L g1333 ( 
.A(n_1278),
.B(n_1225),
.C(n_1224),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1230),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1287),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1279),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1237),
.B(n_1226),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1301),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1275),
.B(n_172),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1246),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1289),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1264),
.B(n_175),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1249),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1306),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1271),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1308),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1299),
.B(n_177),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1302),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1285),
.A2(n_1283),
.B1(n_1274),
.B2(n_1280),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1307),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1232),
.B(n_178),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1286),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1282),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1247),
.B(n_179),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1297),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1243),
.B(n_180),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1294),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1304),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1236),
.B(n_16),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1251),
.B(n_17),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1248),
.B(n_1255),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1305),
.Y(n_1363)
);

OR2x4_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_18),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1256),
.B(n_19),
.Y(n_1365)
);

INVx5_ASAP7_75t_L g1366 ( 
.A(n_1233),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1250),
.B(n_1265),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1260),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1241),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1303),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1257),
.Y(n_1371)
);

CKINVDCx8_ASAP7_75t_R g1372 ( 
.A(n_1300),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_R g1374 ( 
.A(n_1270),
.B(n_181),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1288),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1258),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1293),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1295),
.Y(n_1378)
);

XNOR2xp5_ASAP7_75t_L g1379 ( 
.A(n_1245),
.B(n_20),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1291),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1380)
);

CKINVDCx8_ASAP7_75t_R g1381 ( 
.A(n_1281),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1276),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1254),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1273),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1342),
.A2(n_1267),
.B(n_1296),
.C(n_1298),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1331),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1359),
.B(n_1272),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1353),
.A2(n_1266),
.B1(n_23),
.B2(n_21),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1362),
.A2(n_183),
.B(n_182),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1356),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1310),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1311),
.A2(n_185),
.B(n_184),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1350),
.A2(n_188),
.B(n_186),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1318),
.A2(n_192),
.B(n_189),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1313),
.Y(n_1395)
);

INVx3_ASAP7_75t_SL g1396 ( 
.A(n_1328),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1356),
.B(n_24),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1370),
.A2(n_195),
.A3(n_196),
.B(n_194),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1326),
.B(n_25),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1366),
.B(n_198),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1382),
.A2(n_199),
.B(n_197),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1383),
.A2(n_201),
.B(n_200),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1338),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1361),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1377),
.A2(n_203),
.B(n_202),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1330),
.B(n_27),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1314),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1384),
.A2(n_208),
.B(n_207),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1368),
.B(n_28),
.Y(n_1411)
);

O2A1O1Ixp5_ASAP7_75t_L g1412 ( 
.A1(n_1360),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1365),
.A2(n_210),
.B(n_209),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1335),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1325),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1337),
.A2(n_212),
.B(n_211),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1375),
.A2(n_215),
.B(n_213),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1367),
.A2(n_217),
.B(n_216),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1378),
.A2(n_219),
.B(n_218),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_221),
.B(n_220),
.Y(n_1420)
);

BUFx4f_ASAP7_75t_SL g1421 ( 
.A(n_1369),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1330),
.B(n_29),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1351),
.A2(n_223),
.B(n_222),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1341),
.B(n_31),
.Y(n_1424)
);

NAND2x1_ASAP7_75t_L g1425 ( 
.A(n_1323),
.B(n_1320),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1344),
.B(n_32),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1366),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1347),
.B(n_32),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1357),
.A2(n_225),
.B(n_224),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1376),
.B(n_33),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1317),
.A2(n_227),
.B(n_226),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1348),
.A2(n_229),
.B(n_228),
.Y(n_1432)
);

AO21x1_ASAP7_75t_L g1433 ( 
.A1(n_1355),
.A2(n_35),
.B(n_34),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_SL g1434 ( 
.A(n_1319),
.B(n_231),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1333),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1366),
.B(n_238),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1334),
.A2(n_1343),
.B(n_1340),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1321),
.A2(n_234),
.B(n_233),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1345),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1346),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1312),
.B(n_236),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1332),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_SL g1443 ( 
.A1(n_1380),
.A2(n_240),
.B(n_237),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1316),
.A2(n_1354),
.B(n_1381),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1324),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1324),
.A2(n_242),
.B(n_241),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1323),
.Y(n_1447)
);

INVx5_ASAP7_75t_L g1448 ( 
.A(n_1320),
.Y(n_1448)
);

BUFx4f_ASAP7_75t_L g1449 ( 
.A(n_1327),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1339),
.A2(n_245),
.B(n_244),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1324),
.A2(n_247),
.B(n_246),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1372),
.A2(n_249),
.B(n_248),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1329),
.B(n_36),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1336),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1379),
.A2(n_251),
.B(n_250),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1327),
.B(n_257),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1315),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1352),
.B(n_36),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1374),
.B(n_37),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1322),
.A2(n_254),
.B(n_253),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1364),
.B(n_37),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1315),
.A2(n_256),
.B(n_255),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1322),
.Y(n_1463)
);

AO21x1_ASAP7_75t_L g1464 ( 
.A1(n_1379),
.A2(n_40),
.B(n_39),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1458),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1393),
.A2(n_662),
.B(n_661),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1416),
.A2(n_259),
.B(n_258),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1395),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_SL g1469 ( 
.A(n_1427),
.B(n_41),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1388),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1399),
.B(n_42),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1385),
.A2(n_47),
.B(n_43),
.C(n_46),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1389),
.A2(n_261),
.B(n_260),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1449),
.Y(n_1474)
);

NOR3xp33_ASAP7_75t_L g1475 ( 
.A(n_1459),
.B(n_1444),
.C(n_1406),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1404),
.B(n_46),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1420),
.A2(n_1423),
.B(n_1410),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1430),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1450),
.A2(n_263),
.B(n_262),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1415),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1387),
.A2(n_265),
.B(n_264),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1437),
.A2(n_269),
.B(n_266),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1394),
.A2(n_271),
.B(n_270),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_273),
.B(n_272),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1409),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1391),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1442),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_1457),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1440),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1439),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1407),
.A2(n_276),
.B(n_274),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1402),
.A2(n_278),
.B(n_277),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_SL g1493 ( 
.A(n_1464),
.B(n_51),
.C(n_52),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1417),
.A2(n_281),
.B(n_280),
.Y(n_1494)
);

AO31x2_ASAP7_75t_L g1495 ( 
.A1(n_1433),
.A2(n_283),
.A3(n_284),
.B(n_282),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1392),
.A2(n_1451),
.B(n_1438),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1419),
.A2(n_1403),
.B(n_1432),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1424),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_SL g1499 ( 
.A1(n_1435),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1426),
.Y(n_1500)
);

AOI221x1_ASAP7_75t_L g1501 ( 
.A1(n_1390),
.A2(n_1413),
.B1(n_1455),
.B2(n_1431),
.C(n_1443),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1460),
.A2(n_1452),
.B(n_1446),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1462),
.A2(n_286),
.B(n_285),
.Y(n_1503)
);

AO31x2_ASAP7_75t_L g1504 ( 
.A1(n_1429),
.A2(n_1428),
.A3(n_1463),
.B(n_1445),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1441),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1412),
.A2(n_56),
.B(n_53),
.C(n_54),
.Y(n_1506)
);

INVx8_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1386),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_SL g1509 ( 
.A(n_1405),
.B(n_56),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1401),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1396),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1448),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1421),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1434),
.A2(n_673),
.B(n_288),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1400),
.A2(n_672),
.B(n_289),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1436),
.A2(n_671),
.B(n_292),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1456),
.A2(n_293),
.B(n_287),
.Y(n_1517)
);

AO31x2_ASAP7_75t_L g1518 ( 
.A1(n_1447),
.A2(n_296),
.A3(n_298),
.B(n_294),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1425),
.A2(n_302),
.B(n_299),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1408),
.A2(n_306),
.B(n_303),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1461),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1521)
);

AO31x2_ASAP7_75t_L g1522 ( 
.A1(n_1398),
.A2(n_308),
.A3(n_309),
.B(n_307),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1454),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1441),
.A2(n_313),
.B(n_312),
.Y(n_1524)
);

AOI21xp33_ASAP7_75t_L g1525 ( 
.A1(n_1414),
.A2(n_60),
.B(n_61),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1448),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1422),
.A2(n_315),
.B(n_314),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1453),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1455),
.A2(n_317),
.B(n_316),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_R g1530 ( 
.A(n_1411),
.B(n_1397),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1398),
.A2(n_321),
.B(n_320),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1399),
.B(n_62),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1457),
.B(n_322),
.Y(n_1533)
);

O2A1O1Ixp5_ASAP7_75t_L g1534 ( 
.A1(n_1393),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1430),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1401),
.B(n_324),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1393),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1395),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_SL g1539 ( 
.A1(n_1393),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1396),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1385),
.A2(n_71),
.B(n_72),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1393),
.A2(n_670),
.B(n_326),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1393),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1386),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1442),
.B(n_75),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1404),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1404),
.B(n_78),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1395),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1449),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1395),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1389),
.A2(n_327),
.B(n_325),
.Y(n_1551)
);

AO31x2_ASAP7_75t_L g1552 ( 
.A1(n_1433),
.A2(n_330),
.A3(n_331),
.B(n_329),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1389),
.A2(n_333),
.B(n_332),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1395),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1395),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1393),
.A2(n_335),
.B(n_334),
.Y(n_1556)
);

AO21x2_ASAP7_75t_L g1557 ( 
.A1(n_1393),
.A2(n_337),
.B(n_336),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1393),
.A2(n_669),
.B(n_342),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1449),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1393),
.A2(n_667),
.B(n_343),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1406),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1561)
);

AO31x2_ASAP7_75t_L g1562 ( 
.A1(n_1433),
.A2(n_344),
.A3(n_346),
.B(n_340),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1401),
.B(n_347),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1393),
.A2(n_666),
.B(n_349),
.Y(n_1564)
);

AOI221x1_ASAP7_75t_L g1565 ( 
.A1(n_1406),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_SL g1566 ( 
.A1(n_1393),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_SL g1567 ( 
.A1(n_1393),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1391),
.B(n_348),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1395),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1393),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1399),
.B(n_87),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1399),
.B(n_88),
.Y(n_1572)
);

AO31x2_ASAP7_75t_L g1573 ( 
.A1(n_1433),
.A2(n_352),
.A3(n_353),
.B(n_351),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1414),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1437),
.A2(n_355),
.B(n_354),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1395),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1508),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1485),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1480),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_356),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1511),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1489),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1541),
.A2(n_1477),
.B1(n_1563),
.B2(n_1536),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1468),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1548),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1465),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1587)
);

CKINVDCx6p67_ASAP7_75t_R g1588 ( 
.A(n_1526),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1523),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1498),
.B(n_90),
.Y(n_1590)
);

CKINVDCx16_ASAP7_75t_R g1591 ( 
.A(n_1488),
.Y(n_1591)
);

BUFx4f_ASAP7_75t_SL g1592 ( 
.A(n_1505),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1474),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1540),
.Y(n_1594)
);

BUFx8_ASAP7_75t_SL g1595 ( 
.A(n_1513),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1574),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1507),
.Y(n_1597)
);

BUFx10_ASAP7_75t_L g1598 ( 
.A(n_1533),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1545),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1479),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1507),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1500),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1475),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1550),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1466),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1555),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1576),
.Y(n_1607)
);

BUFx10_ASAP7_75t_L g1608 ( 
.A(n_1549),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1493),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1509),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1470),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1535),
.A2(n_105),
.B1(n_102),
.B2(n_104),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1538),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1542),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1554),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1546),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1616)
);

BUFx2_ASAP7_75t_R g1617 ( 
.A(n_1512),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1558),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1559),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1569),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1490),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1504),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1537),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1560),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1624)
);

AOI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1561),
.A2(n_112),
.B(n_113),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1564),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1530),
.Y(n_1627)
);

CKINVDCx16_ASAP7_75t_R g1628 ( 
.A(n_1471),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1557),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1486),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1467),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1631)
);

CKINVDCx11_ASAP7_75t_R g1632 ( 
.A(n_1487),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1532),
.B(n_357),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1504),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1476),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1571),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1547),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1469),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1525),
.A2(n_1572),
.B1(n_1529),
.B2(n_1556),
.Y(n_1639)
);

INVx6_ASAP7_75t_L g1640 ( 
.A(n_1568),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1481),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1524),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1515),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1521),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1517),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1543),
.A2(n_1570),
.B(n_1565),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1501),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_1647)
);

CKINVDCx20_ASAP7_75t_R g1648 ( 
.A(n_1514),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1522),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1483),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1522),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1518),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1516),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1499),
.B(n_125),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1519),
.B(n_358),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1484),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1482),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1510),
.Y(n_1658)
);

BUFx4f_ASAP7_75t_SL g1659 ( 
.A(n_1520),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1518),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1497),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1495),
.Y(n_1662)
);

CKINVDCx11_ASAP7_75t_R g1663 ( 
.A(n_1478),
.Y(n_1663)
);

BUFx8_ASAP7_75t_L g1664 ( 
.A(n_1528),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1527),
.Y(n_1665)
);

INVx6_ASAP7_75t_L g1666 ( 
.A(n_1472),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1503),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1495),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1506),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1531),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1552),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1502),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1575),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1552),
.Y(n_1674)
);

CKINVDCx20_ASAP7_75t_R g1675 ( 
.A(n_1539),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_SL g1676 ( 
.A(n_1566),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1578),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1585),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1582),
.Y(n_1679)
);

CKINVDCx16_ASAP7_75t_R g1680 ( 
.A(n_1591),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1601),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1673),
.A2(n_1496),
.B(n_1473),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1577),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1594),
.B(n_359),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1583),
.A2(n_1567),
.B(n_1534),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1589),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1586),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1604),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1606),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1630),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1607),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1620),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1622),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1615),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1596),
.B(n_133),
.Y(n_1695)
);

AOI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1652),
.A2(n_1660),
.B(n_1651),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1595),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1579),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1613),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1635),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1649),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1663),
.A2(n_1494),
.B1(n_1492),
.B2(n_1491),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1621),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1630),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1581),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1634),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1657),
.A2(n_1553),
.B(n_1551),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1637),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1668),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1671),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1584),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1593),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1644),
.A2(n_1573),
.B1(n_1562),
.B2(n_136),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1645),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1665),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1590),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_SL g1719 ( 
.A(n_1619),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1628),
.B(n_1562),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1667),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1654),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1676),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1667),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1659),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1667),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1658),
.A2(n_1573),
.B1(n_136),
.B2(n_134),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1630),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1639),
.A2(n_1625),
.B(n_1641),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1597),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1666),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1640),
.Y(n_1732)
);

AO21x1_ASAP7_75t_SL g1733 ( 
.A1(n_1603),
.A2(n_135),
.B(n_137),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1666),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1636),
.B(n_135),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1640),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1675),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1647),
.A2(n_1646),
.B(n_1587),
.C(n_1623),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1608),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1655),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1597),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1650),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1633),
.B(n_137),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1588),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1598),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1653),
.B(n_138),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1599),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1643),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1648),
.A2(n_361),
.B(n_360),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1602),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1670),
.A2(n_365),
.B(n_363),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1580),
.B(n_366),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1617),
.B(n_138),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1664),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1669),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1638),
.B(n_665),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1661),
.A2(n_368),
.B(n_367),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1610),
.Y(n_1758)
);

INVx4_ASAP7_75t_SL g1759 ( 
.A(n_1592),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1627),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1629),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1632),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1631),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1672),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1642),
.B(n_139),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1605),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1614),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_L g1768 ( 
.A1(n_1618),
.A2(n_140),
.B(n_141),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1626),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1600),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1656),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1609),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1624),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_SL g1774 ( 
.A(n_1612),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1616),
.B(n_140),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1611),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1577),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_SL g1778 ( 
.A1(n_1676),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1585),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1622),
.A2(n_142),
.B(n_144),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1578),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1635),
.B(n_144),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1578),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1578),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1589),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1578),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1578),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1585),
.Y(n_1788)
);

AND2x4_ASAP7_75t_SL g1789 ( 
.A(n_1596),
.B(n_369),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1585),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1601),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1589),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1578),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1635),
.B(n_145),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1585),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1585),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1585),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1589),
.Y(n_1798)
);

AO21x2_ASAP7_75t_L g1799 ( 
.A1(n_1652),
.A2(n_145),
.B(n_146),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1630),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1579),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1578),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1635),
.B(n_147),
.Y(n_1803)
);

AOI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1652),
.A2(n_147),
.B(n_148),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1579),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1585),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1578),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1578),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1647),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1700),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1677),
.Y(n_1811)
);

AO21x2_ASAP7_75t_L g1812 ( 
.A1(n_1696),
.A2(n_149),
.B(n_150),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1678),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1687),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1679),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1781),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1692),
.B(n_1785),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1688),
.Y(n_1818)
);

AO21x1_ASAP7_75t_L g1819 ( 
.A1(n_1738),
.A2(n_151),
.B(n_152),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1779),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1783),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1784),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1790),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1792),
.Y(n_1825)
);

OA21x2_ASAP7_75t_L g1826 ( 
.A1(n_1682),
.A2(n_152),
.B(n_153),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1795),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1680),
.B(n_153),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1798),
.B(n_154),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1801),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1744),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1796),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1801),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1686),
.B(n_370),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1681),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1786),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1797),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1806),
.Y(n_1838)
);

AO21x2_ASAP7_75t_L g1839 ( 
.A1(n_1696),
.A2(n_371),
.B(n_372),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1724),
.B(n_373),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1787),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1793),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1802),
.Y(n_1843)
);

AO21x2_ASAP7_75t_L g1844 ( 
.A1(n_1804),
.A2(n_375),
.B(n_377),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1804),
.A2(n_378),
.B(n_379),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1807),
.Y(n_1846)
);

BUFx2_ASAP7_75t_L g1847 ( 
.A(n_1725),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1742),
.B(n_380),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1805),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1720),
.B(n_382),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1805),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1683),
.B(n_384),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1808),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1691),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1689),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1707),
.A2(n_385),
.B(n_386),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1713),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1694),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1708),
.A2(n_387),
.B(n_388),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1706),
.Y(n_1860)
);

AO21x2_ASAP7_75t_L g1861 ( 
.A1(n_1710),
.A2(n_389),
.B(n_390),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1701),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1698),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1699),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1697),
.B(n_391),
.Y(n_1865)
);

AO21x2_ASAP7_75t_L g1866 ( 
.A1(n_1711),
.A2(n_392),
.B(n_394),
.Y(n_1866)
);

OA21x2_ASAP7_75t_L g1867 ( 
.A1(n_1693),
.A2(n_664),
.B(n_395),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1703),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1709),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1716),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1763),
.A2(n_399),
.B1(n_396),
.B2(n_397),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1718),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1717),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1721),
.B(n_401),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1712),
.B(n_402),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1693),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1809),
.A2(n_1766),
.B1(n_1769),
.B2(n_1763),
.C(n_1768),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1715),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1780),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1722),
.B(n_403),
.Y(n_1880)
);

AO21x2_ASAP7_75t_L g1881 ( 
.A1(n_1726),
.A2(n_404),
.B(n_405),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1728),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1777),
.B(n_406),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1748),
.A2(n_1685),
.B(n_1702),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1780),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1799),
.Y(n_1886)
);

BUFx12f_ASAP7_75t_L g1887 ( 
.A(n_1705),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1732),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1717),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1729),
.A2(n_407),
.B(n_408),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1736),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1729),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1690),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1747),
.B(n_409),
.Y(n_1894)
);

OA21x2_ASAP7_75t_L g1895 ( 
.A1(n_1714),
.A2(n_660),
.B(n_410),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1810),
.B(n_1723),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1889),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1825),
.B(n_1817),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1892),
.B(n_1782),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1892),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1873),
.B(n_1754),
.Y(n_1901)
);

INVxp67_ASAP7_75t_SL g1902 ( 
.A(n_1849),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1889),
.B(n_1737),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1811),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1876),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1891),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1830),
.B(n_1744),
.Y(n_1907)
);

OAI211xp5_ASAP7_75t_L g1908 ( 
.A1(n_1877),
.A2(n_1778),
.B(n_1727),
.C(n_1746),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1811),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1847),
.B(n_1791),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1815),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1815),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1816),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1870),
.B(n_1794),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1816),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1882),
.B(n_1760),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1821),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1841),
.B(n_1803),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1830),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1819),
.A2(n_1770),
.B1(n_1767),
.B2(n_1756),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1857),
.B(n_1731),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1821),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1872),
.B(n_1869),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1888),
.B(n_1833),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1888),
.B(n_1762),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1833),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1829),
.Y(n_1927)
);

NOR2x1_ASAP7_75t_L g1928 ( 
.A(n_1867),
.B(n_1741),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1822),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1851),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1851),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1884),
.B(n_1704),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1858),
.B(n_1743),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1893),
.B(n_1800),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1813),
.B(n_1735),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1814),
.B(n_1758),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1822),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1836),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1857),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1836),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1842),
.Y(n_1941)
);

BUFx2_ASAP7_75t_SL g1942 ( 
.A(n_1831),
.Y(n_1942)
);

NOR2x1_ASAP7_75t_SL g1943 ( 
.A(n_1879),
.B(n_1885),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1818),
.B(n_1730),
.Y(n_1944)
);

INVxp67_ASAP7_75t_SL g1945 ( 
.A(n_1842),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1820),
.B(n_1750),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1879),
.A2(n_1684),
.B(n_1734),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1843),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1843),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1823),
.B(n_1730),
.Y(n_1950)
);

INVx3_ASAP7_75t_SL g1951 ( 
.A(n_1857),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1835),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1860),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1846),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1890),
.A2(n_1765),
.B(n_1761),
.C(n_1695),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1887),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1824),
.B(n_1745),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1831),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1886),
.B(n_1755),
.C(n_1749),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1846),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1827),
.B(n_1739),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1853),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1853),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1868),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1895),
.A2(n_1774),
.B1(n_1756),
.B2(n_1772),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1860),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1855),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1863),
.B(n_1864),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1832),
.B(n_1753),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1895),
.A2(n_1773),
.B1(n_1764),
.B2(n_1771),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1837),
.B(n_1759),
.Y(n_1971)
);

INVx4_ASAP7_75t_L g1972 ( 
.A(n_1867),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1855),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1838),
.B(n_1759),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1932),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1953),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1951),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1966),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1904),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1932),
.B(n_1862),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1943),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1947),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_SL g1983 ( 
.A1(n_1965),
.A2(n_1828),
.B1(n_1812),
.B2(n_1775),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1910),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1940),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1898),
.B(n_1854),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1901),
.B(n_1886),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1909),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1948),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1924),
.B(n_1885),
.Y(n_1990)
);

OR2x2_ASAP7_75t_SL g1991 ( 
.A(n_1935),
.B(n_1826),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1896),
.B(n_1878),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1945),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1911),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1912),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1927),
.B(n_1862),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1913),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1907),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1915),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1903),
.B(n_1850),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1917),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1922),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1923),
.B(n_1826),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1949),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1900),
.Y(n_2005)
);

NOR2x1_ASAP7_75t_L g2006 ( 
.A(n_1928),
.B(n_1839),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1906),
.B(n_1894),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1956),
.B(n_1719),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1929),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1907),
.B(n_1834),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1952),
.B(n_1852),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1958),
.B(n_1875),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1937),
.A2(n_1845),
.B(n_1844),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1902),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1925),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1944),
.B(n_1883),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1938),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1900),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1936),
.B(n_1880),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1941),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1960),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1954),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1962),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1979),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1975),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2014),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1988),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1998),
.B(n_2010),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1975),
.Y(n_2029)
);

BUFx3_ASAP7_75t_L g2030 ( 
.A(n_2008),
.Y(n_2030)
);

OR2x2_ASAP7_75t_SL g2031 ( 
.A(n_1981),
.B(n_1899),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1994),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1980),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1998),
.B(n_1971),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2010),
.B(n_1974),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_SL g2036 ( 
.A(n_1977),
.B(n_1972),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1980),
.B(n_1972),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1987),
.B(n_1939),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_2005),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1995),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1990),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2015),
.B(n_1916),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1983),
.B(n_1970),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1997),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_2018),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1984),
.B(n_1969),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2012),
.B(n_1950),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1996),
.B(n_1961),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1999),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2003),
.B(n_1957),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2001),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1985),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2019),
.B(n_1957),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2016),
.B(n_1942),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2007),
.B(n_1942),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1976),
.B(n_1934),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1993),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1976),
.B(n_1934),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1986),
.B(n_1933),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1982),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2002),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2009),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1992),
.B(n_1905),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1989),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1978),
.B(n_1921),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2004),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2024),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2034),
.B(n_2000),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2035),
.B(n_1978),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2024),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2043),
.B(n_1993),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2026),
.B(n_1991),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2027),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2027),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2059),
.B(n_1918),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2039),
.Y(n_2076)
);

AOI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2036),
.A2(n_1908),
.B(n_1955),
.C(n_1959),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_2030),
.B(n_2017),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2028),
.B(n_2020),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_2065),
.B(n_2006),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2045),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_2065),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2048),
.B(n_1920),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2050),
.B(n_1946),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2040),
.Y(n_2085)
);

NAND2x1p5_ASAP7_75t_L g2086 ( 
.A(n_2037),
.B(n_1905),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2031),
.B(n_2052),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2055),
.B(n_2022),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2040),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2061),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2056),
.A2(n_2013),
.B1(n_1865),
.B2(n_2011),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2042),
.B(n_2023),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_SL g2093 ( 
.A(n_2082),
.B(n_2076),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2078),
.B(n_2053),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_SL g2095 ( 
.A(n_2081),
.B(n_2060),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2077),
.B(n_2056),
.Y(n_2096)
);

NOR2x1_ASAP7_75t_L g2097 ( 
.A(n_2080),
.B(n_2060),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2083),
.B(n_2058),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2071),
.B(n_2046),
.Y(n_2099)
);

NAND2xp33_ASAP7_75t_SL g2100 ( 
.A(n_2087),
.B(n_2054),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2068),
.B(n_2033),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2072),
.B(n_2057),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2092),
.B(n_2058),
.Y(n_2103)
);

AO221x2_ASAP7_75t_L g2104 ( 
.A1(n_2067),
.A2(n_2029),
.B1(n_2025),
.B2(n_2062),
.C(n_2061),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_2080),
.Y(n_2105)
);

NOR2x1_ASAP7_75t_L g2106 ( 
.A(n_2070),
.B(n_2037),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_2091),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_2073),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_SL g2109 ( 
.A1(n_2086),
.A2(n_1752),
.B1(n_2044),
.B2(n_2032),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2075),
.A2(n_2041),
.B1(n_2051),
.B2(n_2049),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2074),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2106),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2105),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_2104),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2111),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2102),
.B(n_2069),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2099),
.B(n_2079),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2104),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2101),
.B(n_2088),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2097),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2103),
.B(n_2084),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_2107),
.A2(n_2085),
.B1(n_2090),
.B2(n_2089),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2108),
.B(n_2064),
.Y(n_2123)
);

NAND3xp33_ASAP7_75t_L g2124 ( 
.A(n_2095),
.B(n_2062),
.C(n_2066),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2110),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_2109),
.B(n_2047),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2098),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2096),
.B(n_2063),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2113),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2116),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2119),
.B(n_2094),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2125),
.B(n_2093),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2115),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2118),
.Y(n_2134)
);

O2A1O1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_2118),
.A2(n_2100),
.B(n_2013),
.C(n_1752),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2112),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_2128),
.B(n_2038),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2120),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2122),
.B(n_1871),
.C(n_1848),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_2124),
.B(n_1914),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2114),
.Y(n_2141)
);

INVx1_ASAP7_75t_SL g2142 ( 
.A(n_2121),
.Y(n_2142)
);

NAND3xp33_ASAP7_75t_L g2143 ( 
.A(n_2127),
.B(n_1776),
.C(n_1840),
.Y(n_2143)
);

NOR2x1_ASAP7_75t_L g2144 ( 
.A(n_2129),
.B(n_2123),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2130),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2142),
.B(n_2126),
.Y(n_2146)
);

O2A1O1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_2132),
.A2(n_2117),
.B(n_1856),
.C(n_1866),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2134),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2141),
.Y(n_2149)
);

OAI31xp33_ASAP7_75t_L g2150 ( 
.A1(n_2135),
.A2(n_1789),
.A3(n_1926),
.B(n_1840),
.Y(n_2150)
);

INVxp67_ASAP7_75t_L g2151 ( 
.A(n_2131),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2136),
.B(n_2021),
.Y(n_2152)
);

AOI322xp5_ASAP7_75t_L g2153 ( 
.A1(n_2140),
.A2(n_1897),
.A3(n_1967),
.B1(n_1963),
.B2(n_1930),
.C1(n_1919),
.C2(n_1931),
.Y(n_2153)
);

AOI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_2138),
.A2(n_1968),
.B1(n_1964),
.B2(n_1973),
.C(n_1861),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2133),
.Y(n_2155)
);

AOI211xp5_ASAP7_75t_L g2156 ( 
.A1(n_2139),
.A2(n_1751),
.B(n_1874),
.C(n_1757),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2143),
.Y(n_2157)
);

AOI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_2147),
.A2(n_2137),
.B(n_1740),
.Y(n_2158)
);

NAND3xp33_ASAP7_75t_L g2159 ( 
.A(n_2146),
.B(n_1874),
.C(n_1733),
.Y(n_2159)
);

OAI31xp33_ASAP7_75t_L g2160 ( 
.A1(n_2150),
.A2(n_1733),
.A3(n_1881),
.B(n_1859),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2149),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_2151),
.B(n_2157),
.Y(n_2162)
);

OAI211xp5_ASAP7_75t_L g2163 ( 
.A1(n_2144),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2145),
.Y(n_2164)
);

OAI322xp33_ASAP7_75t_L g2165 ( 
.A1(n_2148),
.A2(n_414),
.A3(n_415),
.B1(n_416),
.B2(n_417),
.C1(n_419),
.C2(n_420),
.Y(n_2165)
);

OAI211xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2155),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2152),
.B(n_424),
.Y(n_2167)
);

OAI221xp5_ASAP7_75t_L g2168 ( 
.A1(n_2156),
.A2(n_428),
.B1(n_425),
.B2(n_426),
.C(n_429),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2154),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2162),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2161),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2164),
.Y(n_2172)
);

NAND2xp33_ASAP7_75t_L g2173 ( 
.A(n_2167),
.B(n_2169),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2158),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2159),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2163),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2165),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2168),
.Y(n_2178)
);

INVxp67_ASAP7_75t_L g2179 ( 
.A(n_2166),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2160),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2162),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_2162),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2162),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_2167),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2173),
.A2(n_2153),
.B(n_433),
.Y(n_2185)
);

AO22x2_ASAP7_75t_L g2186 ( 
.A1(n_2174),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2170),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_2182),
.A2(n_437),
.B(n_438),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2181),
.Y(n_2189)
);

NOR2xp67_ASAP7_75t_L g2190 ( 
.A(n_2183),
.B(n_2171),
.Y(n_2190)
);

NOR2xp67_ASAP7_75t_L g2191 ( 
.A(n_2172),
.B(n_439),
.Y(n_2191)
);

NAND3xp33_ASAP7_75t_L g2192 ( 
.A(n_2180),
.B(n_2175),
.C(n_2176),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2184),
.Y(n_2193)
);

AOI211xp5_ASAP7_75t_L g2194 ( 
.A1(n_2177),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_2194)
);

NOR2xp67_ASAP7_75t_L g2195 ( 
.A(n_2179),
.B(n_444),
.Y(n_2195)
);

OAI211xp5_ASAP7_75t_L g2196 ( 
.A1(n_2192),
.A2(n_2178),
.B(n_448),
.C(n_446),
.Y(n_2196)
);

AOI221x1_ASAP7_75t_L g2197 ( 
.A1(n_2186),
.A2(n_447),
.B1(n_450),
.B2(n_451),
.C(n_452),
.Y(n_2197)
);

O2A1O1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_2193),
.A2(n_457),
.B(n_454),
.C(n_456),
.Y(n_2198)
);

AOI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2190),
.A2(n_462),
.B(n_458),
.C(n_460),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_2187),
.B(n_463),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_2185),
.A2(n_464),
.B(n_465),
.Y(n_2201)
);

A2O1A1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2191),
.A2(n_2195),
.B(n_2189),
.C(n_2188),
.Y(n_2202)
);

AOI211xp5_ASAP7_75t_L g2203 ( 
.A1(n_2194),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_2203)
);

NAND3xp33_ASAP7_75t_SL g2204 ( 
.A(n_2194),
.B(n_472),
.C(n_473),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_2192),
.B(n_475),
.C(n_477),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2202),
.B(n_478),
.Y(n_2206)
);

NOR3xp33_ASAP7_75t_L g2207 ( 
.A(n_2196),
.B(n_480),
.C(n_481),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_2200),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2201),
.B(n_482),
.Y(n_2209)
);

NAND3xp33_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_2203),
.C(n_2205),
.Y(n_2210)
);

AOI221xp5_ASAP7_75t_L g2211 ( 
.A1(n_2204),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.C(n_487),
.Y(n_2211)
);

NAND3xp33_ASAP7_75t_L g2212 ( 
.A(n_2199),
.B(n_488),
.C(n_489),
.Y(n_2212)
);

NAND3xp33_ASAP7_75t_L g2213 ( 
.A(n_2198),
.B(n_490),
.C(n_491),
.Y(n_2213)
);

NAND3xp33_ASAP7_75t_L g2214 ( 
.A(n_2197),
.B(n_492),
.C(n_493),
.Y(n_2214)
);

NOR3xp33_ASAP7_75t_L g2215 ( 
.A(n_2196),
.B(n_494),
.C(n_495),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2204),
.A2(n_499),
.B1(n_496),
.B2(n_497),
.Y(n_2216)
);

OAI321xp33_ASAP7_75t_L g2217 ( 
.A1(n_2196),
.A2(n_500),
.A3(n_501),
.B1(n_502),
.B2(n_503),
.C(n_504),
.Y(n_2217)
);

NAND3xp33_ASAP7_75t_L g2218 ( 
.A(n_2197),
.B(n_507),
.C(n_508),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2206),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2208),
.B(n_510),
.Y(n_2220)
);

OAI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_2210),
.A2(n_511),
.B(n_512),
.Y(n_2221)
);

NOR4xp25_ASAP7_75t_L g2222 ( 
.A(n_2214),
.B(n_516),
.C(n_513),
.D(n_515),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2218),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_2209),
.B(n_517),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2216),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2212),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2207),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2215),
.A2(n_521),
.B1(n_518),
.B2(n_519),
.Y(n_2228)
);

NOR4xp75_ASAP7_75t_L g2229 ( 
.A(n_2217),
.B(n_523),
.C(n_527),
.D(n_528),
.Y(n_2229)
);

NOR2x1_ASAP7_75t_L g2230 ( 
.A(n_2213),
.B(n_529),
.Y(n_2230)
);

NAND4xp75_ASAP7_75t_L g2231 ( 
.A(n_2211),
.B(n_530),
.C(n_532),
.D(n_533),
.Y(n_2231)
);

NOR2x1_ASAP7_75t_L g2232 ( 
.A(n_2214),
.B(n_534),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_2219),
.B(n_535),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2232),
.B(n_536),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2224),
.B(n_537),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2231),
.Y(n_2236)
);

NAND3xp33_ASAP7_75t_L g2237 ( 
.A(n_2221),
.B(n_538),
.C(n_539),
.Y(n_2237)
);

NOR2x1_ASAP7_75t_L g2238 ( 
.A(n_2220),
.B(n_659),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2227),
.A2(n_540),
.B1(n_541),
.B2(n_543),
.Y(n_2239)
);

INVx4_ASAP7_75t_L g2240 ( 
.A(n_2223),
.Y(n_2240)
);

NAND3x1_ASAP7_75t_L g2241 ( 
.A(n_2230),
.B(n_544),
.C(n_546),
.Y(n_2241)
);

NAND4xp75_ASAP7_75t_SL g2242 ( 
.A(n_2229),
.B(n_547),
.C(n_551),
.D(n_552),
.Y(n_2242)
);

XNOR2x1_ASAP7_75t_L g2243 ( 
.A(n_2226),
.B(n_553),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_2225),
.B(n_554),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2228),
.Y(n_2245)
);

AND3x2_ASAP7_75t_L g2246 ( 
.A(n_2222),
.B(n_555),
.C(n_556),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2220),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2232),
.B(n_557),
.Y(n_2248)
);

XNOR2xp5_ASAP7_75t_L g2249 ( 
.A(n_2229),
.B(n_558),
.Y(n_2249)
);

AOI21xp5_ASAP7_75t_SL g2250 ( 
.A1(n_2221),
.A2(n_560),
.B(n_561),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_R g2251 ( 
.A(n_2249),
.B(n_562),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_2240),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2236),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2242),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2246),
.B(n_567),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2247),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2233),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2250),
.A2(n_2235),
.B(n_2243),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2238),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2234),
.B(n_568),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2244),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2248),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2241),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2252),
.A2(n_2256),
.B1(n_2245),
.B2(n_2261),
.Y(n_2264)
);

NAND4xp25_ASAP7_75t_L g2265 ( 
.A(n_2258),
.B(n_2237),
.C(n_2239),
.D(n_571),
.Y(n_2265)
);

BUFx3_ASAP7_75t_L g2266 ( 
.A(n_2252),
.Y(n_2266)
);

AO22x2_ASAP7_75t_L g2267 ( 
.A1(n_2259),
.A2(n_569),
.B1(n_570),
.B2(n_572),
.Y(n_2267)
);

AOI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2254),
.A2(n_573),
.B1(n_575),
.B2(n_576),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2255),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.Y(n_2269)
);

OAI22x1_ASAP7_75t_L g2270 ( 
.A1(n_2263),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_2270)
);

OAI22x1_ASAP7_75t_L g2271 ( 
.A1(n_2257),
.A2(n_583),
.B1(n_584),
.B2(n_585),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2260),
.Y(n_2272)
);

OAI22x1_ASAP7_75t_L g2273 ( 
.A1(n_2262),
.A2(n_2253),
.B1(n_2251),
.B2(n_589),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2266),
.Y(n_2274)
);

OAI22x1_ASAP7_75t_L g2275 ( 
.A1(n_2264),
.A2(n_586),
.B1(n_587),
.B2(n_590),
.Y(n_2275)
);

XNOR2xp5_ASAP7_75t_L g2276 ( 
.A(n_2273),
.B(n_591),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2272),
.A2(n_592),
.B1(n_594),
.B2(n_595),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2265),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2274),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_SL g2280 ( 
.A1(n_2276),
.A2(n_2269),
.B(n_2268),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2278),
.A2(n_2267),
.B1(n_2270),
.B2(n_2271),
.Y(n_2281)
);

CKINVDCx20_ASAP7_75t_R g2282 ( 
.A(n_2279),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2281),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2283),
.A2(n_2280),
.B(n_2275),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2282),
.Y(n_2285)
);

AOI211xp5_ASAP7_75t_L g2286 ( 
.A1(n_2285),
.A2(n_2277),
.B(n_2267),
.C(n_601),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_SL g2287 ( 
.A1(n_2284),
.A2(n_599),
.B1(n_600),
.B2(n_602),
.Y(n_2287)
);

AO21x2_ASAP7_75t_L g2288 ( 
.A1(n_2287),
.A2(n_603),
.B(n_605),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2286),
.A2(n_607),
.B(n_608),
.Y(n_2289)
);

AOI21x1_ASAP7_75t_L g2290 ( 
.A1(n_2289),
.A2(n_658),
.B(n_610),
.Y(n_2290)
);

AOI221xp5_ASAP7_75t_L g2291 ( 
.A1(n_2288),
.A2(n_609),
.B1(n_611),
.B2(n_612),
.C(n_613),
.Y(n_2291)
);

AOI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_2291),
.A2(n_614),
.B1(n_615),
.B2(n_617),
.C(n_618),
.Y(n_2292)
);

OA22x2_ASAP7_75t_L g2293 ( 
.A1(n_2292),
.A2(n_2290),
.B1(n_619),
.B2(n_620),
.Y(n_2293)
);


endmodule