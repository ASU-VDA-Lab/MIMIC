module fake_aes_3159_n_15 (n_3, n_1, n_2, n_0, n_15);
input n_3;
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_7), .B(n_0), .Y(n_10) );
AO21x2_ASAP7_75t_L g11 ( .A1(n_6), .A2(n_1), .B(n_3), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
NOR3xp33_ASAP7_75t_L g13 ( .A(n_12), .B(n_10), .C(n_8), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
AOI21xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_11), .B(n_1), .Y(n_15) );
endmodule