module fake_netlist_1_4315_n_489 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_489);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_489;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_6), .Y(n_75) );
NOR2xp33_ASAP7_75t_L g76 ( .A(n_5), .B(n_46), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_71), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_26), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_3), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_17), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_37), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_62), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_9), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_67), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_64), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_36), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_0), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_5), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_11), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_56), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_70), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_32), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_51), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_30), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_3), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_88), .B(n_0), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_84), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_80), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_106), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_75), .B(n_1), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_82), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_78), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_84), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_75), .B(n_1), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_86), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_2), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_108), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
NOR2xp67_ASAP7_75t_L g127 ( .A(n_101), .B(n_4), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_79), .B(n_4), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_90), .B(n_6), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_83), .B(n_7), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_119), .B(n_90), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_119), .A2(n_97), .B1(n_94), .B2(n_95), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_126), .B(n_92), .Y(n_137) );
OAI22xp33_ASAP7_75t_SL g138 ( .A1(n_117), .A2(n_111), .B1(n_94), .B2(n_95), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_113), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_115), .B(n_100), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_125), .B(n_115), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_125), .B(n_111), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_125), .B(n_97), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_126), .B(n_105), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_128), .B(n_92), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_113), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_128), .B(n_109), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_129), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_132), .A2(n_105), .B1(n_93), .B2(n_96), .Y(n_155) );
XOR2xp5_ASAP7_75t_L g156 ( .A(n_155), .B(n_114), .Y(n_156) );
NOR3xp33_ASAP7_75t_SL g157 ( .A(n_140), .B(n_116), .C(n_124), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
NOR2xp33_ASAP7_75t_R g160 ( .A(n_146), .B(n_123), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_143), .B(n_132), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_154), .B(n_118), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_145), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_146), .B(n_123), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_145), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_141), .B(n_118), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_141), .Y(n_169) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_143), .B(n_132), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
CKINVDCx11_ASAP7_75t_R g174 ( .A(n_143), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_154), .B(n_112), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_143), .Y(n_177) );
NOR2xp33_ASAP7_75t_R g178 ( .A(n_151), .B(n_129), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVxp67_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_144), .B(n_112), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
AOI21xp33_ASAP7_75t_L g186 ( .A1(n_163), .A2(n_144), .B(n_155), .Y(n_186) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_181), .Y(n_187) );
BUFx4_ASAP7_75t_SL g188 ( .A(n_161), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_181), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_183), .B(n_144), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_181), .B(n_147), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_170), .B(n_147), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_168), .B(n_138), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_170), .B(n_147), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_183), .A2(n_150), .B(n_137), .Y(n_199) );
CKINVDCx8_ASAP7_75t_R g200 ( .A(n_161), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_177), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
INVxp33_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_162), .B(n_147), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_168), .A2(n_138), .B(n_117), .C(n_121), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_162), .Y(n_211) );
INVx8_ASAP7_75t_L g212 ( .A(n_162), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_180), .Y(n_213) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_131), .A3(n_134), .B(n_137), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_184), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_198), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_200), .B(n_180), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_198), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_192), .B(n_169), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_215), .Y(n_220) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_207), .B(n_174), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_192), .B(n_172), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_192), .B(n_172), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_194), .A2(n_175), .B1(n_147), .B2(n_135), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_215), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_191), .B(n_185), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_192), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_186), .A2(n_135), .B1(n_121), .B2(n_131), .C(n_134), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_206), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_200), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_205), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_205), .A2(n_156), .B1(n_172), .B2(n_179), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_214), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_189), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_189), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_193), .A2(n_156), .B1(n_150), .B2(n_127), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_214), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_226), .B(n_193), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g243 ( .A1(n_239), .A2(n_203), .B1(n_197), .B2(n_157), .C(n_209), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_218), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g245 ( .A1(n_239), .A2(n_203), .B1(n_197), .B2(n_207), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_213), .B1(n_148), .B2(n_211), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_236), .A2(n_199), .B(n_152), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_226), .B(n_205), .Y(n_248) );
NOR2xp33_ASAP7_75t_R g249 ( .A(n_221), .B(n_190), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_236), .B(n_214), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_216), .Y(n_251) );
OAI221xp5_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_211), .B1(n_187), .B2(n_208), .C(n_210), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_213), .B1(n_148), .B2(n_212), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_219), .A2(n_205), .B1(n_212), .B2(n_190), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_230), .B(n_130), .C(n_120), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_205), .B1(n_212), .B2(n_196), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_218), .Y(n_258) );
OAI33xp33_ASAP7_75t_L g259 ( .A1(n_240), .A2(n_81), .A3(n_107), .B1(n_104), .B2(n_85), .B3(n_87), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_233), .B(n_205), .Y(n_261) );
OAI31xp33_ASAP7_75t_L g262 ( .A1(n_253), .A2(n_219), .A3(n_227), .B(n_229), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_258), .A2(n_240), .B(n_238), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_244), .Y(n_264) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_256), .A2(n_238), .B(n_237), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_256), .B(n_230), .C(n_130), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_250), .B(n_220), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_251), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_253), .A2(n_221), .B1(n_219), .B2(n_233), .Y(n_269) );
OAI31xp33_ASAP7_75t_SL g270 ( .A1(n_246), .A2(n_217), .A3(n_220), .B(n_223), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_250), .B(n_225), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_244), .B(n_225), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_251), .B(n_214), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_244), .Y(n_274) );
AOI211xp5_ASAP7_75t_L g275 ( .A1(n_243), .A2(n_232), .B(n_227), .C(n_127), .Y(n_275) );
OAI21xp5_ASAP7_75t_SL g276 ( .A1(n_246), .A2(n_222), .B(n_223), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_254), .B(n_214), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_260), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_260), .B(n_225), .Y(n_279) );
NAND2x1_ASAP7_75t_L g280 ( .A(n_260), .B(n_228), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_241), .B(n_225), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_267), .B(n_247), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_267), .B(n_247), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_276), .A2(n_245), .B1(n_241), .B2(n_221), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_278), .Y(n_289) );
OAI31xp33_ASAP7_75t_L g290 ( .A1(n_262), .A2(n_248), .A3(n_252), .B(n_261), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_271), .B(n_242), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_273), .B(n_242), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_271), .B(n_248), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_273), .B(n_261), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_262), .A2(n_249), .B1(n_259), .B2(n_261), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
AOI322xp5_ASAP7_75t_L g297 ( .A1(n_269), .A2(n_255), .A3(n_257), .B1(n_261), .B2(n_87), .C1(n_99), .C2(n_81), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_277), .B(n_234), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_278), .B(n_85), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_268), .B(n_98), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_234), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_282), .B(n_234), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_282), .B(n_237), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_281), .B(n_237), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_270), .B(n_238), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_272), .B(n_98), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_272), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_276), .B(n_231), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_291), .B(n_270), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_281), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_292), .B(n_263), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_296), .B(n_275), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_291), .B(n_272), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_303), .B(n_272), .Y(n_318) );
AOI31xp67_ASAP7_75t_SL g319 ( .A1(n_307), .A2(n_275), .A3(n_102), .B(n_103), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_301), .B(n_279), .Y(n_320) );
NAND2xp33_ASAP7_75t_SL g321 ( .A(n_303), .B(n_280), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_299), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_301), .B(n_279), .Y(n_324) );
BUFx2_ASAP7_75t_SL g325 ( .A(n_299), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_293), .B(n_263), .Y(n_326) );
NOR2x1p5_ASAP7_75t_L g327 ( .A(n_307), .B(n_266), .Y(n_327) );
NAND2x1_ASAP7_75t_L g328 ( .A(n_285), .B(n_279), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_286), .B(n_265), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_297), .A2(n_266), .B(n_77), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_308), .B(n_279), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_310), .B(n_99), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_287), .B(n_233), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_293), .B(n_302), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_302), .B(n_280), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_286), .B(n_265), .Y(n_341) );
OAI211xp5_ASAP7_75t_L g342 ( .A1(n_287), .A2(n_233), .B(n_76), .C(n_110), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_308), .B(n_102), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_300), .B(n_103), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_283), .B(n_265), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_298), .B(n_265), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_298), .B(n_306), .Y(n_347) );
NAND2x1p5_ASAP7_75t_SL g348 ( .A(n_300), .B(n_109), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_304), .B(n_104), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_339), .B(n_284), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_290), .B(n_295), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_309), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_323), .B(n_304), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_336), .A2(n_295), .B1(n_309), .B2(n_304), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_336), .A2(n_329), .B(n_338), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_342), .A2(n_349), .B(n_315), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_334), .Y(n_359) );
NOR2x1_ASAP7_75t_L g360 ( .A(n_342), .B(n_284), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_318), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_337), .A2(n_289), .B1(n_288), .B2(n_284), .Y(n_363) );
NAND4xp25_ASAP7_75t_SL g364 ( .A(n_311), .B(n_297), .C(n_290), .D(n_110), .Y(n_364) );
AOI322xp5_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_107), .A3(n_288), .B1(n_289), .B2(n_120), .C1(n_113), .C2(n_12), .Y(n_365) );
OAI322xp33_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_306), .A3(n_120), .B1(n_113), .B2(n_289), .C1(n_288), .C2(n_12), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_319), .A2(n_265), .B1(n_223), .B2(n_222), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_347), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_333), .B(n_328), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_319), .A2(n_223), .B1(n_222), .B2(n_212), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_332), .A2(n_120), .B1(n_113), .B2(n_222), .C1(n_10), .C2(n_11), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_333), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_312), .B(n_7), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_325), .A2(n_228), .B1(n_120), .B2(n_178), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_326), .B(n_8), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_343), .B(n_8), .Y(n_378) );
XNOR2xp5_ASAP7_75t_L g379 ( .A(n_348), .B(n_9), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_314), .B(n_13), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_320), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_333), .A2(n_228), .B1(n_120), .B2(n_195), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
INVxp33_ASAP7_75t_L g385 ( .A(n_335), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_344), .A2(n_120), .B1(n_133), .B2(n_139), .C(n_149), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_331), .B(n_13), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_321), .B(n_14), .C(n_15), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_333), .B(n_14), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_327), .A2(n_228), .B1(n_202), .B2(n_201), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_341), .B(n_346), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_341), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_348), .A2(n_15), .B(n_16), .C(n_18), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_381), .B(n_16), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_395), .B(n_18), .C(n_133), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_351), .B(n_133), .C(n_139), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_389), .B(n_19), .C(n_23), .Y(n_401) );
NOR2x1p5_ASAP7_75t_L g402 ( .A(n_362), .B(n_228), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_387), .B(n_24), .Y(n_405) );
AOI322xp5_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_139), .A3(n_149), .B1(n_152), .B2(n_153), .C1(n_164), .C2(n_179), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_360), .A2(n_228), .B(n_204), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_393), .B(n_25), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_392), .B(n_27), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_383), .B(n_153), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_355), .B(n_153), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_388), .B(n_152), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_384), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_353), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_352), .B(n_28), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_359), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_370), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_354), .B(n_171), .C(n_164), .D(n_173), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_358), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_390), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_357), .Y(n_423) );
OAI21xp33_ASAP7_75t_SL g424 ( .A1(n_373), .A2(n_31), .B(n_33), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_385), .B(n_35), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_363), .B(n_38), .Y(n_426) );
XNOR2x2_ASAP7_75t_L g427 ( .A(n_379), .B(n_40), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g428 ( .A1(n_370), .A2(n_195), .B(n_189), .Y(n_428) );
NAND2x1_ASAP7_75t_L g429 ( .A(n_390), .B(n_204), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_391), .B(n_204), .Y(n_430) );
NOR4xp25_ASAP7_75t_SL g431 ( .A(n_356), .B(n_42), .C(n_43), .D(n_44), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_356), .B(n_45), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_419), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_423), .B(n_378), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_421), .Y(n_437) );
NAND4xp75_ASAP7_75t_L g438 ( .A(n_424), .B(n_386), .C(n_364), .D(n_366), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_433), .A2(n_371), .B1(n_367), .B2(n_391), .C(n_382), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_427), .A2(n_372), .B1(n_367), .B2(n_371), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_422), .A2(n_372), .B(n_365), .C(n_376), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_432), .A2(n_404), .B1(n_396), .B2(n_413), .C1(n_403), .C2(n_415), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g443 ( .A(n_427), .B(n_47), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_414), .B(n_418), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g445 ( .A1(n_402), .A2(n_173), .A3(n_172), .B(n_185), .Y(n_445) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_397), .B(n_48), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_434), .B(n_50), .Y(n_447) );
AOI221x1_ASAP7_75t_L g448 ( .A1(n_398), .A2(n_204), .B1(n_195), .B2(n_185), .C(n_165), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_401), .B(n_430), .C(n_428), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
OA22x2_ASAP7_75t_L g452 ( .A1(n_408), .A2(n_52), .B1(n_54), .B2(n_55), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_401), .A2(n_165), .B(n_195), .C(n_167), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_430), .A2(n_165), .A3(n_60), .B(n_61), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_420), .A2(n_182), .B1(n_159), .B2(n_158), .C(n_167), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_429), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_426), .B(n_159), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_442), .B(n_400), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g459 ( .A1(n_443), .A2(n_408), .B(n_426), .Y(n_459) );
NOR3xp33_ASAP7_75t_SL g460 ( .A(n_441), .B(n_425), .C(n_412), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
OAI21xp33_ASAP7_75t_SL g462 ( .A1(n_442), .A2(n_416), .B(n_405), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_449), .A2(n_408), .B(n_426), .Y(n_463) );
HB1xp67_ASAP7_75t_SL g464 ( .A(n_435), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_453), .A2(n_411), .B(n_431), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_440), .A2(n_409), .B(n_406), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_456), .B(n_407), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_439), .A2(n_410), .B1(n_158), .B2(n_167), .Y(n_468) );
NAND4xp75_ASAP7_75t_L g469 ( .A(n_439), .B(n_58), .C(n_65), .D(n_66), .Y(n_469) );
AOI322xp5_ASAP7_75t_L g470 ( .A1(n_436), .A2(n_68), .A3(n_72), .B1(n_73), .B2(n_74), .C1(n_182), .C2(n_167), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_438), .B(n_158), .C(n_182), .Y(n_471) );
OAI222xp33_ASAP7_75t_L g472 ( .A1(n_452), .A2(n_167), .B1(n_457), .B2(n_450), .C1(n_451), .C2(n_447), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_455), .B(n_167), .C(n_446), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_452), .A2(n_445), .B1(n_454), .B2(n_448), .Y(n_474) );
AOI221x1_ASAP7_75t_L g475 ( .A1(n_449), .A2(n_436), .B1(n_389), .B2(n_437), .C(n_423), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_440), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_476), .A2(n_462), .B1(n_460), .B2(n_459), .Y(n_477) );
AO22x2_ASAP7_75t_L g478 ( .A1(n_475), .A2(n_458), .B1(n_459), .B2(n_463), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_461), .B(n_471), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_468), .B(n_466), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_480), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_479), .Y(n_483) );
NAND5xp2_ASAP7_75t_L g484 ( .A(n_477), .B(n_473), .C(n_465), .D(n_470), .E(n_469), .Y(n_484) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_482), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_482), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_486), .Y(n_487) );
AOI322xp5_ASAP7_75t_L g488 ( .A1(n_487), .A2(n_485), .A3(n_483), .B1(n_481), .B2(n_478), .C1(n_484), .C2(n_467), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_488), .A2(n_472), .B(n_474), .Y(n_489) );
endmodule