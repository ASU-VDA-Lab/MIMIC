module fake_jpeg_3265_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_16),
.B(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_50),
.B1(n_51),
.B2(n_73),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_61),
.B1(n_64),
.B2(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_54),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_50),
.B1(n_55),
.B2(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_47),
.B1(n_49),
.B2(n_26),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_92),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_65),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_99),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_68),
.B(n_66),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_101),
.C(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_61),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_79),
.Y(n_115)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_116),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_114),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_22),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_64),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_113),
.B1(n_118),
.B2(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_47),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_15),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_90),
.B1(n_97),
.B2(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_21),
.B1(n_44),
.B2(n_42),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_147),
.B(n_9),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_144),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_20),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_29),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_0),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_13),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_157),
.B1(n_140),
.B2(n_146),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_4),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_165),
.B(n_166),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_161),
.B(n_167),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_34),
.B(n_41),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_18),
.C1(n_27),
.C2(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_157),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_149),
.CI(n_144),
.CON(n_170),
.SN(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_158),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_129),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_151),
.C(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_177),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_182),
.C(n_175),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_155),
.B(n_156),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_150),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_168),
.B(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_33),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_178),
.B1(n_188),
.B2(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_191),
.A3(n_176),
.B1(n_173),
.B2(n_129),
.C1(n_39),
.C2(n_35),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_37),
.C(n_38),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_193),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_189),
.Y(n_195)
);


endmodule