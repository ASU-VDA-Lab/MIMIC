module fake_jpeg_13514_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_70),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_37),
.B(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_51),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_42),
.C(n_46),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_6),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_52),
.B1(n_37),
.B2(n_46),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_67),
.B1(n_75),
.B2(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_20),
.Y(n_86)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_0),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_4),
.Y(n_106)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_24),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_23),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_106),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_12),
.Y(n_121)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_77),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_78),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_97),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_120),
.C(n_118),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_91),
.C(n_111),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_119),
.C(n_116),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_113),
.A3(n_108),
.B1(n_122),
.B2(n_125),
.C1(n_103),
.C2(n_126),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_108),
.B1(n_14),
.B2(n_19),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

AOI321xp33_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_13),
.A3(n_25),
.B1(n_28),
.B2(n_31),
.C(n_32),
.Y(n_136)
);

XNOR2x2_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_34),
.Y(n_137)
);


endmodule