module real_jpeg_11697_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_33),
.B1(n_52),
.B2(n_55),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_36),
.B(n_37),
.C(n_43),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_4),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_40),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_4),
.A2(n_40),
.B(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_25),
.C(n_85),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_39),
.B1(n_52),
.B2(n_55),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_4),
.A2(n_24),
.B1(n_27),
.B2(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_61),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_25),
.B1(n_31),
.B2(n_49),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_8),
.A2(n_30),
.B1(n_52),
.B2(n_55),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_52),
.B1(n_55),
.B2(n_67),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_10),
.A2(n_25),
.B1(n_31),
.B2(n_67),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_25),
.B1(n_31),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_11),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_52),
.B1(n_55),
.B2(n_79),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_52),
.B1(n_55),
.B2(n_69),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_13),
.A2(n_25),
.B1(n_31),
.B2(n_69),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_25),
.B1(n_31),
.B2(n_60),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_14),
.A2(n_52),
.B1(n_55),
.B2(n_60),
.Y(n_117)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_109),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.C(n_62),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_21),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_22),
.A2(n_34),
.B1(n_35),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_22),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_23),
.A2(n_76),
.B(n_97),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_23),
.A2(n_28),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_24),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_24),
.A2(n_27),
.B1(n_190),
.B2(n_198),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_24),
.A2(n_75),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_25),
.A2(n_31),
.B1(n_85),
.B2(n_86),
.Y(n_88)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_27),
.B(n_39),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_28),
.A2(n_29),
.B(n_77),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_31),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_40),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_39),
.B(n_88),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_56)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_SL g162 ( 
.A(n_41),
.B(n_53),
.C(n_55),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_62),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_57),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_59),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_50),
.A2(n_51),
.B1(n_121),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_50),
.A2(n_51),
.B1(n_145),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_55),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_52),
.A2(n_54),
.B(n_160),
.C(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_52),
.B(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_61),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_66),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_92),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_80),
.B2(n_91),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_88),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_83),
.A2(n_89),
.B1(n_155),
.B2(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_83),
.A2(n_89),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_83),
.A2(n_89),
.B1(n_177),
.B2(n_187),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_117),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_98),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_127),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_110),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_112),
.B(n_127),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.C(n_122),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_114),
.B1(n_119),
.B2(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B(n_118),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_226),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_221),
.B(n_222),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_165),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_150),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_135),
.B(n_150),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_139),
.B(n_146),
.C(n_148),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_157),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_163),
.B1(n_164),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_178),
.B(n_220),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_170),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.C(n_176),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_214),
.B(n_219),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_204),
.B(n_213),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_193),
.B(n_203),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_188),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_202),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_209),
.C(n_212),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_218),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);


endmodule