module fake_jpeg_9535_n_114 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_32),
.B(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_34),
.Y(n_37)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_6),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_34),
.B1(n_28),
.B2(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_20),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_61),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_11),
.Y(n_77)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_72),
.B1(n_73),
.B2(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_77),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_56),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_86),
.B(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_50),
.C(n_59),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_68),
.C(n_76),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_61),
.B1(n_46),
.B2(n_47),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_82),
.B(n_78),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_66),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_73),
.C(n_55),
.Y(n_94)
);

AOI31xp67_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_46),
.A3(n_86),
.B(n_81),
.Y(n_95)
);

AOI321xp33_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_14),
.A3(n_11),
.B1(n_63),
.B2(n_30),
.C(n_64),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_100),
.B(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_69),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_84),
.A3(n_65),
.B1(n_69),
.B2(n_53),
.C(n_23),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_67),
.B1(n_22),
.B2(n_12),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_93),
.B(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_57),
.B1(n_7),
.B2(n_8),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_101),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_108),
.C(n_7),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_109),
.C(n_10),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_112),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule