module fake_jpeg_24903_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_0),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_75),
.B1(n_84),
.B2(n_85),
.Y(n_98)
);

INVxp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_67),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_64),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_62),
.B1(n_72),
.B2(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_18),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_34),
.B1(n_33),
.B2(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_82),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_34),
.B1(n_33),
.B2(n_35),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_19),
.B1(n_24),
.B2(n_38),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_15),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_30),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_92),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_106),
.Y(n_125)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_31),
.B1(n_20),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_59),
.B1(n_79),
.B2(n_72),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_49),
.B(n_48),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_62),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_1),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_20),
.C(n_37),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_15),
.B(n_17),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_111),
.A3(n_17),
.B1(n_16),
.B2(n_3),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_115),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_15),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_1),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_57),
.B(n_13),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_137),
.B(n_147),
.Y(n_158)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_133),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_153),
.Y(n_166)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_53),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_135),
.Y(n_157)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_89),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_97),
.B(n_1),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_56),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_61),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_63),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_54),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_54),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_90),
.B(n_97),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_96),
.B(n_1),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_109),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_98),
.B1(n_113),
.B2(n_128),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_88),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_92),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_113),
.B1(n_145),
.B2(n_87),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_117),
.C(n_110),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_29),
.C(n_2),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_171),
.A2(n_143),
.B(n_7),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_88),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_178),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_87),
.B1(n_90),
.B2(n_95),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_90),
.B1(n_121),
.B2(n_88),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_140),
.B1(n_90),
.B2(n_124),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_186),
.B1(n_147),
.B2(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_106),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_115),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_102),
.B(n_119),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_188),
.B(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_3),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_119),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_83),
.B1(n_93),
.B2(n_100),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_185),
.A2(n_132),
.B1(n_135),
.B2(n_129),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_120),
.B1(n_109),
.B2(n_100),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_126),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_196),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_201),
.B(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_137),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_193),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_129),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_199),
.B1(n_180),
.B2(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_130),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_204),
.C(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_130),
.C(n_139),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_206),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_146),
.B1(n_139),
.B2(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_203),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_37),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_36),
.B1(n_31),
.B2(n_29),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_212),
.B1(n_217),
.B2(n_156),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_11),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_143),
.B1(n_29),
.B2(n_2),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_185),
.B1(n_217),
.B2(n_166),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_218),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_177),
.Y(n_216)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_227),
.B1(n_165),
.B2(n_179),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_160),
.B1(n_158),
.B2(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_231),
.B1(n_208),
.B2(n_181),
.Y(n_255)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_164),
.Y(n_233)
);

NOR4xp25_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_186),
.C(n_171),
.D(n_169),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_191),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_174),
.C(n_173),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_189),
.C(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_208),
.B(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_181),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_248),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_232),
.B(n_220),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_193),
.Y(n_248)
);

XOR2x1_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_189),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_249),
.A2(n_259),
.B1(n_261),
.B2(n_220),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_251),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_214),
.Y(n_251)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_229),
.B1(n_225),
.B2(n_208),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_229),
.B1(n_228),
.B2(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_256),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_198),
.C(n_165),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_260),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_188),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_155),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_155),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_265),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_277),
.B1(n_240),
.B2(n_253),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_219),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_206),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_253),
.B(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_261),
.C(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_275),
.C(n_273),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_251),
.C(n_224),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_285),
.C(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_223),
.C(n_256),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_230),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_241),
.B1(n_242),
.B2(n_230),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_273),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_264),
.B(n_268),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_280),
.B(n_161),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_274),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_277),
.B1(n_291),
.B2(n_283),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_274),
.B(n_262),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_287),
.B1(n_284),
.B2(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_294),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_306),
.B(n_308),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_295),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_294),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_234),
.A3(n_161),
.B(n_8),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_13),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_316),
.B1(n_311),
.B2(n_8),
.C(n_16),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_308),
.A3(n_307),
.B1(n_234),
.B2(n_16),
.C1(n_5),
.C2(n_9),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_5),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_307),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_17),
.Y(n_321)
);


endmodule