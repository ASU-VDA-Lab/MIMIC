module real_jpeg_12860_n_19 (n_17, n_8, n_0, n_93, n_2, n_10, n_9, n_12, n_92, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_94, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_93;
input n_2;
input n_10;
input n_9;
input n_12;
input n_92;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_94;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_0),
.A2(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_0),
.B(n_9),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_4),
.B1(n_25),
.B2(n_49),
.Y(n_48)
);

AOI221xp5_ASAP7_75t_L g50 ( 
.A1(n_0),
.A2(n_1),
.B1(n_25),
.B2(n_51),
.C(n_52),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_0),
.A2(n_18),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_92),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_57),
.B1(n_59),
.B2(n_70),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_21),
.B1(n_54),
.B2(n_55),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_8),
.A2(n_54),
.B1(n_74),
.B2(n_84),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_9),
.B(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_9),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_12),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_93),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_94),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

AOI221xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_56),
.B1(n_73),
.B2(n_85),
.C(n_89),
.Y(n_19)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

OAI211xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_36),
.C(n_45),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_35),
.C(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_34),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_35),
.A2(n_42),
.B(n_78),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_37),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_77),
.C(n_83),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_61),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_66),
.B(n_69),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);


endmodule