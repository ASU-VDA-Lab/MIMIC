module real_aes_6830_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_1), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_1), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_2), .A2(n_134), .B(n_139), .C(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_3), .A2(n_129), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g498 ( .A(n_4), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_5), .B(n_167), .Y(n_233) );
AOI21xp33_ASAP7_75t_L g505 ( .A1(n_6), .A2(n_129), .B(n_506), .Y(n_505) );
AND2x6_ASAP7_75t_L g134 ( .A(n_7), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_8), .A2(n_264), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g146 ( .A(n_9), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_10), .B(n_43), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_11), .A2(n_33), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_11), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_12), .B(n_144), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_13), .B(n_191), .Y(n_477) );
INVx1_ASAP7_75t_L g510 ( .A(n_14), .Y(n_510) );
INVx1_ASAP7_75t_L g127 ( .A(n_15), .Y(n_127) );
INVx1_ASAP7_75t_L g489 ( .A(n_16), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_17), .A2(n_147), .B(n_161), .C(n_165), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_18), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_19), .B(n_468), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_20), .B(n_129), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_21), .B(n_273), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_22), .A2(n_191), .B(n_192), .C(n_194), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_23), .B(n_167), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_24), .B(n_144), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_25), .A2(n_163), .B(n_165), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_26), .B(n_144), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_27), .Y(n_215) );
INVx1_ASAP7_75t_L g203 ( .A(n_28), .Y(n_203) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_29), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_30), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_31), .B(n_144), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_32), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g453 ( .A(n_33), .Y(n_453) );
INVx1_ASAP7_75t_L g269 ( .A(n_34), .Y(n_269) );
INVx1_ASAP7_75t_L g518 ( .A(n_35), .Y(n_518) );
INVx2_ASAP7_75t_L g132 ( .A(n_36), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_37), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_38), .A2(n_191), .B(n_229), .C(n_231), .Y(n_228) );
INVxp67_ASAP7_75t_L g270 ( .A(n_39), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_40), .A2(n_139), .B(n_202), .C(n_208), .Y(n_201) );
CKINVDCx14_ASAP7_75t_R g227 ( .A(n_41), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_42), .A2(n_134), .B(n_139), .C(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g517 ( .A(n_44), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_45), .A2(n_143), .B(n_145), .C(n_148), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_46), .B(n_144), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_47), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_48), .Y(n_266) );
INVx1_ASAP7_75t_L g189 ( .A(n_49), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_50), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_51), .B(n_129), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_52), .A2(n_139), .B1(n_194), .B2(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_53), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_54), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g137 ( .A(n_55), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_56), .A2(n_143), .B(n_231), .C(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_57), .Y(n_555) );
INVx1_ASAP7_75t_L g507 ( .A(n_58), .Y(n_507) );
INVx1_ASAP7_75t_L g135 ( .A(n_59), .Y(n_135) );
INVx1_ASAP7_75t_L g126 ( .A(n_60), .Y(n_126) );
INVx1_ASAP7_75t_SL g230 ( .A(n_61), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_62), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_63), .B(n_167), .Y(n_196) );
INVx1_ASAP7_75t_L g218 ( .A(n_64), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_SL g526 ( .A1(n_65), .A2(n_231), .B(n_468), .C(n_527), .Y(n_526) );
INVxp67_ASAP7_75t_L g528 ( .A(n_66), .Y(n_528) );
INVx1_ASAP7_75t_L g442 ( .A(n_67), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_68), .A2(n_129), .B(n_136), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_69), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_70), .A2(n_129), .B(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_71), .Y(n_521) );
INVx1_ASAP7_75t_L g549 ( .A(n_72), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_73), .A2(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g159 ( .A(n_74), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_75), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_76), .A2(n_77), .B1(n_430), .B2(n_431), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_76), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_77), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_78), .A2(n_134), .B(n_139), .C(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_SL g444 ( .A1(n_79), .A2(n_107), .B1(n_445), .B2(n_739), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_80), .A2(n_129), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g162 ( .A(n_81), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_82), .B(n_204), .Y(n_466) );
INVx2_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
INVx1_ASAP7_75t_L g178 ( .A(n_84), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_85), .B(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_86), .A2(n_134), .B(n_139), .C(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g106 ( .A(n_87), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g737 ( .A(n_87), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_88), .A2(n_139), .B(n_217), .C(n_220), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_89), .A2(n_91), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_89), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_90), .B(n_123), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_91), .A2(n_104), .B1(n_436), .B2(n_443), .C1(n_742), .C2(n_746), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_91), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_92), .A2(n_134), .B(n_139), .C(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_93), .Y(n_481) );
INVx1_ASAP7_75t_L g525 ( .A(n_94), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_95), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_96), .B(n_204), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_97), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_98), .B(n_152), .Y(n_490) );
INVx2_ASAP7_75t_L g193 ( .A(n_99), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_100), .B(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_101), .A2(n_447), .B1(n_448), .B2(n_449), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_101), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_102), .A2(n_129), .B(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_111), .B(n_433), .Y(n_104) );
INVx1_ASAP7_75t_SL g745 ( .A(n_105), .Y(n_745) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_106), .Y(n_435) );
BUFx2_ASAP7_75t_L g748 ( .A(n_106), .Y(n_748) );
NOR2x2_ASAP7_75t_L g741 ( .A(n_107), .B(n_737), .Y(n_741) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_115), .B1(n_116), .B2(n_432), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_112), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_113), .B(n_172), .Y(n_501) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
XOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_429), .Y(n_116) );
INVx2_ASAP7_75t_L g738 ( .A(n_117), .Y(n_738) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_359), .Y(n_117) );
NAND5xp2_ASAP7_75t_L g118 ( .A(n_119), .B(n_274), .C(n_306), .D(n_323), .E(n_346), .Y(n_118) );
AOI221xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_197), .B1(n_234), .B2(n_238), .C(n_242), .Y(n_119) );
INVx1_ASAP7_75t_L g386 ( .A(n_120), .Y(n_386) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_169), .Y(n_120) );
AND3x2_ASAP7_75t_L g361 ( .A(n_121), .B(n_171), .C(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_154), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_122), .B(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g249 ( .A(n_122), .Y(n_249) );
AND2x2_ASAP7_75t_L g253 ( .A(n_122), .B(n_185), .Y(n_253) );
INVx2_ASAP7_75t_L g283 ( .A(n_122), .Y(n_283) );
OR2x2_ASAP7_75t_L g294 ( .A(n_122), .B(n_186), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_122), .B(n_170), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_122), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g373 ( .A(n_122), .B(n_186), .Y(n_373) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_151), .Y(n_122) );
INVx1_ASAP7_75t_L g172 ( .A(n_123), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_123), .A2(n_175), .B(n_200), .C(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g223 ( .A(n_123), .Y(n_223) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_123), .A2(n_484), .B(n_490), .Y(n_483) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_L g153 ( .A(n_124), .B(n_125), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx2_ASAP7_75t_L g264 ( .A(n_129), .Y(n_264) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_130), .B(n_134), .Y(n_175) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx1_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx1_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_133), .Y(n_144) );
INVx3_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
INVx1_ASAP7_75t_L g468 ( .A(n_133), .Y(n_468) );
INVx4_ASAP7_75t_SL g150 ( .A(n_134), .Y(n_150) );
BUFx3_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_138), .B(n_142), .C(n_150), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_SL g158 ( .A1(n_138), .A2(n_150), .B(n_159), .C(n_160), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_138), .A2(n_150), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_138), .A2(n_150), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_138), .A2(n_150), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_138), .A2(n_150), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_138), .A2(n_150), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_138), .A2(n_150), .B(n_525), .C(n_526), .Y(n_524) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g149 ( .A(n_140), .Y(n_149) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_140), .Y(n_232) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx5_ASAP7_75t_L g204 ( .A(n_147), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_147), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_147), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_150), .A2(n_175), .B1(n_515), .B2(n_519), .Y(n_514) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_152), .Y(n_156) );
INVx4_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_523), .B(n_529), .Y(n_522) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g261 ( .A(n_153), .Y(n_261) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_154), .Y(n_252) );
AND2x2_ASAP7_75t_L g314 ( .A(n_154), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_154), .B(n_170), .Y(n_333) );
INVx1_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
OR2x2_ASAP7_75t_L g241 ( .A(n_155), .B(n_170), .Y(n_241) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_155), .Y(n_248) );
AND2x2_ASAP7_75t_L g300 ( .A(n_155), .B(n_186), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_155), .B(n_169), .C(n_283), .Y(n_325) );
AND2x2_ASAP7_75t_L g390 ( .A(n_155), .B(n_171), .Y(n_390) );
AND2x2_ASAP7_75t_L g424 ( .A(n_155), .B(n_170), .Y(n_424) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_166), .Y(n_155) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_156), .A2(n_187), .B(n_196), .Y(n_186) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_156), .A2(n_225), .B(n_233), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_163), .B(n_193), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_163), .A2(n_204), .B1(n_269), .B2(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_163), .B(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g516 ( .A1(n_164), .A2(n_180), .B1(n_517), .B2(n_518), .Y(n_516) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_167), .A2(n_505), .B(n_511), .Y(n_504) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_168), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_168), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_168), .A2(n_214), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_SL g469 ( .A(n_168), .B(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_185), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_170), .B(n_283), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_170), .B(n_314), .Y(n_322) );
AND2x2_ASAP7_75t_L g372 ( .A(n_170), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g400 ( .A(n_170), .Y(n_400) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g307 ( .A(n_171), .B(n_300), .Y(n_307) );
BUFx3_ASAP7_75t_L g339 ( .A(n_171), .Y(n_339) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_183), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_172), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_172), .B(n_555), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_175), .A2(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_175), .A2(n_495), .B(n_496), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_175), .A2(n_549), .B(n_550), .Y(n_548) );
O2A1O1Ixp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_181), .C(n_182), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_179), .A2(n_182), .B(n_218), .C(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_182), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_182), .A2(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g315 ( .A(n_185), .Y(n_315) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_191), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g500 ( .A(n_194), .Y(n_500) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_197), .A2(n_375), .B1(n_377), .B2(n_378), .Y(n_374) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_211), .Y(n_197) );
AND2x2_ASAP7_75t_L g234 ( .A(n_198), .B(n_235), .Y(n_234) );
INVx3_ASAP7_75t_SL g245 ( .A(n_198), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_198), .B(n_278), .Y(n_310) );
OR2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_212), .Y(n_329) );
AND2x2_ASAP7_75t_L g334 ( .A(n_198), .B(n_286), .Y(n_334) );
AND2x2_ASAP7_75t_L g337 ( .A(n_198), .B(n_279), .Y(n_337) );
AND2x2_ASAP7_75t_L g349 ( .A(n_198), .B(n_224), .Y(n_349) );
AND2x2_ASAP7_75t_L g365 ( .A(n_198), .B(n_213), .Y(n_365) );
AND2x4_ASAP7_75t_L g368 ( .A(n_198), .B(n_236), .Y(n_368) );
OR2x2_ASAP7_75t_L g385 ( .A(n_198), .B(n_321), .Y(n_385) );
OR2x2_ASAP7_75t_L g416 ( .A(n_198), .B(n_258), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_198), .B(n_344), .Y(n_418) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_204), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_207), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g292 ( .A(n_211), .B(n_256), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_211), .B(n_279), .Y(n_411) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_224), .Y(n_211) );
AND2x2_ASAP7_75t_L g244 ( .A(n_212), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g278 ( .A(n_212), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g286 ( .A(n_212), .B(n_258), .Y(n_286) );
AND2x2_ASAP7_75t_L g304 ( .A(n_212), .B(n_236), .Y(n_304) );
OR2x2_ASAP7_75t_L g321 ( .A(n_212), .B(n_279), .Y(n_321) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
AND2x2_ASAP7_75t_L g344 ( .A(n_213), .B(n_224), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx1_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_223), .A2(n_473), .B(n_480), .Y(n_472) );
INVx2_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
INVx1_ASAP7_75t_L g356 ( .A(n_224), .Y(n_356) );
AND2x2_ASAP7_75t_L g406 ( .A(n_224), .B(n_245), .Y(n_406) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_232), .Y(n_478) );
AND2x2_ASAP7_75t_L g255 ( .A(n_235), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g290 ( .A(n_235), .B(n_245), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_235), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AND2x2_ASAP7_75t_L g277 ( .A(n_236), .B(n_245), .Y(n_277) );
OR2x2_ASAP7_75t_L g393 ( .A(n_237), .B(n_367), .Y(n_393) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_240), .B(n_373), .Y(n_379) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OAI32xp33_ASAP7_75t_L g335 ( .A1(n_241), .A2(n_336), .A3(n_338), .B1(n_340), .B2(n_341), .Y(n_335) );
OR2x2_ASAP7_75t_L g352 ( .A(n_241), .B(n_294), .Y(n_352) );
OAI21xp33_ASAP7_75t_SL g377 ( .A1(n_241), .A2(n_251), .B(n_282), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .B1(n_251), .B2(n_254), .Y(n_242) );
INVxp33_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_244), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_245), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g403 ( .A(n_245), .B(n_344), .Y(n_403) );
OR2x2_ASAP7_75t_L g427 ( .A(n_245), .B(n_321), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_246), .A2(n_309), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g287 ( .A(n_248), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_248), .B(n_253), .Y(n_305) );
AND2x2_ASAP7_75t_L g327 ( .A(n_249), .B(n_300), .Y(n_327) );
INVx1_ASAP7_75t_L g340 ( .A(n_249), .Y(n_340) );
OR2x2_ASAP7_75t_L g345 ( .A(n_249), .B(n_279), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_252), .B(n_294), .Y(n_293) );
OAI22xp33_ASAP7_75t_L g275 ( .A1(n_253), .A2(n_276), .B1(n_281), .B2(n_285), .Y(n_275) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_256), .A2(n_318), .B1(n_325), .B2(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g402 ( .A(n_256), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_258), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g421 ( .A(n_258), .B(n_304), .Y(n_421) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B(n_271), .Y(n_258) );
INVx1_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_259), .A2(n_548), .B(n_554), .Y(n_547) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_260), .A2(n_463), .B(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_261), .A2(n_494), .B(n_501), .Y(n_493) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_261), .A2(n_514), .B(n_520), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_261), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_263), .A2(n_272), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_287), .B1(n_288), .B2(n_293), .C(n_295), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_277), .B(n_279), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_277), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_278), .A2(n_384), .B(n_385), .C(n_386), .Y(n_383) );
AND2x2_ASAP7_75t_L g388 ( .A(n_278), .B(n_368), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_SL g426 ( .A1(n_278), .A2(n_367), .B(n_427), .C(n_428), .Y(n_426) );
BUFx3_ASAP7_75t_L g318 ( .A(n_279), .Y(n_318) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_282), .B(n_339), .Y(n_382) );
AOI211xp5_ASAP7_75t_L g401 ( .A1(n_282), .A2(n_402), .B(n_404), .C(n_410), .Y(n_401) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVxp67_ASAP7_75t_L g362 ( .A(n_284), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_286), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AOI211xp5_ASAP7_75t_L g306 ( .A1(n_290), .A2(n_307), .B(n_308), .C(n_316), .Y(n_306) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g391 ( .A(n_294), .Y(n_391) );
OR2x2_ASAP7_75t_L g408 ( .A(n_294), .B(n_338), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B1(n_302), .B2(n_305), .Y(n_295) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_297), .A2(n_309), .B1(n_310), .B2(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
OR2x2_ASAP7_75t_L g395 ( .A(n_299), .B(n_339), .Y(n_395) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g350 ( .A(n_300), .B(n_340), .Y(n_350) );
INVx1_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_304), .B(n_318), .Y(n_366) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_314), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g423 ( .A(n_315), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B(n_322), .Y(n_316) );
INVx1_ASAP7_75t_L g353 ( .A(n_317), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_318), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_318), .B(n_349), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_318), .B(n_344), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_318), .B(n_365), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_318), .A2(n_328), .B(n_368), .C(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AOI221xp5_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_328), .B1(n_330), .B2(n_334), .C(n_335), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_332), .B(n_340), .Y(n_414) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g425 ( .A1(n_334), .A2(n_349), .B(n_351), .C(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_337), .B(n_344), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_338), .B(n_391), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
INVxp33_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AOI21xp33_ASAP7_75t_SL g354 ( .A1(n_343), .A2(n_355), .B(n_357), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_343), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_344), .B(n_398), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_350), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
NAND5xp2_ASAP7_75t_L g359 ( .A(n_360), .B(n_387), .C(n_401), .D(n_412), .E(n_425), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_370), .C(n_383), .Y(n_360) );
INVx2_ASAP7_75t_SL g407 ( .A(n_361), .Y(n_407) );
NAND4xp25_ASAP7_75t_SL g363 ( .A(n_364), .B(n_366), .C(n_367), .D(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_369), .A2(n_371), .B(n_374), .C(n_380), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_372), .A2(n_413), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI221xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B1(n_392), .B2(n_394), .C(n_396), .Y(n_387) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_418), .B1(n_420), .B2(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_SL g744 ( .A(n_439), .B(n_441), .Y(n_744) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_439), .A2(n_440), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
XOR2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_735), .B1(n_736), .B2(n_738), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_704), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_597), .C(n_670), .Y(n_457) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_491), .B(n_530), .C(n_581), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_471), .Y(n_460) );
AND2x2_ASAP7_75t_L g546 ( .A(n_461), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g564 ( .A(n_461), .Y(n_564) );
INVx2_ASAP7_75t_L g579 ( .A(n_461), .Y(n_579) );
INVx1_ASAP7_75t_L g609 ( .A(n_461), .Y(n_609) );
AND2x2_ASAP7_75t_L g659 ( .A(n_461), .B(n_580), .Y(n_659) );
AOI32xp33_ASAP7_75t_L g686 ( .A1(n_461), .A2(n_614), .A3(n_687), .B1(n_689), .B2(n_690), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_461), .B(n_536), .Y(n_692) );
AND2x2_ASAP7_75t_L g719 ( .A(n_461), .B(n_562), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_461), .B(n_728), .Y(n_727) );
OR2x6_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
AND2x2_ASAP7_75t_L g608 ( .A(n_471), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g630 ( .A(n_471), .Y(n_630) );
AND2x2_ASAP7_75t_L g715 ( .A(n_471), .B(n_546), .Y(n_715) );
AND2x2_ASAP7_75t_L g718 ( .A(n_471), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
INVx2_ASAP7_75t_L g538 ( .A(n_472), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_472), .B(n_562), .Y(n_568) );
AND2x2_ASAP7_75t_L g578 ( .A(n_472), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g614 ( .A(n_472), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_479), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_478), .Y(n_475) );
AND2x2_ASAP7_75t_L g556 ( .A(n_482), .B(n_538), .Y(n_556) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
AND2x2_ASAP7_75t_L g580 ( .A(n_483), .B(n_562), .Y(n_580) );
AND2x2_ASAP7_75t_L g649 ( .A(n_483), .B(n_547), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
OR2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_513), .Y(n_544) );
INVx1_ASAP7_75t_L g622 ( .A(n_492), .Y(n_622) );
AND2x2_ASAP7_75t_L g636 ( .A(n_492), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_492), .B(n_512), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_492), .B(n_634), .Y(n_688) );
AND2x2_ASAP7_75t_L g696 ( .A(n_492), .B(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AND2x2_ASAP7_75t_L g603 ( .A(n_493), .B(n_513), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_502), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g730 ( .A(n_502), .Y(n_730) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_503), .B(n_574), .Y(n_596) );
OR2x2_ASAP7_75t_L g625 ( .A(n_503), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g657 ( .A(n_503), .B(n_637), .Y(n_657) );
INVx1_ASAP7_75t_SL g677 ( .A(n_503), .Y(n_677) );
AND2x2_ASAP7_75t_L g681 ( .A(n_503), .B(n_543), .Y(n_681) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_SL g535 ( .A(n_504), .B(n_512), .Y(n_535) );
AND2x2_ASAP7_75t_L g542 ( .A(n_504), .B(n_522), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_504), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_566), .Y(n_584) );
INVx1_ASAP7_75t_SL g591 ( .A(n_504), .Y(n_591) );
BUFx2_ASAP7_75t_L g602 ( .A(n_504), .Y(n_602) );
AND2x2_ASAP7_75t_L g618 ( .A(n_504), .B(n_534), .Y(n_618) );
AND2x2_ASAP7_75t_L g633 ( .A(n_504), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g697 ( .A(n_504), .B(n_513), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_512), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g621 ( .A(n_512), .B(n_622), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_512), .A2(n_639), .B1(n_642), .B2(n_645), .C(n_650), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_512), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
INVx3_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
BUFx2_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
AND2x2_ASAP7_75t_L g590 ( .A(n_522), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
OR2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_566), .Y(n_626) );
INVx3_ASAP7_75t_L g634 ( .A(n_522), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_522), .B(n_566), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_536), .B1(n_540), .B2(n_545), .C(n_557), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_533), .B(n_606), .Y(n_731) );
OR2x2_ASAP7_75t_L g734 ( .A(n_533), .B(n_565), .Y(n_734) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_534), .A2(n_558), .B1(n_565), .B2(n_567), .C(n_570), .Y(n_557) );
AND2x2_ASAP7_75t_L g574 ( .A(n_534), .B(n_566), .Y(n_574) );
AND2x2_ASAP7_75t_L g582 ( .A(n_534), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_534), .B(n_590), .Y(n_589) );
NAND2x1_ASAP7_75t_L g632 ( .A(n_534), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g684 ( .A(n_534), .B(n_626), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_536), .A2(n_644), .B1(n_673), .B2(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AOI322xp5_ASAP7_75t_L g581 ( .A1(n_537), .A2(n_546), .A3(n_582), .B1(n_585), .B2(n_588), .C1(n_592), .C2(n_595), .Y(n_581) );
OR2x2_ASAP7_75t_L g593 ( .A(n_537), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_538), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g572 ( .A(n_538), .B(n_547), .Y(n_572) );
INVx1_ASAP7_75t_L g587 ( .A(n_538), .Y(n_587) );
AND2x2_ASAP7_75t_L g653 ( .A(n_538), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g563 ( .A(n_539), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g654 ( .A(n_539), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_539), .B(n_562), .Y(n_728) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_543), .B(n_677), .Y(n_676) );
INVx3_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g628 ( .A(n_544), .B(n_575), .Y(n_628) );
OR2x2_ASAP7_75t_L g725 ( .A(n_544), .B(n_576), .Y(n_725) );
INVx1_ASAP7_75t_L g706 ( .A(n_545), .Y(n_706) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
INVx4_ASAP7_75t_L g594 ( .A(n_546), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_546), .B(n_613), .Y(n_619) );
INVx2_ASAP7_75t_L g562 ( .A(n_547), .Y(n_562) );
INVx1_ASAP7_75t_L g644 ( .A(n_556), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_556), .B(n_616), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_558), .A2(n_632), .B(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g616 ( .A(n_562), .Y(n_616) );
INVx1_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
INVx1_ASAP7_75t_L g569 ( .A(n_563), .Y(n_569) );
AND2x2_ASAP7_75t_L g571 ( .A(n_563), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g667 ( .A(n_564), .B(n_653), .Y(n_667) );
AND2x2_ASAP7_75t_L g689 ( .A(n_564), .B(n_649), .Y(n_689) );
BUFx2_ASAP7_75t_L g641 ( .A(n_566), .Y(n_641) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AOI32xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .A3(n_574), .B1(n_575), .B2(n_577), .Y(n_570) );
INVx1_ASAP7_75t_L g651 ( .A(n_571), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_571), .A2(n_699), .B1(n_700), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_574), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_574), .B(n_633), .Y(n_674) );
AND2x2_ASAP7_75t_L g721 ( .A(n_574), .B(n_606), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_575), .B(n_622), .Y(n_669) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g722 ( .A(n_577), .Y(n_722) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g647 ( .A(n_578), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_580), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g694 ( .A(n_580), .B(n_614), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_580), .B(n_609), .Y(n_701) );
INVx1_ASAP7_75t_SL g683 ( .A(n_582), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_583), .B(n_634), .Y(n_661) );
NOR4xp25_ASAP7_75t_L g707 ( .A(n_583), .B(n_606), .C(n_708), .D(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_584), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_L g664 ( .A(n_587), .Y(n_664) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_590), .A2(n_681), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g606 ( .A(n_591), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g655 ( .A(n_594), .Y(n_655) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND4xp25_ASAP7_75t_SL g597 ( .A(n_598), .B(n_623), .C(n_638), .D(n_658), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_604), .B(n_608), .C(n_610), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g690 ( .A(n_603), .B(n_633), .Y(n_690) );
AND2x2_ASAP7_75t_L g699 ( .A(n_603), .B(n_677), .Y(n_699) );
INVx3_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_606), .B(n_641), .Y(n_703) );
AND2x2_ASAP7_75t_L g615 ( .A(n_609), .B(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_617), .B1(n_619), .B2(n_620), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
AND2x2_ASAP7_75t_L g713 ( .A(n_613), .B(n_659), .Y(n_713) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_615), .B(n_664), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_616), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_629), .C(n_631), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_624), .A2(n_659), .B1(n_660), .B2(n_662), .C(n_665), .Y(n_658) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_632), .A2(n_717), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_633), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_641), .B(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g671 ( .A(n_643), .Y(n_671) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_646), .A2(n_666), .B1(n_668), .B2(n_669), .Y(n_665) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_655), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_666), .A2(n_692), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g711 ( .A(n_668), .Y(n_711) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_672), .B(n_678), .C(n_698), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B(n_682), .C(n_691), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_685), .C(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g710 ( .A(n_688), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_689), .A2(n_715), .B(n_733), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B(n_695), .Y(n_691) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_701), .A2(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_716), .C(n_729), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_712), .C(n_714), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
CKINVDCx14_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
NAND2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
endmodule