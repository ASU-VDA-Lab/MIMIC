module fake_jpeg_12673_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_61),
.B(n_62),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_71),
.B(n_98),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_13),
.Y(n_114)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_89),
.Y(n_128)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g160 ( 
.A(n_92),
.Y(n_160)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_8),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_35),
.B1(n_27),
.B2(n_50),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_102),
.Y(n_149)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_49),
.Y(n_153)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_54),
.A2(n_19),
.B1(n_30),
.B2(n_48),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_116),
.B(n_104),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_51),
.B1(n_37),
.B2(n_48),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_109),
.A2(n_119),
.B1(n_122),
.B2(n_136),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_167),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_69),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_85),
.A2(n_51),
.B1(n_46),
.B2(n_48),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_127),
.A2(n_133),
.B1(n_141),
.B2(n_159),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_46),
.B1(n_33),
.B2(n_28),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_52),
.B1(n_24),
.B2(n_33),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_52),
.B1(n_34),
.B2(n_36),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_146),
.B1(n_148),
.B2(n_45),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_90),
.B1(n_102),
.B2(n_63),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_53),
.A2(n_52),
.B1(n_34),
.B2(n_36),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_68),
.A2(n_52),
.B1(n_47),
.B2(n_96),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_10),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_39),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_155),
.B(n_156),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_57),
.B(n_39),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_42),
.B1(n_38),
.B2(n_50),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_64),
.A2(n_49),
.B1(n_42),
.B2(n_35),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_91),
.B1(n_83),
.B2(n_100),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_70),
.A2(n_47),
.B1(n_19),
.B2(n_45),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_78),
.B(n_0),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_168),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_169),
.A2(n_183),
.B1(n_192),
.B2(n_227),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_171),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_173),
.A2(n_188),
.B1(n_212),
.B2(n_221),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_175),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_92),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_176),
.B(n_181),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_103),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_177),
.B(n_217),
.Y(n_248)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g273 ( 
.A1(n_179),
.A2(n_121),
.B(n_144),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_105),
.Y(n_180)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_15),
.Y(n_181)
);

BUFx6f_ASAP7_75t_SL g182 ( 
.A(n_165),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_72),
.B1(n_73),
.B2(n_81),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_183),
.A2(n_189),
.B(n_128),
.Y(n_250)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_81),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_186),
.B(n_187),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_147),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_106),
.A2(n_76),
.B1(n_86),
.B2(n_88),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_93),
.B1(n_80),
.B2(n_45),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_196),
.C(n_215),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_8),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_204),
.Y(n_265)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_45),
.B1(n_8),
.B2(n_3),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_206),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_276)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_207),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_210),
.B1(n_214),
.B2(n_216),
.Y(n_231)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_209),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_211),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_107),
.A2(n_45),
.B1(n_12),
.B2(n_3),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_213),
.Y(n_280)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_108),
.B(n_18),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_138),
.Y(n_271)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_126),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_108),
.A2(n_7),
.B1(n_15),
.B2(n_3),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_134),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_142),
.A2(n_7),
.B1(n_15),
.B2(n_4),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_162),
.A2(n_6),
.B1(n_14),
.B2(n_4),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_225),
.A2(n_0),
.B1(n_2),
.B2(n_224),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_227),
.B1(n_157),
.B2(n_164),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_142),
.A2(n_6),
.B1(n_14),
.B2(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_118),
.B(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_128),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_152),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_238),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_111),
.B(n_145),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_234),
.A2(n_214),
.B(n_208),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_152),
.B1(n_147),
.B2(n_135),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_235),
.A2(n_249),
.B1(n_261),
.B2(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_135),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_162),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_268),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_200),
.A2(n_166),
.B1(n_132),
.B2(n_131),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_216),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_190),
.A2(n_166),
.B1(n_131),
.B2(n_126),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_177),
.B(n_160),
.C(n_128),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_193),
.C(n_184),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_170),
.B(n_121),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_207),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_190),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_254),
.B1(n_246),
.B2(n_242),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_277),
.B1(n_180),
.B2(n_220),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_188),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_225),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_169),
.A2(n_0),
.B1(n_2),
.B2(n_189),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_219),
.B(n_2),
.CI(n_189),
.CON(n_282),
.SN(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_174),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_284),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_182),
.C(n_178),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_285),
.B(n_314),
.C(n_316),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_286),
.B(n_288),
.Y(n_367)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_287),
.Y(n_372)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_294),
.A2(n_299),
.B1(n_301),
.B2(n_315),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_171),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_235),
.B1(n_232),
.B2(n_261),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g301 ( 
.A1(n_250),
.A2(n_198),
.B(n_197),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_272),
.B(n_205),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_303),
.B(n_320),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_230),
.A2(n_168),
.B1(n_226),
.B2(n_210),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_306),
.A2(n_293),
.B1(n_324),
.B2(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_209),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_248),
.A2(n_204),
.B(n_203),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_310),
.A2(n_297),
.B(n_312),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_243),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_311),
.B(n_312),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_248),
.B(n_239),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_313),
.A2(n_327),
.B(n_330),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_250),
.A2(n_2),
.B1(n_230),
.B2(n_258),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_238),
.C(n_259),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_274),
.C(n_248),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_250),
.A2(n_279),
.B1(n_282),
.B2(n_252),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_318),
.A2(n_315),
.B1(n_294),
.B2(n_295),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_252),
.B(n_264),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_323),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_240),
.B(n_269),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_237),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_326),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_322),
.A2(n_254),
.B1(n_246),
.B2(n_242),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_257),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_324),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_254),
.Y(n_325)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_263),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_276),
.A2(n_244),
.B(n_269),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_233),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_328),
.B(n_329),
.Y(n_359)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_236),
.A2(n_263),
.B(n_270),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_253),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_236),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_257),
.B(n_231),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_346),
.B1(n_352),
.B2(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_351),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_318),
.A2(n_266),
.B1(n_270),
.B2(n_253),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_280),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_290),
.A2(n_266),
.B1(n_265),
.B2(n_233),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_300),
.B(n_309),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_290),
.A2(n_266),
.B1(n_265),
.B2(n_255),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_295),
.A2(n_255),
.B1(n_246),
.B2(n_245),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_355),
.A2(n_369),
.B1(n_354),
.B2(n_352),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_301),
.B1(n_329),
.B2(n_305),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_241),
.B1(n_297),
.B2(n_311),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_362),
.A2(n_371),
.B1(n_301),
.B2(n_285),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_326),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_366),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_299),
.A2(n_241),
.B1(n_301),
.B2(n_283),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_309),
.B1(n_327),
.B2(n_316),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_331),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_373),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_304),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_360),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_380),
.B1(n_383),
.B2(n_385),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_301),
.B1(n_300),
.B2(n_307),
.Y(n_380)
);

AOI21xp33_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_307),
.B(n_330),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_381),
.B(n_335),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_314),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_401),
.C(n_405),
.Y(n_419)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_371),
.A2(n_317),
.B1(n_302),
.B2(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_344),
.A2(n_310),
.B(n_289),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_392),
.A2(n_393),
.B(n_394),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_308),
.B(n_325),
.Y(n_393)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_365),
.A2(n_293),
.B(n_291),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_338),
.A2(n_341),
.B1(n_334),
.B2(n_353),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_399),
.B1(n_337),
.B2(n_356),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_342),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_406),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_397),
.A2(n_400),
.B(n_404),
.Y(n_416)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_338),
.A2(n_334),
.B1(n_370),
.B2(n_335),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_343),
.A2(n_336),
.B(n_362),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_364),
.A2(n_373),
.B(n_359),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_367),
.C(n_359),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_350),
.A2(n_349),
.B(n_369),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_350),
.A2(n_348),
.B(n_368),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g412 ( 
.A1(n_407),
.A2(n_368),
.B(n_356),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_355),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_376),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_413),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_386),
.A2(n_357),
.B1(n_348),
.B2(n_337),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_411),
.A2(n_428),
.B1(n_429),
.B2(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_412),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_418),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_438),
.C(n_401),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_421),
.A2(n_422),
.B1(n_427),
.B2(n_432),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_361),
.B1(n_358),
.B2(n_372),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_377),
.B(n_361),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_425),
.B(n_407),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_358),
.B1(n_372),
.B2(n_333),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_386),
.A2(n_333),
.B1(n_372),
.B2(n_339),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_388),
.A2(n_397),
.B1(n_396),
.B2(n_405),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_430),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_395),
.A2(n_380),
.B1(n_389),
.B2(n_405),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_376),
.B1(n_385),
.B2(n_408),
.Y(n_433)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_433),
.Y(n_440)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_374),
.Y(n_435)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_436),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_382),
.B(n_401),
.C(n_375),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_382),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_420),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_442),
.B(n_444),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_393),
.C(n_394),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_448),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_404),
.Y(n_444)
);

AOI211xp5_ASAP7_75t_L g471 ( 
.A1(n_445),
.A2(n_437),
.B(n_412),
.C(n_416),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_377),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_446),
.B(n_459),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_425),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_416),
.A2(n_400),
.B(n_406),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_457),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_455),
.A2(n_463),
.B1(n_420),
.B2(n_432),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_391),
.Y(n_456)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_464),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_379),
.C(n_381),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_384),
.C(n_387),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_460),
.B(n_461),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_398),
.C(n_402),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_429),
.A2(n_403),
.B1(n_410),
.B2(n_411),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_470),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_479),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_463),
.A2(n_413),
.B1(n_422),
.B2(n_436),
.Y(n_469)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_444),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_477),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_428),
.B1(n_423),
.B2(n_424),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_472),
.A2(n_480),
.B1(n_481),
.B2(n_439),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_415),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_483),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_434),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_434),
.B1(n_423),
.B2(n_424),
.Y(n_479)
);

INVx11_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_450),
.A2(n_415),
.B1(n_426),
.B2(n_431),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_459),
.B(n_426),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_470),
.C(n_466),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_487),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_460),
.C(n_443),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_461),
.C(n_440),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_492),
.C(n_483),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_440),
.C(n_449),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_465),
.A2(n_462),
.B1(n_452),
.B2(n_439),
.Y(n_493)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_484),
.A2(n_462),
.B(n_456),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_476),
.B1(n_430),
.B2(n_435),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_467),
.B(n_454),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_498),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_476),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_465),
.A2(n_454),
.B1(n_447),
.B2(n_431),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_447),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_481),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_500),
.A2(n_478),
.B1(n_480),
.B2(n_472),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_493),
.B1(n_498),
.B2(n_496),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_508),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_489),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_482),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_500),
.A2(n_474),
.B(n_471),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_510),
.B(n_511),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_474),
.C(n_477),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_491),
.C(n_489),
.Y(n_511)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_512),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_514),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_513),
.A2(n_490),
.B1(n_488),
.B2(n_492),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_523),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_505),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_508),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_509),
.A2(n_499),
.B(n_504),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_506),
.B(n_511),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_502),
.A2(n_499),
.B1(n_510),
.B2(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_524),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_527),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_519),
.B(n_507),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_521),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_524),
.B(n_516),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_529),
.A2(n_520),
.B(n_526),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_533),
.B(n_530),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_515),
.C(n_523),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_535),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_517),
.B(n_505),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_518),
.Y(n_538)
);


endmodule