module fake_netlist_6_3253_n_2078 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2078);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2078;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_0),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_61),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_31),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_27),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_38),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_55),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_161),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_28),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_0),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_37),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_86),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_56),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_61),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_27),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_154),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_59),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_128),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_47),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_94),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_55),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_155),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_45),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_140),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_58),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_111),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_76),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_7),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_58),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_64),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_82),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_96),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_181),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_172),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_54),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_131),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_116),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_68),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_71),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_56),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_49),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_180),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_60),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_20),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_84),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_70),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_182),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_18),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_113),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_4),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_21),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_99),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_174),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_98),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_97),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_122),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_193),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_189),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_177),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_126),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_39),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_63),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_74),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_18),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_109),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_57),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_78),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_83),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_42),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_102),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_32),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_52),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_19),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_152),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_103),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_133),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_149),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_117),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_5),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_138),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_21),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_62),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_9),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_120),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_101),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_74),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_10),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_41),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_194),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_11),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_26),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_157),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_184),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_16),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_31),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_188),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_80),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_123),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_10),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_173),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_39),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_121),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_59),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_72),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_11),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_175),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_7),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_36),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_185),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_70),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_46),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_144),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_44),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_187),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_33),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_196),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_63),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_171),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_77),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_20),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_41),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_143),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_112),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_72),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_124),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_45),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_169),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_119),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_165),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_48),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_110),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_8),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_6),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_141),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_34),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_23),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_1),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_24),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_89),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_148),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_12),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_191),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_230),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_203),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_215),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_216),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_229),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_224),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_224),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_211),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_270),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_288),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_232),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_291),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_211),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_299),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_233),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_304),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_350),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_234),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_350),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_236),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_214),
.B(n_1),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_224),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_233),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_308),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

BUFx2_ASAP7_75t_SL g422 ( 
.A(n_202),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_237),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_240),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_228),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_242),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_248),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_228),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_247),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_249),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_228),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_251),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_256),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_251),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_251),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_200),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_258),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_259),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_308),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_261),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_263),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_258),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_324),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_258),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_264),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_269),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_262),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_301),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_301),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_277),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_348),
.B(n_2),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_281),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_262),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_235),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_341),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_284),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_207),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_235),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_214),
.B(n_2),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_235),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_341),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_201),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_286),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_201),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_290),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_293),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_205),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_205),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_294),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_218),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_307),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_218),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_311),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_221),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_314),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_221),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_318),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_323),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_204),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_239),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_239),
.B(n_246),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_253),
.B(n_3),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_329),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_346),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_360),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_371),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_207),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_434),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_393),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_422),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_469),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_395),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_469),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_398),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_472),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_413),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_399),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_451),
.A2(n_199),
.B(n_197),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_458),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_463),
.B(n_253),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_400),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_407),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_414),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_416),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_458),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_473),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_458),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_423),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_463),
.B(n_347),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_426),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_396),
.B(n_285),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_415),
.B(n_347),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_405),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_402),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_475),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_475),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_427),
.B(n_248),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_403),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_429),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_477),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_397),
.B(n_248),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_433),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_406),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_403),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_397),
.B(n_332),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_408),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_440),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_479),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_449),
.B(n_332),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_454),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_468),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_470),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_471),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_476),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_412),
.B(n_231),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_481),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_488),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_437),
.B(n_202),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_446),
.A2(n_198),
.B1(n_208),
.B2(n_206),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_489),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_401),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_410),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_490),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_424),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_422),
.B(n_220),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_485),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_401),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_446),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_494),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_511),
.B(n_465),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_533),
.B(n_332),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_547),
.B(n_491),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_498),
.B(n_412),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_430),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_498),
.B(n_404),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_500),
.B(n_409),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_528),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_366),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_533),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_499),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_499),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_502),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_505),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_538),
.A2(n_441),
.B1(n_444),
.B2(n_420),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_526),
.B(n_462),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_538),
.B(n_542),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_532),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_508),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_220),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_518),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_507),
.B(n_462),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_438),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_526),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_568),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_538),
.B(n_255),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_527),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_538),
.B(n_262),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_518),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_511),
.B(n_465),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_527),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_518),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_518),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_527),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_542),
.B(n_255),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_542),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_571),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_542),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_555),
.B(n_486),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_503),
.B(n_492),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_520),
.B(n_459),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_518),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

BUFx10_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_486),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_510),
.B(n_366),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_510),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_532),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_564),
.B(n_274),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_514),
.B(n_492),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_532),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_532),
.B(n_364),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_517),
.A2(n_455),
.B1(n_436),
.B2(n_419),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_540),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_544),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_532),
.B(n_364),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_522),
.B(n_459),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_564),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_442),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_519),
.B(n_443),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_497),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_523),
.B(n_448),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_497),
.Y(n_652)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_559),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_564),
.Y(n_654)
);

OAI21xp33_ASAP7_75t_L g655 ( 
.A1(n_531),
.A2(n_421),
.B(n_460),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_532),
.B(n_366),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_495),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_564),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_565),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_535),
.B(n_456),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_531),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_539),
.B(n_461),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_564),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_545),
.B(n_474),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_570),
.B(n_370),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_559),
.A2(n_213),
.B1(n_313),
.B2(n_300),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_525),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_524),
.B(n_285),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_536),
.B(n_425),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_567),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_506),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_548),
.B(n_549),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_506),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_501),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_570),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_570),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_550),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

CKINVDCx8_ASAP7_75t_R g686 ( 
.A(n_551),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_552),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_553),
.B(n_370),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_557),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_537),
.B(n_419),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_495),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_546),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_546),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_553),
.B(n_370),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_495),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_524),
.B(n_285),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_495),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_554),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_556),
.B(n_436),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_553),
.B(n_210),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_516),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_556),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_516),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_560),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_569),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_572),
.Y(n_710)
);

INVx6_ASAP7_75t_L g711 ( 
.A(n_495),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_572),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_516),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_495),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_504),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_553),
.B(n_331),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_504),
.B(n_197),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_504),
.B(n_274),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_493),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_509),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_493),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_504),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_496),
.B(n_428),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_562),
.B(n_478),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_566),
.B(n_480),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_605),
.A2(n_483),
.B1(n_482),
.B2(n_336),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_691),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_691),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_595),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_595),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_605),
.B(n_504),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_574),
.A2(n_250),
.B1(n_265),
.B2(n_246),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_580),
.B(n_466),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_701),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_623),
.B(n_411),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_574),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_577),
.B(n_504),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_595),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_589),
.A2(n_590),
.B(n_598),
.C(n_575),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_589),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_590),
.A2(n_467),
.B(n_319),
.C(n_292),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_594),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_661),
.B(n_496),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_661),
.B(n_710),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_598),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_608),
.B(n_373),
.Y(n_747)
);

NOR2x2_ASAP7_75t_L g748 ( 
.A(n_621),
.B(n_274),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_618),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_608),
.A2(n_697),
.B1(n_706),
.B2(n_687),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_673),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_L g753 ( 
.A1(n_639),
.A2(n_417),
.B1(n_487),
.B2(n_464),
.C(n_309),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_578),
.B(n_209),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_584),
.B(n_285),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_579),
.A2(n_280),
.B1(n_231),
.B2(n_268),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_620),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_710),
.B(n_199),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_621),
.A2(n_375),
.B1(n_376),
.B2(n_382),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_594),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_SL g762 ( 
.A(n_686),
.B(n_231),
.Y(n_762)
);

AND2x6_ASAP7_75t_SL g763 ( 
.A(n_602),
.B(n_250),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_701),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_584),
.B(n_285),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_723),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_687),
.B(n_219),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_697),
.B(n_219),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_SL g769 ( 
.A1(n_668),
.A2(n_303),
.B1(n_276),
.B2(n_337),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_686),
.B(n_231),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_704),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_704),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_578),
.B(n_358),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_706),
.B(n_222),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_688),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_643),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_707),
.B(n_285),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_688),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_707),
.B(n_222),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_708),
.B(n_225),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_608),
.A2(n_712),
.B1(n_708),
.B2(n_611),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_623),
.B(n_207),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_592),
.B(n_655),
.C(n_643),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_585),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_723),
.Y(n_786)
);

AND2x2_ASAP7_75t_SL g787 ( 
.A(n_670),
.B(n_322),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_586),
.B(n_225),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_709),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_603),
.B(n_359),
.C(n_417),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_670),
.B(n_322),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_621),
.A2(n_384),
.B1(n_389),
.B2(n_390),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_621),
.A2(n_392),
.B1(n_344),
.B2(n_340),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_587),
.B(n_226),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_576),
.A2(n_275),
.B1(n_226),
.B2(n_244),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_673),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_588),
.B(n_244),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_702),
.B(n_322),
.Y(n_798)
);

BUFx8_ASAP7_75t_L g799 ( 
.A(n_681),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_716),
.B(n_354),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_625),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_721),
.B(n_212),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_625),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_630),
.Y(n_804)
);

BUFx8_ASAP7_75t_L g805 ( 
.A(n_681),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_671),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_608),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_606),
.B(n_617),
.Y(n_808)
);

BUFx6f_ASAP7_75t_SL g809 ( 
.A(n_627),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_591),
.B(n_354),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_593),
.B(n_217),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_597),
.B(n_245),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_631),
.B(n_633),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_608),
.A2(n_312),
.B1(n_309),
.B2(n_305),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_676),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_630),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_599),
.A2(n_387),
.B(n_312),
.C(n_265),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_608),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_629),
.A2(n_354),
.B1(n_339),
.B2(n_340),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_245),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_223),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_576),
.B(n_464),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_646),
.B(n_275),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_575),
.A2(n_378),
.B1(n_349),
.B2(n_352),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_593),
.B(n_227),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_287),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_629),
.B(n_238),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_671),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_649),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_684),
.B(n_287),
.Y(n_830)
);

BUFx5_ASAP7_75t_L g831 ( 
.A(n_632),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_693),
.B(n_306),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_694),
.B(n_306),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_700),
.B(n_320),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_611),
.A2(n_378),
.B(n_266),
.C(n_271),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_576),
.B(n_320),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_649),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_647),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_629),
.B(n_241),
.Y(n_839)
);

NAND2x1_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_524),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_583),
.A2(n_273),
.B1(n_296),
.B2(n_282),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_581),
.B(n_207),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_662),
.B(n_325),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_662),
.B(n_325),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_583),
.A2(n_380),
.B1(n_377),
.B2(n_362),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_583),
.B(n_339),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_652),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_573),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_719),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_627),
.B(n_268),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_672),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_656),
.A2(n_509),
.B(n_521),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_664),
.B(n_666),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_652),
.Y(n_854)
);

BUFx5_ASAP7_75t_L g855 ( 
.A(n_632),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_664),
.B(n_344),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_630),
.B(n_345),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_669),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_627),
.B(n_268),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_667),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_669),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_672),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_675),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_628),
.B(n_268),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_628),
.B(n_355),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_666),
.B(n_345),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_619),
.A2(n_601),
.B1(n_635),
.B2(n_622),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_634),
.B(n_524),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_662),
.B(n_607),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_674),
.B(n_243),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_679),
.B(n_357),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_653),
.B(n_252),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_675),
.Y(n_873)
);

AND2x6_ASAP7_75t_SL g874 ( 
.A(n_648),
.B(n_266),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_654),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_678),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_689),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_718),
.A2(n_272),
.B1(n_352),
.B2(n_349),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_607),
.B(n_254),
.Y(n_879)
);

AND2x6_ASAP7_75t_L g880 ( 
.A(n_604),
.B(n_357),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_610),
.A2(n_362),
.B1(n_377),
.B2(n_380),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_678),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_679),
.B(n_563),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_695),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_718),
.A2(n_271),
.B1(n_273),
.B2(n_282),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_682),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_628),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_610),
.B(n_521),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_640),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_612),
.B(n_521),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_654),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_612),
.B(n_563),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_682),
.Y(n_893)
);

AND2x6_ASAP7_75t_SL g894 ( 
.A(n_663),
.B(n_272),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_613),
.B(n_260),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_573),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_613),
.B(n_563),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_736),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_SL g899 ( 
.A(n_769),
.B(n_753),
.C(n_872),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_755),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_807),
.Y(n_901)
);

AND2x2_ASAP7_75t_SL g902 ( 
.A(n_732),
.B(n_665),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_733),
.B(n_616),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_752),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_775),
.Y(n_906)
);

NOR2x1_ASAP7_75t_R g907 ( 
.A(n_778),
.B(n_582),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_807),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_730),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_735),
.B(n_724),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_807),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_755),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_889),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_R g914 ( 
.A(n_848),
.B(n_582),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_796),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_766),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_818),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_SL g919 ( 
.A1(n_838),
.A2(n_690),
.B1(n_659),
.B2(n_641),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_730),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_736),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_766),
.Y(n_922)
);

AND3x1_ASAP7_75t_SL g923 ( 
.A(n_763),
.B(n_305),
.C(n_296),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_R g924 ( 
.A(n_887),
.B(n_641),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_815),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_650),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_818),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_733),
.B(n_616),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_741),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_858),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_786),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_818),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_896),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_872),
.B(n_660),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_818),
.Y(n_935)
);

BUFx8_ASAP7_75t_L g936 ( 
.A(n_809),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_804),
.B(n_725),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_746),
.B(n_626),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_782),
.B(n_662),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_729),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_727),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_738),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_741),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_849),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_728),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_734),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_743),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_887),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_776),
.B(n_659),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_SL g950 ( 
.A1(n_851),
.A2(n_690),
.B1(n_279),
.B2(n_372),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_764),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_801),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_SL g953 ( 
.A(n_821),
.B(n_278),
.C(n_267),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_732),
.A2(n_824),
.B1(n_787),
.B2(n_791),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_743),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_801),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_816),
.B(n_722),
.Y(n_957)
);

AO22x1_ASAP7_75t_L g958 ( 
.A1(n_870),
.A2(n_328),
.B1(n_310),
.B2(n_302),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_840),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_803),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_803),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_740),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_829),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_829),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_745),
.B(n_626),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_811),
.B(n_283),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_837),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_782),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_SL g969 ( 
.A(n_821),
.B(n_295),
.C(n_289),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_837),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_877),
.B(n_645),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_771),
.B(n_722),
.Y(n_972)
);

INVx3_ASAP7_75t_SL g973 ( 
.A(n_748),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_809),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_822),
.Y(n_975)
);

OR2x6_ASAP7_75t_SL g976 ( 
.A(n_819),
.B(n_297),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_749),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_847),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_761),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_754),
.B(n_645),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_750),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_875),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_884),
.B(n_806),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_862),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_799),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_824),
.A2(n_391),
.B1(n_387),
.B2(n_334),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_822),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_857),
.B(n_717),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_799),
.B(n_298),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_805),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_758),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_828),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_827),
.B(n_316),
.C(n_315),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_857),
.B(n_717),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_875),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_808),
.A2(n_680),
.B1(n_685),
.B2(n_683),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_808),
.A2(n_680),
.B1(n_685),
.B2(n_683),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_785),
.B(n_860),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_SL g999 ( 
.A(n_827),
.B(n_321),
.C(n_317),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_847),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_805),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_813),
.B(n_658),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_854),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_787),
.A2(n_391),
.B1(n_388),
.B2(n_334),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_772),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_781),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_857),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_744),
.B(n_658),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_789),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_751),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_731),
.B(n_677),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_754),
.B(n_355),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_802),
.B(n_677),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_863),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_873),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_873),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_783),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_839),
.B(n_327),
.C(n_326),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_751),
.B(n_662),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_861),
.Y(n_1022)
);

OAI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_793),
.A2(n_487),
.B1(n_717),
.B2(n_374),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_784),
.B(n_714),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_802),
.B(n_692),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_861),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_876),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_850),
.B(n_654),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_853),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_882),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_882),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_773),
.A2(n_870),
.B1(n_846),
.B2(n_836),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_773),
.B(n_714),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_886),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_886),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_SL g1036 ( 
.A(n_859),
.B(n_654),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_893),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_879),
.B(n_692),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_893),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_864),
.Y(n_1040)
);

OR2x2_ASAP7_75t_SL g1041 ( 
.A(n_825),
.B(n_367),
.Y(n_1041)
);

BUFx4f_ASAP7_75t_L g1042 ( 
.A(n_865),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_888),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_842),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_726),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_879),
.B(n_692),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_895),
.B(n_696),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_890),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_739),
.A2(n_388),
.B(n_385),
.C(n_374),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_839),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_739),
.A2(n_715),
.B1(n_604),
.B2(n_614),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_788),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_790),
.B(n_355),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_867),
.B(n_330),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_895),
.B(n_696),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_760),
.A2(n_715),
.B1(n_696),
.B2(n_711),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_892),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_762),
.B(n_355),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_874),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_792),
.A2(n_711),
.B1(n_615),
.B2(n_609),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_835),
.B(n_654),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_759),
.B(n_609),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_897),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_880),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_770),
.B(n_657),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_894),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_R g1067 ( 
.A(n_737),
.B(n_333),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_830),
.B(n_614),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_791),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_830),
.B(n_624),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_856),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_747),
.B(n_335),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_757),
.B(n_338),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_866),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_871),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_742),
.B(n_711),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_841),
.A2(n_385),
.B(n_367),
.C(n_431),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_767),
.B(n_609),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_768),
.B(n_615),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_798),
.A2(n_615),
.B1(n_624),
.B2(n_634),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_832),
.B(n_657),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_832),
.B(n_657),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_883),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_869),
.B(n_699),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_774),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_779),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_780),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_841),
.A2(n_379),
.B(n_342),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_794),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_817),
.B(n_386),
.C(n_343),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_954),
.A2(n_814),
.B(n_795),
.C(n_845),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1051),
.A2(n_852),
.B(n_765),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_939),
.A2(n_891),
.B(n_869),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1024),
.A2(n_756),
.B(n_765),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_939),
.A2(n_636),
.B(n_814),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_980),
.B(n_797),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1038),
.A2(n_756),
.B(n_800),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1024),
.A2(n_800),
.B(n_798),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_921),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_917),
.B(n_812),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1064),
.A2(n_810),
.B(n_823),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_904),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_934),
.B(n_820),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_1049),
.A2(n_777),
.B(n_810),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1049),
.A2(n_834),
.A3(n_833),
.B(n_826),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_967),
.B(n_964),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_914),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_934),
.B(n_881),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_980),
.B(n_878),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1064),
.A2(n_777),
.B(n_843),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_SL g1111 ( 
.A1(n_968),
.A2(n_699),
.B(n_600),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_910),
.B(n_843),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_998),
.B(n_878),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_984),
.B(n_885),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_SL g1115 ( 
.A1(n_1024),
.A2(n_1025),
.B(n_1046),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1014),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_1033),
.A2(n_637),
.A3(n_642),
.B(n_703),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1021),
.A2(n_844),
.B(n_868),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_921),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1033),
.B(n_885),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_898),
.A2(n_636),
.B(n_596),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1047),
.A2(n_596),
.B(n_638),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1064),
.A2(n_844),
.B(n_703),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_929),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1012),
.A2(n_705),
.B(n_713),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_929),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1084),
.A2(n_705),
.B(n_713),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_906),
.B(n_85),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1055),
.A2(n_596),
.B(n_638),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_943),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1087),
.B(n_880),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1045),
.A2(n_356),
.B1(n_353),
.B2(n_383),
.C(n_361),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1011),
.A2(n_928),
.B(n_903),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_SL g1134 ( 
.A1(n_954),
.A2(n_720),
.B(n_452),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1083),
.A2(n_453),
.A3(n_431),
.B(n_432),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1013),
.B(n_365),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_918),
.A2(n_720),
.B(n_453),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1089),
.B(n_880),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1085),
.B(n_880),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_906),
.B(n_87),
.Y(n_1140)
);

AOI221x1_ASAP7_75t_L g1141 ( 
.A1(n_1028),
.A2(n_445),
.B1(n_428),
.B2(n_452),
.C(n_432),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_943),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_902),
.A2(n_699),
.B1(n_600),
.B2(n_381),
.Y(n_1143)
);

NAND2x1_ASAP7_75t_L g1144 ( 
.A(n_982),
.B(n_699),
.Y(n_1144)
);

INVxp67_ASAP7_75t_SL g1145 ( 
.A(n_995),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_902),
.B(n_880),
.Y(n_1146)
);

BUFx4_ASAP7_75t_SL g1147 ( 
.A(n_913),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_915),
.B(n_435),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1042),
.B(n_855),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1002),
.A2(n_600),
.B(n_699),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1043),
.A2(n_698),
.B(n_718),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_983),
.B(n_831),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1073),
.A2(n_368),
.B1(n_369),
.B2(n_435),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1086),
.B(n_831),
.Y(n_1154)
);

OAI22x1_ASAP7_75t_L g1155 ( 
.A1(n_1058),
.A2(n_439),
.B1(n_445),
.B2(n_447),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_908),
.B(n_927),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_901),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_944),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_900),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_963),
.A2(n_541),
.B(n_529),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_952),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_917),
.B(n_913),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_1050),
.B(n_90),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_941),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1048),
.A2(n_698),
.B(n_718),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_952),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1084),
.A2(n_439),
.B(n_447),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_988),
.A2(n_600),
.B(n_831),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1078),
.A2(n_450),
.B(n_543),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_901),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_912),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_899),
.A2(n_450),
.B(n_543),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1086),
.B(n_831),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1067),
.A2(n_1054),
.B(n_1019),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_988),
.A2(n_600),
.B(n_855),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1005),
.A2(n_543),
.B1(n_541),
.B2(n_534),
.C(n_529),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_925),
.B(n_529),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1057),
.B(n_831),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_946),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1079),
.A2(n_541),
.B(n_534),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1063),
.A2(n_718),
.B(n_634),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1083),
.A2(n_534),
.A3(n_634),
.B(n_718),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_916),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_996),
.A2(n_509),
.B(n_831),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_933),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_997),
.A2(n_509),
.B(n_855),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_922),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_963),
.A2(n_855),
.B(n_634),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_948),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1042),
.B(n_280),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_964),
.A2(n_855),
.B(n_634),
.Y(n_1191)
);

AO21x1_ASAP7_75t_L g1192 ( 
.A1(n_1028),
.A2(n_280),
.B(n_8),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_918),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_964),
.A2(n_855),
.B(n_139),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1071),
.B(n_524),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_945),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_988),
.A2(n_524),
.B(n_137),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_995),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_967),
.A2(n_142),
.B(n_93),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1074),
.B(n_524),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_3),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_967),
.A2(n_136),
.B(n_183),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_931),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1003),
.A2(n_135),
.B(n_176),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_992),
.B(n_12),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_988),
.A2(n_130),
.B(n_168),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1005),
.B(n_13),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_994),
.A2(n_115),
.B(n_167),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_994),
.A2(n_114),
.B(n_164),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_994),
.A2(n_107),
.B(n_159),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1003),
.A2(n_106),
.B(n_158),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_940),
.B(n_942),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1008),
.B(n_14),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1008),
.B(n_14),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1003),
.A2(n_1030),
.B(n_1004),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_994),
.A2(n_151),
.B(n_147),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_971),
.A2(n_280),
.B(n_105),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_965),
.B(n_17),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1062),
.A2(n_104),
.B(n_91),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_918),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1004),
.A2(n_28),
.B(n_29),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1068),
.A2(n_29),
.B(n_30),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_956),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_951),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_948),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_995),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_930),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1004),
.A2(n_30),
.B(n_32),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_935),
.A2(n_982),
.B(n_1056),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1030),
.A2(n_33),
.B(n_35),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_966),
.B(n_35),
.Y(n_1231)
);

AND2x2_ASAP7_75t_SL g1232 ( 
.A(n_1065),
.B(n_40),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1030),
.A2(n_40),
.B(n_42),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_901),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1015),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_982),
.A2(n_938),
.B(n_995),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_956),
.A2(n_43),
.B(n_44),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_962),
.B(n_43),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1077),
.A2(n_46),
.A3(n_47),
.B(n_48),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_977),
.B(n_50),
.Y(n_1240)
);

AOI211x1_ASAP7_75t_L g1241 ( 
.A1(n_1088),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_960),
.A2(n_1035),
.B(n_1027),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1009),
.A2(n_53),
.B(n_57),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_960),
.A2(n_53),
.B(n_60),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_935),
.A2(n_932),
.B1(n_927),
.B2(n_908),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_961),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1077),
.A2(n_62),
.A3(n_65),
.B(n_66),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_909),
.A2(n_66),
.B(n_67),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_981),
.B(n_67),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_908),
.B(n_68),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1016),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_961),
.A2(n_69),
.A3(n_73),
.B(n_75),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_991),
.B(n_69),
.Y(n_1253)
);

CKINVDCx16_ASAP7_75t_R g1254 ( 
.A(n_914),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1091),
.A2(n_1023),
.B(n_1018),
.C(n_1034),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1164),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1158),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1212),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1189),
.B(n_975),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_1065),
.B1(n_926),
.B2(n_937),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1091),
.A2(n_1037),
.B(n_1010),
.C(n_1060),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1097),
.A2(n_1146),
.B(n_1150),
.Y(n_1262)
);

NAND2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1198),
.B(n_908),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1111),
.B(n_1229),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1103),
.B(n_1040),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1108),
.A2(n_1068),
.B(n_1070),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1103),
.B(n_1040),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1164),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1096),
.B(n_1044),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1232),
.A2(n_973),
.B1(n_926),
.B2(n_1053),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1189),
.B(n_975),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1099),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1196),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1115),
.A2(n_1017),
.B(n_1039),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1133),
.A2(n_1068),
.B(n_1070),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1217),
.A2(n_1072),
.B(n_1080),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1180),
.A2(n_970),
.B(n_1035),
.Y(n_1277)
);

AOI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1136),
.A2(n_1067),
.B(n_949),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1116),
.A2(n_1072),
.B(n_1082),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1115),
.A2(n_1194),
.B(n_1125),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1125),
.A2(n_1027),
.B(n_978),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1236),
.A2(n_1036),
.B(n_920),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1225),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1180),
.A2(n_978),
.B(n_1000),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1169),
.A2(n_1031),
.B(n_1000),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1198),
.B(n_1106),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1099),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1235),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1251),
.Y(n_1289)
);

INVx8_ASAP7_75t_L g1290 ( 
.A(n_1198),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1185),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1112),
.B(n_1007),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1112),
.B(n_1007),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1119),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1162),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1113),
.B(n_987),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_1082),
.B(n_1081),
.Y(n_1298)
);

AO21x2_ASAP7_75t_L g1299 ( 
.A1(n_1134),
.A2(n_1082),
.B(n_1081),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1242),
.A2(n_1039),
.B(n_1031),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1109),
.A2(n_926),
.B1(n_937),
.B2(n_976),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1161),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1242),
.A2(n_970),
.B(n_1017),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1120),
.A2(n_1070),
.B(n_1081),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1166),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1124),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1126),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1184),
.A2(n_920),
.B(n_909),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1130),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1102),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1232),
.B(n_972),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1193),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1098),
.A2(n_1020),
.B(n_999),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1142),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1166),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1222),
.A2(n_986),
.B(n_1036),
.C(n_993),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1184),
.A2(n_920),
.B(n_909),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1159),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1095),
.A2(n_972),
.B(n_1076),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1207),
.A2(n_973),
.B1(n_926),
.B2(n_937),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1223),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1157),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1225),
.B(n_987),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1198),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1223),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1246),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1224),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1174),
.A2(n_937),
.B1(n_1006),
.B2(n_979),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1246),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1179),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1171),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1183),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1193),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1135),
.Y(n_1334)
);

BUFx2_ASAP7_75t_R g1335 ( 
.A(n_1149),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1094),
.A2(n_986),
.B(n_969),
.C(n_953),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1139),
.A2(n_976),
.B(n_1069),
.C(n_1090),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1187),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1203),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_1029),
.B(n_1061),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1177),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1092),
.A2(n_972),
.B(n_957),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1201),
.B(n_1029),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1135),
.Y(n_1344)
);

CKINVDCx6p67_ASAP7_75t_R g1345 ( 
.A(n_1254),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1192),
.A2(n_1208),
.B(n_1206),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1135),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1172),
.A2(n_1205),
.B(n_1218),
.C(n_1163),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1114),
.B(n_1029),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1141),
.A2(n_1143),
.A3(n_1155),
.B(n_1093),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1153),
.A2(n_935),
.A3(n_1061),
.B(n_1069),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1135),
.Y(n_1352)
);

CKINVDCx6p67_ASAP7_75t_R g1353 ( 
.A(n_1162),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1186),
.A2(n_1076),
.B(n_1061),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1215),
.A2(n_1029),
.B(n_1061),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1127),
.A2(n_1076),
.B(n_927),
.Y(n_1356)
);

AOI21xp33_ASAP7_75t_L g1357 ( 
.A1(n_1107),
.A2(n_919),
.B(n_907),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1107),
.B(n_950),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1162),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1226),
.B(n_957),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1138),
.B(n_958),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1190),
.B(n_957),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1127),
.A2(n_1076),
.B(n_927),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1160),
.A2(n_932),
.B(n_1069),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1227),
.A2(n_1066),
.B1(n_1059),
.B2(n_1140),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1157),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1148),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1092),
.A2(n_932),
.B(n_979),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1238),
.B(n_979),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1188),
.A2(n_932),
.B(n_979),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1100),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1157),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1179),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1188),
.A2(n_955),
.B(n_947),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1176),
.A2(n_1244),
.B(n_1233),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1191),
.A2(n_955),
.B(n_947),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1167),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1100),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1231),
.A2(n_1132),
.B1(n_1131),
.B2(n_1213),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1240),
.B(n_1041),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1118),
.A2(n_911),
.B(n_905),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1105),
.B(n_955),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_SL g1383 ( 
.A1(n_1220),
.A2(n_923),
.B(n_947),
.C(n_955),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1191),
.A2(n_947),
.B(n_911),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1123),
.A2(n_911),
.B(n_901),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1100),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1105),
.B(n_911),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1214),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1249),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1152),
.A2(n_974),
.B(n_1059),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1105),
.B(n_905),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1123),
.A2(n_905),
.B(n_959),
.Y(n_1392)
);

INVx8_ASAP7_75t_L g1393 ( 
.A(n_1157),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1170),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1226),
.B(n_905),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1167),
.A2(n_959),
.B(n_924),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1244),
.A2(n_974),
.B(n_959),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1147),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1137),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1204),
.A2(n_959),
.B(n_924),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1145),
.B(n_1001),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1145),
.A2(n_985),
.B1(n_1026),
.B2(n_1022),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1149),
.B(n_1052),
.Y(n_1404)
);

AO21x1_ASAP7_75t_L g1405 ( 
.A1(n_1221),
.A2(n_75),
.B(n_76),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1248),
.A2(n_990),
.B(n_1001),
.C(n_1022),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1221),
.A2(n_1233),
.B(n_1228),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1237),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1228),
.A2(n_1052),
.B(n_78),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1211),
.A2(n_936),
.B(n_990),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1178),
.B(n_985),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1151),
.A2(n_936),
.B(n_989),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1110),
.A2(n_936),
.B(n_989),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1170),
.B(n_1234),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1209),
.A2(n_1210),
.B(n_1216),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1154),
.B(n_1173),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1250),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1110),
.A2(n_1202),
.B(n_1199),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1147),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1156),
.A2(n_1168),
.B1(n_1175),
.B2(n_1245),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1128),
.A2(n_1250),
.B1(n_1200),
.B2(n_1195),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1241),
.B(n_1144),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1165),
.A2(n_1104),
.B1(n_1181),
.B2(n_1234),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1252),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1199),
.B(n_1202),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1170),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1273),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1272),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1270),
.A2(n_1380),
.B(n_1278),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1402),
.B(n_1234),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1282),
.A2(n_1156),
.B(n_1129),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1320),
.A2(n_1234),
.B1(n_1170),
.B2(n_1104),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1402),
.B(n_1182),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1290),
.B(n_1230),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1328),
.A2(n_1104),
.B1(n_1197),
.B2(n_1121),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1257),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1272),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1260),
.A2(n_1122),
.B1(n_1105),
.B2(n_1239),
.C(n_1247),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1283),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1301),
.A2(n_1389),
.B1(n_1399),
.B2(n_1388),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1288),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1266),
.A2(n_1243),
.B1(n_1230),
.B2(n_1101),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1311),
.B(n_1367),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1287),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1265),
.A2(n_1243),
.B1(n_1219),
.B2(n_1101),
.Y(n_1445)
);

OAI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1379),
.A2(n_1243),
.B(n_1239),
.C(n_1247),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_R g1447 ( 
.A1(n_1403),
.A2(n_1239),
.B(n_1247),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_1182),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1289),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1312),
.B(n_1182),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1318),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1341),
.B(n_1239),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1258),
.B(n_1269),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1331),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1267),
.B(n_1252),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1276),
.A2(n_1252),
.B1(n_1117),
.B2(n_1182),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1273),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1332),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1292),
.B(n_1117),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1349),
.B(n_1117),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1276),
.A2(n_1117),
.B1(n_1252),
.B2(n_1293),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1297),
.A2(n_1365),
.B1(n_1362),
.B2(n_1353),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1346),
.A2(n_1280),
.B(n_1408),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1276),
.A2(n_1319),
.B(n_1279),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1313),
.A2(n_1358),
.B1(n_1304),
.B2(n_1404),
.Y(n_1465)
);

CKINVDCx16_ASAP7_75t_R g1466 ( 
.A(n_1359),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1313),
.A2(n_1279),
.B1(n_1295),
.B2(n_1405),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1256),
.B(n_1268),
.Y(n_1468)
);

OAI222xp33_ASAP7_75t_L g1469 ( 
.A1(n_1422),
.A2(n_1343),
.B1(n_1361),
.B2(n_1369),
.C1(n_1338),
.C2(n_1339),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1291),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1411),
.B(n_1330),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1391),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1330),
.B(n_1373),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1313),
.A2(n_1279),
.B1(n_1295),
.B2(n_1405),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1373),
.B(n_1259),
.Y(n_1475)
);

AOI221xp5_ASAP7_75t_L g1476 ( 
.A1(n_1316),
.A2(n_1336),
.B1(n_1255),
.B2(n_1348),
.C(n_1261),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1327),
.Y(n_1477)
);

OR2x6_ASAP7_75t_L g1478 ( 
.A(n_1290),
.B(n_1264),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1310),
.B(n_1390),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1391),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1316),
.A2(n_1336),
.B1(n_1255),
.B2(n_1348),
.C(n_1261),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1353),
.A2(n_1359),
.B1(n_1345),
.B2(n_1422),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1287),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1264),
.A2(n_1275),
.B(n_1415),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1294),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1371),
.A2(n_1345),
.B1(n_1412),
.B2(n_1357),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1424),
.A2(n_1347),
.A3(n_1334),
.B(n_1352),
.Y(n_1487)
);

AO31x2_ASAP7_75t_L g1488 ( 
.A1(n_1334),
.A2(n_1347),
.A3(n_1352),
.B(n_1344),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1306),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1371),
.A2(n_1409),
.B1(n_1422),
.B2(n_1386),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1378),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1493)
);

OAI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1406),
.A2(n_1378),
.B(n_1337),
.C(n_1383),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1314),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1290),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1335),
.A2(n_1423),
.B1(n_1406),
.B2(n_1417),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1283),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1264),
.A2(n_1259),
.B1(n_1271),
.B2(n_1323),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1296),
.Y(n_1500)
);

OAI211xp5_ASAP7_75t_L g1501 ( 
.A1(n_1337),
.A2(n_1383),
.B(n_1409),
.C(n_1419),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1271),
.B(n_1323),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1264),
.A2(n_1323),
.B1(n_1324),
.B2(n_1422),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1409),
.A2(n_1386),
.B1(n_1290),
.B2(n_1324),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1296),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1382),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1366),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1421),
.A2(n_1398),
.B1(n_1416),
.B2(n_1400),
.C(n_1420),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1302),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1324),
.A2(n_1360),
.B1(n_1387),
.B2(n_1382),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1305),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1315),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1413),
.B(n_1324),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1360),
.A2(n_1387),
.B1(n_1312),
.B2(n_1333),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1280),
.A2(n_1356),
.B(n_1363),
.Y(n_1516)
);

OAI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1416),
.A2(n_1262),
.B1(n_1425),
.B2(n_1354),
.C(n_1312),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1386),
.A2(n_1299),
.B1(n_1315),
.B2(n_1325),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1360),
.A2(n_1333),
.B1(n_1263),
.B2(n_1395),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1381),
.A2(n_1397),
.B1(n_1299),
.B2(n_1396),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1321),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1356),
.A2(n_1363),
.B(n_1285),
.Y(n_1522)
);

CKINVDCx8_ASAP7_75t_R g1523 ( 
.A(n_1393),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1366),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1321),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1333),
.A2(n_1263),
.B1(n_1395),
.B2(n_1329),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1351),
.B(n_1414),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1342),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1325),
.A2(n_1329),
.B1(n_1326),
.B2(n_1372),
.Y(n_1529)
);

OAI211xp5_ASAP7_75t_L g1530 ( 
.A1(n_1413),
.A2(n_1397),
.B(n_1407),
.C(n_1326),
.Y(n_1530)
);

CKINVDCx11_ASAP7_75t_R g1531 ( 
.A(n_1393),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1299),
.A2(n_1342),
.B1(n_1381),
.B2(n_1397),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1274),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1372),
.B(n_1322),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1351),
.B(n_1395),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1396),
.A2(n_1401),
.B1(n_1407),
.B2(n_1342),
.Y(n_1536)
);

NOR3xp33_ASAP7_75t_SL g1537 ( 
.A(n_1351),
.B(n_1410),
.C(n_1393),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1263),
.A2(n_1286),
.B1(n_1394),
.B2(n_1426),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1375),
.A2(n_1298),
.B1(n_1407),
.B2(n_1274),
.Y(n_1539)
);

INVxp33_ASAP7_75t_SL g1540 ( 
.A(n_1410),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1351),
.B(n_1414),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1351),
.B(n_1414),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1394),
.B(n_1426),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1322),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1375),
.A2(n_1298),
.B1(n_1340),
.B2(n_1277),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1372),
.A2(n_1286),
.B1(n_1322),
.B2(n_1393),
.Y(n_1546)
);

AO21x2_ASAP7_75t_L g1547 ( 
.A1(n_1418),
.A2(n_1377),
.B(n_1298),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1401),
.A2(n_1375),
.B1(n_1355),
.B2(n_1425),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1322),
.B(n_1350),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1300),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1322),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1286),
.A2(n_1425),
.B1(n_1377),
.B2(n_1277),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1300),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1303),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1303),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1355),
.A2(n_1340),
.B1(n_1368),
.B2(n_1364),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1277),
.A2(n_1350),
.B1(n_1368),
.B2(n_1392),
.Y(n_1557)
);

BUFx8_ASAP7_75t_L g1558 ( 
.A(n_1350),
.Y(n_1558)
);

BUFx8_ASAP7_75t_L g1559 ( 
.A(n_1350),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1364),
.B(n_1317),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1285),
.A2(n_1281),
.B1(n_1284),
.B2(n_1308),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1350),
.A2(n_1392),
.B1(n_1385),
.B2(n_1308),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1374),
.A2(n_1376),
.B1(n_1317),
.B2(n_1370),
.Y(n_1563)
);

AOI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1418),
.A2(n_1284),
.B(n_1281),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1565)
);

NOR3xp33_ASAP7_75t_SL g1566 ( 
.A(n_1384),
.B(n_1385),
.C(n_1370),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1384),
.A2(n_934),
.B1(n_1108),
.B2(n_872),
.C(n_769),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1260),
.A2(n_1232),
.B1(n_902),
.B2(n_668),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1345),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1270),
.A2(n_1108),
.B1(n_902),
.B2(n_934),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1282),
.A2(n_1111),
.B(n_1133),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1380),
.A2(n_934),
.B(n_757),
.C(n_899),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1260),
.A2(n_1232),
.B1(n_902),
.B2(n_668),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1380),
.A2(n_934),
.B1(n_579),
.B2(n_567),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1260),
.B(n_1232),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1291),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1282),
.A2(n_1111),
.B(n_1133),
.Y(n_1577)
);

BUFx12f_ASAP7_75t_L g1578 ( 
.A(n_1295),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1270),
.A2(n_1108),
.B1(n_902),
.B2(n_934),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1257),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1270),
.A2(n_1108),
.B1(n_902),
.B2(n_934),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1283),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_R g1583 ( 
.A(n_1290),
.B(n_906),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1272),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1269),
.B(n_1349),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1272),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1380),
.A2(n_1232),
.B1(n_902),
.B2(n_1108),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1272),
.Y(n_1588)
);

INVx4_ASAP7_75t_L g1589 ( 
.A(n_1290),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1380),
.A2(n_934),
.B1(n_579),
.B2(n_567),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1257),
.Y(n_1591)
);

NOR3xp33_ASAP7_75t_SL g1592 ( 
.A(n_1412),
.B(n_1059),
.C(n_1301),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1272),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1345),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_L g1595 ( 
.A(n_1453),
.B(n_1501),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1496),
.Y(n_1596)
);

AOI222xp33_ASAP7_75t_L g1597 ( 
.A1(n_1570),
.A2(n_1581),
.B1(n_1579),
.B2(n_1587),
.C1(n_1575),
.C2(n_1572),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1575),
.B2(n_1587),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1468),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1436),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1465),
.B2(n_1567),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1439),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1574),
.A2(n_1590),
.B1(n_1429),
.B2(n_1462),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1476),
.A2(n_1481),
.B1(n_1465),
.B2(n_1440),
.C(n_1462),
.Y(n_1604)
);

AOI222xp33_ASAP7_75t_L g1605 ( 
.A1(n_1497),
.A2(n_1440),
.B1(n_1443),
.B2(n_1479),
.C1(n_1471),
.C2(n_1477),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1506),
.B(n_1527),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1494),
.A2(n_1583),
.B1(n_1503),
.B2(n_1578),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1542),
.B(n_1455),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1508),
.A2(n_1486),
.B1(n_1482),
.B2(n_1491),
.Y(n_1609)
);

AOI222xp33_ASAP7_75t_L g1610 ( 
.A1(n_1470),
.A2(n_1576),
.B1(n_1473),
.B2(n_1467),
.C1(n_1474),
.C2(n_1427),
.Y(n_1610)
);

OAI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1467),
.A2(n_1474),
.B(n_1446),
.C(n_1490),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1571),
.A2(n_1577),
.B(n_1464),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1484),
.A2(n_1431),
.B(n_1529),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1439),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1457),
.Y(n_1615)
);

A2O1A1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1592),
.A2(n_1490),
.B(n_1438),
.C(n_1504),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1482),
.A2(n_1493),
.B1(n_1475),
.B2(n_1585),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1583),
.A2(n_1559),
.B1(n_1558),
.B2(n_1466),
.Y(n_1618)
);

OAI33xp33_ASAP7_75t_L g1619 ( 
.A1(n_1441),
.A2(n_1449),
.A3(n_1591),
.B1(n_1451),
.B2(n_1580),
.B3(n_1458),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1569),
.A2(n_1594),
.B1(n_1502),
.B2(n_1592),
.Y(n_1620)
);

OAI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1504),
.A2(n_1461),
.B(n_1459),
.C(n_1442),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1499),
.A2(n_1452),
.B1(n_1559),
.B2(n_1558),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1529),
.A2(n_1478),
.B(n_1435),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1433),
.A2(n_1448),
.B1(n_1511),
.B2(n_1459),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1478),
.B(n_1433),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1539),
.A2(n_1561),
.B(n_1545),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1515),
.A2(n_1460),
.B1(n_1432),
.B2(n_1478),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1535),
.A2(n_1430),
.B1(n_1582),
.B2(n_1498),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1582),
.A2(n_1447),
.B1(n_1518),
.B2(n_1454),
.Y(n_1629)
);

AOI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1445),
.A2(n_1434),
.B(n_1552),
.Y(n_1630)
);

BUFx12f_ASAP7_75t_L g1631 ( 
.A(n_1531),
.Y(n_1631)
);

AOI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1461),
.A2(n_1517),
.B(n_1442),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1469),
.A2(n_1518),
.B1(n_1489),
.B2(n_1495),
.C(n_1485),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1430),
.A2(n_1540),
.B1(n_1541),
.B2(n_1549),
.Y(n_1634)
);

AOI222xp33_ASAP7_75t_L g1635 ( 
.A1(n_1469),
.A2(n_1512),
.B1(n_1510),
.B2(n_1505),
.C1(n_1513),
.C2(n_1519),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1492),
.A2(n_1523),
.B1(n_1589),
.B2(n_1496),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1507),
.A2(n_1524),
.B1(n_1531),
.B2(n_1526),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1530),
.A2(n_1563),
.B(n_1562),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1520),
.A2(n_1514),
.B1(n_1551),
.B2(n_1544),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1520),
.A2(n_1532),
.B1(n_1589),
.B2(n_1456),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1487),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1543),
.B(n_1428),
.Y(n_1642)
);

A2O1A1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1532),
.A2(n_1537),
.B(n_1456),
.C(n_1545),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1437),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1514),
.A2(n_1434),
.B1(n_1546),
.B2(n_1556),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1557),
.A2(n_1546),
.B1(n_1528),
.B2(n_1539),
.C(n_1538),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1537),
.A2(n_1536),
.B(n_1566),
.C(n_1548),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1509),
.A2(n_1593),
.B1(n_1444),
.B2(n_1584),
.C1(n_1588),
.C2(n_1483),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1488),
.B(n_1487),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1434),
.A2(n_1586),
.B1(n_1525),
.B2(n_1521),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1500),
.B(n_1450),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1488),
.B(n_1463),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1553),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1534),
.A2(n_1450),
.B1(n_1548),
.B2(n_1536),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1561),
.A2(n_1533),
.B1(n_1560),
.B2(n_1566),
.C(n_1554),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1555),
.A2(n_1550),
.B1(n_1463),
.B2(n_1565),
.C(n_1547),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1565),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1547),
.B(n_1560),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1522),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1560),
.A2(n_1587),
.B1(n_1568),
.B2(n_1573),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1472),
.B(n_1480),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1585),
.B(n_1453),
.Y(n_1666)
);

OAI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1572),
.A2(n_757),
.B(n_1573),
.C(n_1568),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1572),
.A2(n_757),
.B(n_1573),
.C(n_1568),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1468),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1472),
.B(n_1480),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1574),
.A2(n_934),
.B(n_579),
.Y(n_1673)
);

OAI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1572),
.A2(n_757),
.B(n_1573),
.C(n_1568),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1570),
.A2(n_1579),
.B1(n_1581),
.B2(n_1587),
.C1(n_1232),
.C2(n_934),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1585),
.B(n_1453),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1468),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1472),
.Y(n_1679)
);

AOI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1570),
.A2(n_934),
.B(n_1579),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1684)
);

BUFx12f_ASAP7_75t_L g1685 ( 
.A(n_1569),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1570),
.A2(n_1581),
.B1(n_1579),
.B2(n_934),
.C(n_1587),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1585),
.B(n_1453),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1464),
.A2(n_1438),
.B(n_1539),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1570),
.A2(n_1581),
.B1(n_1579),
.B2(n_934),
.C(n_1587),
.Y(n_1691)
);

OAI211xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1572),
.A2(n_1278),
.B(n_899),
.C(n_1574),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1567),
.A2(n_769),
.B1(n_1587),
.B2(n_1579),
.C(n_1581),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1695)
);

BUFx10_ASAP7_75t_L g1696 ( 
.A(n_1594),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1571),
.A2(n_1577),
.B(n_1111),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1496),
.B(n_1198),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1478),
.B(n_1433),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1585),
.B(n_1453),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1436),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1574),
.A2(n_1590),
.B1(n_934),
.B2(n_1587),
.C(n_1572),
.Y(n_1705)
);

OAI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1574),
.A2(n_934),
.B1(n_579),
.B2(n_1590),
.C(n_1573),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1570),
.A2(n_934),
.B(n_1579),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1564),
.A2(n_1280),
.B(n_1516),
.Y(n_1710)
);

INVxp67_ASAP7_75t_R g1711 ( 
.A(n_1471),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1568),
.A2(n_1573),
.B1(n_1579),
.B2(n_1570),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1587),
.A2(n_1568),
.B1(n_1573),
.B2(n_1574),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_SL g1718 ( 
.A(n_1498),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1433),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1531),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1654),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1608),
.B(n_1644),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1608),
.B(n_1644),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1663),
.B(n_1672),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1650),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1659),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1641),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1606),
.B(n_1653),
.Y(n_1728)
);

INVx5_ASAP7_75t_SL g1729 ( 
.A(n_1638),
.Y(n_1729)
);

BUFx8_ASAP7_75t_L g1730 ( 
.A(n_1718),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1658),
.B(n_1621),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1600),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1660),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1689),
.B(n_1626),
.Y(n_1734)
);

CKINVDCx16_ASAP7_75t_R g1735 ( 
.A(n_1631),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1706),
.B(n_1673),
.C(n_1674),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1626),
.B(n_1643),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1679),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1643),
.B(n_1648),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1601),
.A2(n_1598),
.B1(n_1695),
.B2(n_1694),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1648),
.B(n_1638),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1638),
.B(n_1612),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1660),
.B(n_1625),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1657),
.B(n_1630),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1666),
.B(n_1676),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1688),
.B(n_1702),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1662),
.B(n_1678),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1710),
.A2(n_1613),
.B(n_1697),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1683),
.A2(n_1714),
.B(n_1717),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1647),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1632),
.A2(n_1707),
.B(n_1680),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1646),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1599),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1700),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1656),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1719),
.B(n_1634),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1645),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1652),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_SL g1760 ( 
.A(n_1611),
.B(n_1655),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1622),
.B(n_1640),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1670),
.B(n_1677),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1624),
.B(n_1616),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1629),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1616),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1749),
.A2(n_1682),
.B1(n_1713),
.B2(n_1690),
.Y(n_1766)
);

OAI21xp33_ASAP7_75t_L g1767 ( 
.A1(n_1749),
.A2(n_1716),
.B(n_1715),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_R g1768 ( 
.A(n_1735),
.B(n_1631),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1735),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1765),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1738),
.Y(n_1771)
);

AOI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1765),
.A2(n_1595),
.B(n_1620),
.Y(n_1772)
);

AOI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1747),
.A2(n_1687),
.B1(n_1705),
.B2(n_1667),
.C(n_1668),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1733),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1738),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1751),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1736),
.A2(n_1603),
.B(n_1671),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1747),
.A2(n_1681),
.B1(n_1712),
.B2(n_1664),
.Y(n_1778)
);

OAI221xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1736),
.A2(n_1709),
.B1(n_1669),
.B2(n_1708),
.C(n_1684),
.Y(n_1779)
);

AOI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1740),
.A2(n_1703),
.B1(n_1665),
.B2(n_1701),
.C1(n_1699),
.C2(n_1686),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1751),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1722),
.B(n_1723),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1721),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1765),
.A2(n_1609),
.B1(n_1604),
.B2(n_1691),
.C(n_1693),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1739),
.A2(n_1675),
.B1(n_1661),
.B2(n_1597),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1724),
.B(n_1615),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1740),
.A2(n_1607),
.B1(n_1763),
.B2(n_1739),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_R g1788 ( 
.A(n_1739),
.B(n_1642),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1721),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1726),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1732),
.Y(n_1791)
);

AO21x2_ASAP7_75t_L g1792 ( 
.A1(n_1742),
.A2(n_1623),
.B(n_1636),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1732),
.Y(n_1793)
);

OAI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1763),
.A2(n_1692),
.A3(n_1617),
.B(n_1637),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1727),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1745),
.B(n_1610),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1763),
.A2(n_1605),
.B1(n_1618),
.B2(n_1627),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1764),
.A2(n_1635),
.B(n_1633),
.C(n_1628),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1727),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1761),
.A2(n_1764),
.B1(n_1752),
.B2(n_1753),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1727),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1756),
.A2(n_1720),
.B1(n_1639),
.B2(n_1711),
.Y(n_1802)
);

NAND2xp33_ASAP7_75t_SL g1803 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1753),
.A2(n_1619),
.B1(n_1642),
.B2(n_1651),
.C(n_1718),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1737),
.A2(n_1718),
.B1(n_1602),
.B2(n_1614),
.C(n_1720),
.Y(n_1805)
);

OA21x2_ASAP7_75t_L g1806 ( 
.A1(n_1748),
.A2(n_1649),
.B(n_1711),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1746),
.B(n_1614),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_L g1808 ( 
.A(n_1741),
.B(n_1756),
.C(n_1762),
.D(n_1737),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1756),
.A2(n_1741),
.B(n_1761),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1722),
.B(n_1723),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1754),
.Y(n_1811)
);

AOI31xp33_ASAP7_75t_L g1812 ( 
.A1(n_1761),
.A2(n_1698),
.A3(n_1720),
.B(n_1696),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1722),
.B(n_1696),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1752),
.A2(n_1685),
.B1(n_1696),
.B2(n_1596),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1723),
.B(n_1596),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1741),
.B(n_1731),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1782),
.B(n_1737),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1782),
.B(n_1734),
.Y(n_1818)
);

OR2x6_ASAP7_75t_L g1819 ( 
.A(n_1806),
.B(n_1748),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1806),
.B(n_1808),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1810),
.B(n_1734),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1795),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1801),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1729),
.Y(n_1824)
);

OAI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1767),
.A2(n_1750),
.A3(n_1742),
.B(n_1744),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1806),
.B(n_1729),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1774),
.B(n_1742),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1776),
.B(n_1729),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1781),
.B(n_1729),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1767),
.B(n_1760),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1783),
.B(n_1725),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1799),
.B(n_1729),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1790),
.B(n_1743),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1792),
.B(n_1729),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1783),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1789),
.B(n_1725),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1792),
.B(n_1728),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1792),
.B(n_1728),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1790),
.B(n_1728),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1789),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1770),
.B(n_1760),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1815),
.B(n_1744),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1791),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1770),
.B(n_1759),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1843),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1840),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1840),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1811),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1843),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1843),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1809),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1770),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1840),
.Y(n_1855)
);

NOR2xp67_ASAP7_75t_L g1856 ( 
.A(n_1820),
.B(n_1808),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1843),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1820),
.B(n_1771),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1817),
.B(n_1813),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1817),
.B(n_1813),
.Y(n_1860)
);

INVxp67_ASAP7_75t_SL g1861 ( 
.A(n_1845),
.Y(n_1861)
);

INVxp67_ASAP7_75t_SL g1862 ( 
.A(n_1845),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1820),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1835),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1840),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1817),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1840),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1825),
.A2(n_1830),
.B1(n_1777),
.B2(n_1773),
.C(n_1785),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1817),
.B(n_1816),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1835),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1842),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1835),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1820),
.B(n_1775),
.Y(n_1873)
);

NOR2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1824),
.B(n_1769),
.Y(n_1874)
);

AOI32xp33_ASAP7_75t_L g1875 ( 
.A1(n_1830),
.A2(n_1766),
.A3(n_1787),
.B1(n_1778),
.B2(n_1770),
.Y(n_1875)
);

NAND2x1_ASAP7_75t_L g1876 ( 
.A(n_1837),
.B(n_1816),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1835),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1835),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1846),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1823),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1846),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1842),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1823),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1842),
.B(n_1815),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1786),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1846),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1842),
.B(n_1744),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1846),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1847),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1868),
.A2(n_1830),
.B(n_1779),
.C(n_1784),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1837),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1848),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1853),
.B(n_1837),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1847),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1875),
.A2(n_1838),
.B1(n_1800),
.B2(n_1834),
.C(n_1804),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1876),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1851),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_L g1899 ( 
.A(n_1875),
.B(n_1814),
.C(n_1780),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1850),
.B(n_1685),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1888),
.B(n_1838),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1851),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1888),
.B(n_1838),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1852),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1852),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1874),
.B(n_1838),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1869),
.B(n_1818),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1861),
.B(n_1841),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1857),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1854),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1857),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1864),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1869),
.B(n_1834),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1862),
.B(n_1762),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1885),
.B(n_1831),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1885),
.B(n_1831),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1848),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1864),
.Y(n_1918)
);

NOR3xp33_ASAP7_75t_L g1919 ( 
.A(n_1856),
.B(n_1798),
.C(n_1772),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1856),
.B(n_1818),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1870),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1858),
.B(n_1831),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1848),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1870),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1872),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1884),
.B(n_1818),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1859),
.B(n_1796),
.Y(n_1927)
);

AND2x2_ASAP7_75t_SL g1928 ( 
.A(n_1858),
.B(n_1841),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_1876),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1859),
.B(n_1841),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1855),
.Y(n_1931)
);

NAND2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1866),
.B(n_1768),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1860),
.B(n_1754),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1855),
.Y(n_1934)
);

OAI21xp33_ASAP7_75t_L g1935 ( 
.A1(n_1919),
.A2(n_1899),
.B(n_1896),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1932),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1897),
.B(n_1863),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1927),
.B(n_1884),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1907),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1890),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1914),
.B(n_1860),
.Y(n_1941)
);

OAI31xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1900),
.A2(n_1863),
.A3(n_1834),
.B(n_1871),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1892),
.B(n_1854),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1891),
.A2(n_1772),
.B(n_1824),
.Y(n_1944)
);

OAI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1894),
.A2(n_1826),
.B(n_1824),
.Y(n_1945)
);

AOI32xp33_ASAP7_75t_L g1946 ( 
.A1(n_1892),
.A2(n_1882),
.A3(n_1797),
.B1(n_1803),
.B2(n_1873),
.Y(n_1946)
);

NAND2x1_ASAP7_75t_L g1947 ( 
.A(n_1897),
.B(n_1854),
.Y(n_1947)
);

OAI32xp33_ASAP7_75t_L g1948 ( 
.A1(n_1929),
.A2(n_1788),
.A3(n_1873),
.B1(n_1824),
.B2(n_1826),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1906),
.A2(n_1794),
.B(n_1826),
.C(n_1802),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1933),
.B(n_1845),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1908),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1928),
.B(n_1818),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1910),
.B(n_1854),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1890),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1895),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1907),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1920),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1906),
.B(n_1854),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1928),
.A2(n_1812),
.B1(n_1805),
.B2(n_1731),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1897),
.A2(n_1826),
.B(n_1794),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1910),
.B(n_1886),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1895),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1922),
.B(n_1836),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1922),
.B(n_1836),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1898),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1910),
.B(n_1886),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1898),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1913),
.B(n_1849),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1902),
.Y(n_1969)
);

CKINVDCx16_ASAP7_75t_R g1970 ( 
.A(n_1920),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_SL g1971 ( 
.A1(n_1913),
.A2(n_1752),
.B1(n_1730),
.B2(n_1750),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1955),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1935),
.B(n_1930),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1936),
.B(n_1913),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1946),
.B(n_1903),
.C(n_1901),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1941),
.B(n_1915),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1951),
.B(n_1926),
.Y(n_1977)
);

AND4x1_ASAP7_75t_L g1978 ( 
.A(n_1949),
.B(n_1926),
.C(n_1807),
.D(n_1904),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1938),
.B(n_1915),
.Y(n_1979)
);

OAI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1942),
.A2(n_1916),
.B1(n_1819),
.B2(n_1911),
.C(n_1905),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1970),
.B(n_1821),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1957),
.B(n_1916),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1948),
.B(n_1746),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_L g1984 ( 
.A(n_1944),
.B(n_1904),
.C(n_1902),
.Y(n_1984)
);

O2A1O1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1948),
.A2(n_1819),
.B(n_1849),
.C(n_1867),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1947),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1955),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1959),
.A2(n_1752),
.B1(n_1750),
.B2(n_1819),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1971),
.A2(n_1819),
.B1(n_1833),
.B2(n_1755),
.Y(n_1989)
);

NOR3xp33_ASAP7_75t_L g1990 ( 
.A(n_1960),
.B(n_1905),
.C(n_1909),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1937),
.A2(n_1752),
.B1(n_1819),
.B2(n_1730),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1940),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1954),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1950),
.B(n_1827),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1943),
.B(n_1821),
.Y(n_1995)
);

AOI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1945),
.A2(n_1819),
.B1(n_1730),
.B2(n_1757),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1962),
.Y(n_1997)
);

NAND2x1_ASAP7_75t_L g1998 ( 
.A(n_1968),
.B(n_1867),
.Y(n_1998)
);

NAND4xp25_ASAP7_75t_SL g1999 ( 
.A(n_1990),
.B(n_1943),
.C(n_1958),
.D(n_1952),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1998),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_1939),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1972),
.Y(n_2002)
);

XNOR2xp5_ASAP7_75t_L g2003 ( 
.A(n_1978),
.B(n_1958),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1974),
.B(n_1939),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1986),
.B(n_1961),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1982),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1973),
.B(n_1953),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1987),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1981),
.B(n_1995),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1993),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_SL g2011 ( 
.A(n_1985),
.B(n_1953),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1997),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_1984),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1983),
.B(n_1956),
.Y(n_2014)
);

NAND2x1_ASAP7_75t_L g2015 ( 
.A(n_1991),
.B(n_1968),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1992),
.Y(n_2016)
);

OAI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1977),
.A2(n_1956),
.B(n_1961),
.Y(n_2017)
);

AOI211xp5_ASAP7_75t_L g2018 ( 
.A1(n_1980),
.A2(n_1966),
.B(n_1967),
.C(n_1969),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2006),
.B(n_1992),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_2005),
.B(n_1966),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2005),
.B(n_1979),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_2009),
.B(n_1968),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_SL g2023 ( 
.A(n_1999),
.B(n_2007),
.C(n_2017),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_2003),
.B(n_1991),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2009),
.B(n_1976),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_2003),
.B(n_1975),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2008),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_2000),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2008),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2013),
.B(n_1988),
.Y(n_2030)
);

HB1xp67_ASAP7_75t_L g2031 ( 
.A(n_2028),
.Y(n_2031)
);

OAI211xp5_ASAP7_75t_SL g2032 ( 
.A1(n_2023),
.A2(n_2018),
.B(n_2001),
.C(n_2016),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_2026),
.A2(n_2011),
.B1(n_2015),
.B2(n_2014),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_SL g2034 ( 
.A1(n_2024),
.A2(n_2004),
.B1(n_2000),
.B2(n_2010),
.C(n_2012),
.Y(n_2034)
);

AOI222xp33_ASAP7_75t_L g2035 ( 
.A1(n_2024),
.A2(n_1975),
.B1(n_2002),
.B2(n_1989),
.C1(n_1996),
.C2(n_2015),
.Y(n_2035)
);

AND3x1_ASAP7_75t_L g2036 ( 
.A(n_2020),
.B(n_2002),
.C(n_1996),
.Y(n_2036)
);

AO21x1_ASAP7_75t_L g2037 ( 
.A1(n_2027),
.A2(n_2029),
.B(n_2019),
.Y(n_2037)
);

AOI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2030),
.A2(n_1947),
.B1(n_1965),
.B2(n_1994),
.C(n_1924),
.Y(n_2038)
);

NAND4xp25_ASAP7_75t_L g2039 ( 
.A(n_2021),
.B(n_2025),
.C(n_2020),
.D(n_2022),
.Y(n_2039)
);

AOI221xp5_ASAP7_75t_SL g2040 ( 
.A1(n_2022),
.A2(n_1893),
.B1(n_1923),
.B2(n_1934),
.C(n_1931),
.Y(n_2040)
);

NAND3xp33_ASAP7_75t_SL g2041 ( 
.A(n_2028),
.B(n_1964),
.C(n_1963),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2031),
.B(n_1963),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2033),
.B(n_1964),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2037),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_2039),
.B(n_1909),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2032),
.A2(n_1911),
.B1(n_1912),
.B2(n_1730),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2041),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2035),
.A2(n_1730),
.B1(n_1918),
.B2(n_1925),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_2036),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2042),
.Y(n_2050)
);

NOR2x1p5_ASAP7_75t_L g2051 ( 
.A(n_2047),
.B(n_2034),
.Y(n_2051)
);

A2O1A1Ixp33_ASAP7_75t_SL g2052 ( 
.A1(n_2044),
.A2(n_2038),
.B(n_2040),
.C(n_1934),
.Y(n_2052)
);

NAND2xp33_ASAP7_75t_R g2053 ( 
.A(n_2043),
.B(n_1893),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_L g2054 ( 
.A(n_2049),
.B(n_1931),
.C(n_1923),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2045),
.Y(n_2055)
);

OAI211xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2048),
.A2(n_1925),
.B(n_1924),
.C(n_1921),
.Y(n_2056)
);

AND3x4_ASAP7_75t_L g2057 ( 
.A(n_2046),
.B(n_1917),
.C(n_1833),
.Y(n_2057)
);

OAI22x1_ASAP7_75t_L g2058 ( 
.A1(n_2051),
.A2(n_1917),
.B1(n_1855),
.B2(n_1865),
.Y(n_2058)
);

NOR2x1p5_ASAP7_75t_L g2059 ( 
.A(n_2055),
.B(n_1918),
.Y(n_2059)
);

OR3x1_ASAP7_75t_L g2060 ( 
.A(n_2056),
.B(n_1921),
.C(n_1889),
.Y(n_2060)
);

AND4x1_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_1828),
.C(n_1829),
.D(n_1839),
.Y(n_2061)
);

NAND4xp25_ASAP7_75t_L g2062 ( 
.A(n_2052),
.B(n_1786),
.C(n_1596),
.D(n_1757),
.Y(n_2062)
);

NOR3xp33_ASAP7_75t_L g2063 ( 
.A(n_2054),
.B(n_1758),
.C(n_1832),
.Y(n_2063)
);

XOR2xp5_ASAP7_75t_L g2064 ( 
.A(n_2058),
.B(n_2062),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2060),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_2059),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_2061),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2067),
.A2(n_2057),
.B1(n_2053),
.B2(n_2063),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2068),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_2069),
.Y(n_2070)
);

OAI332xp33_ASAP7_75t_L g2071 ( 
.A1(n_2069),
.A2(n_2066),
.A3(n_2065),
.B1(n_2064),
.B2(n_1865),
.B3(n_1887),
.C1(n_1889),
.C2(n_1879),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1865),
.B(n_1878),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2070),
.A2(n_1887),
.B1(n_1877),
.B2(n_1881),
.C(n_1878),
.Y(n_2073)
);

OAI222xp33_ASAP7_75t_L g2074 ( 
.A1(n_2072),
.A2(n_1881),
.B1(n_1879),
.B2(n_1877),
.C1(n_1872),
.C2(n_1880),
.Y(n_2074)
);

AO21x2_ASAP7_75t_L g2075 ( 
.A1(n_2073),
.A2(n_1883),
.B(n_1880),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2075),
.A2(n_1883),
.B1(n_1880),
.B2(n_1839),
.Y(n_2076)
);

AOI221xp5_ASAP7_75t_L g2077 ( 
.A1(n_2076),
.A2(n_2074),
.B1(n_2075),
.B2(n_1883),
.C(n_1822),
.Y(n_2077)
);

AOI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_2077),
.A2(n_1836),
.B(n_1829),
.C(n_1828),
.Y(n_2078)
);


endmodule