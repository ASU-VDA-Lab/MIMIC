module fake_jpeg_22645_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_SL g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_3),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

AO22x1_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_17),
.B1(n_10),
.B2(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_20),
.B1(n_8),
.B2(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_9),
.B1(n_6),
.B2(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_13),
.C(n_15),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_17),
.B1(n_11),
.B2(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_8),
.Y(n_28)
);

XNOR2x1_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_23),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_19),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_5),
.B(n_4),
.Y(n_32)
);

NOR5xp2_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_5),
.C(n_18),
.D(n_31),
.E(n_33),
.Y(n_34)
);


endmodule