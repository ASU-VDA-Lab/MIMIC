module real_jpeg_25966_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_34),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_34),
.B1(n_53),
.B2(n_56),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_34),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_59),
.B(n_201),
.C(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_57),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_38),
.B(n_44),
.C(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_3),
.B(n_25),
.C(n_28),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_3),
.B(n_96),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_167),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_3),
.B(n_27),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_4),
.A2(n_42),
.B1(n_44),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_22),
.B1(n_26),
.B2(n_49),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_49),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_53),
.B1(n_64),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_8),
.A2(n_42),
.B1(n_44),
.B2(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_143),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_143),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_42),
.B1(n_44),
.B2(n_54),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_10),
.A2(n_22),
.B1(n_26),
.B2(n_54),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_54),
.Y(n_163)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_11),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_11),
.B(n_256),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_91),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_89),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_76),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_15),
.B(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_67),
.B2(n_75),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_50),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_18),
.A2(n_35),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_18),
.A2(n_80),
.B1(n_85),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_18),
.A2(n_80),
.B1(n_185),
.B2(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_19),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_20),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_20),
.B(n_33),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_20),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_22),
.B(n_244),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_26),
.A2(n_34),
.B(n_39),
.Y(n_227)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_27),
.B(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_27),
.B(n_231),
.Y(n_241)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_28),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_28),
.B(n_267),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_31),
.B(n_32),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_31),
.A2(n_100),
.B(n_115),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_34),
.A2(n_44),
.B(n_58),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_36),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_40),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_37),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_41),
.B(n_86),
.Y(n_137)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_87),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_45),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_46),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_60),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_53),
.Y(n_203)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_57),
.B(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_57),
.B(n_142),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_61),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_62),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_68),
.B(n_160),
.C(n_170),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_68),
.A2(n_73),
.B1(n_170),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_70),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_72),
.B(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_84),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_77),
.A2(n_81),
.B1(n_105),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.C(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_80),
.B(n_183),
.C(n_185),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_82),
.B(n_171),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_84),
.B(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_88),
.B(n_194),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI211xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_144),
.B(n_149),
.C(n_311),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_121),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_121),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_93),
.B(n_146),
.Y(n_311)
);

FAx1_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.CI(n_107),
.CON(n_93),
.SN(n_93)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_95),
.B(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_96),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_98),
.B(n_229),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_100),
.B(n_241),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B(n_117),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_114),
.B1(n_125),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_108),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_108),
.A2(n_125),
.B1(n_226),
.B2(n_283),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B(n_112),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_109),
.B(n_112),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_109),
.B(n_255),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_116),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_116),
.B(n_230),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.C(n_138),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_129),
.B(n_134),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_130),
.B(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_132),
.A2(n_163),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_132),
.B(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_137),
.B(n_187),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_150),
.C(n_151),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_175),
.B(n_310),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_172),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_153),
.B(n_172),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_154),
.B(n_157),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_159),
.B(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_160),
.A2(n_161),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_168),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_165),
.B(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_170),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_305),
.B(n_309),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_219),
.B(n_292),
.C(n_304),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_207),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_178),
.B(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_191),
.B2(n_206),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_189),
.B2(n_190),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_181),
.B(n_190),
.C(n_206),
.Y(n_293)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_184),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_188),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_193),
.B(n_198),
.C(n_199),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_196),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_204),
.Y(n_213)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_209),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_291),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_235),
.B(n_290),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_232),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_222),
.B(n_232),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_228),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_226),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_285),
.B(n_289),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_276),
.B(n_284),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_258),
.B(n_275),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_239),
.B(n_245),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_242),
.B1(n_243),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_252),
.B2(n_257),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_251),
.C(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_264),
.B(n_274),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_270),
.B(n_273),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_271),
.B(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_301),
.B2(n_302),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_302),
.C(n_303),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_306),
.B(n_307),
.Y(n_309)
);


endmodule