module fake_aes_132_n_672 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_672);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_672;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_38), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_6), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_11), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_8), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_37), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_7), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_56), .Y(n_87) );
CKINVDCx14_ASAP7_75t_R g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_45), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_15), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_21), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_67), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_59), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_69), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_33), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_28), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_0), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_20), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_30), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_54), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_51), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_46), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_36), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_29), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_7), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_24), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_44), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_43), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_9), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_16), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_90), .B(n_1), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_119), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_88), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_106), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_79), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_84), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_106), .B(n_86), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_92), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_102), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_122), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_123), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_77), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_111), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_101), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
BUFx10_ASAP7_75t_L g149 ( .A(n_103), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_87), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_78), .B(n_2), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g154 ( .A(n_85), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_109), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_78), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_80), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_80), .B(n_93), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_93), .B(n_3), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_131), .B(n_121), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_136), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_131), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_146), .B(n_110), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_158), .B(n_108), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_157), .B(n_121), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_126), .Y(n_178) );
OR2x2_ASAP7_75t_SL g179 ( .A(n_154), .B(n_120), .Y(n_179) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_161), .B(n_120), .C(n_98), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_149), .B(n_99), .Y(n_181) );
INVxp67_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_134), .B(n_96), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_158), .B(n_97), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_137), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_141), .B(n_99), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_162), .B(n_97), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_152), .A2(n_116), .B(n_98), .C(n_114), .Y(n_195) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_124), .B(n_105), .C(n_113), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_162), .B(n_113), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_162), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_124), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_139), .B(n_105), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_128), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_128), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_165), .B(n_114), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_138), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_139), .A2(n_117), .B(n_96), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_144), .Y(n_217) );
INVx3_ASAP7_75t_R g218 ( .A(n_150), .Y(n_218) );
INVx8_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_140), .Y(n_222) );
AND2x6_ASAP7_75t_L g223 ( .A(n_163), .B(n_100), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_142), .B(n_117), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_145), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_204), .B(n_142), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_194), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_194), .Y(n_229) );
NAND3xp33_ASAP7_75t_SL g230 ( .A(n_222), .B(n_152), .C(n_132), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_198), .Y(n_231) );
BUFx10_ASAP7_75t_L g232 ( .A(n_223), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_178), .Y(n_235) );
BUFx12f_ASAP7_75t_L g236 ( .A(n_178), .Y(n_236) );
OR2x6_ASAP7_75t_SL g237 ( .A(n_169), .B(n_143), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_197), .B(n_143), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_203), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_179), .B(n_153), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_177), .B(n_153), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_184), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_176), .B(n_155), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_189), .Y(n_246) );
NOR3xp33_ASAP7_75t_SL g247 ( .A(n_180), .B(n_82), .C(n_91), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_219), .B(n_165), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_189), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_169), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_223), .A2(n_164), .B1(n_160), .B2(n_155), .Y(n_252) );
INVx8_ASAP7_75t_L g253 ( .A(n_219), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_223), .A2(n_164), .B1(n_160), .B2(n_156), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_195), .A2(n_156), .B1(n_116), .B2(n_151), .C(n_150), .Y(n_256) );
BUFx4f_ASAP7_75t_L g257 ( .A(n_184), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_200), .B(n_159), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_203), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_206), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_199), .B(n_159), .Y(n_263) );
CKINVDCx11_ASAP7_75t_R g264 ( .A(n_213), .Y(n_264) );
INVx5_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_219), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_219), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_197), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_197), .B(n_159), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_209), .B(n_151), .Y(n_271) );
INVx5_ASAP7_75t_L g272 ( .A(n_184), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_186), .B(n_209), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
NOR3xp33_ASAP7_75t_SL g277 ( .A(n_175), .B(n_118), .C(n_107), .Y(n_277) );
XNOR2xp5_ASAP7_75t_L g278 ( .A(n_213), .B(n_118), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_171), .Y(n_279) );
NOR3xp33_ASAP7_75t_SL g280 ( .A(n_196), .B(n_100), .C(n_104), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_172), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_209), .B(n_151), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_193), .A2(n_214), .B(n_205), .C(n_221), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_182), .Y(n_284) );
CKINVDCx6p67_ASAP7_75t_R g285 ( .A(n_200), .Y(n_285) );
BUFx12f_ASAP7_75t_L g286 ( .A(n_179), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_172), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
AO21x1_ASAP7_75t_L g289 ( .A1(n_242), .A2(n_104), .B(n_112), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_253), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_283), .A2(n_211), .B(n_208), .C(n_210), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_238), .B(n_223), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_238), .B(n_223), .Y(n_296) );
INVx5_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_231), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_236), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_231), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_268), .A2(n_220), .B1(n_183), .B2(n_215), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_264), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_257), .B(n_205), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_253), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_238), .B(n_223), .Y(n_308) );
HAxp5_ASAP7_75t_L g309 ( .A(n_237), .B(n_192), .CON(n_309), .SN(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_236), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_241), .B(n_181), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_227), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_235), .B(n_208), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_264), .Y(n_317) );
O2A1O1Ixp5_ASAP7_75t_L g318 ( .A1(n_283), .A2(n_224), .B(n_168), .C(n_207), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_268), .A2(n_223), .B1(n_184), .B2(n_220), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_226), .A2(n_210), .B1(n_221), .B2(n_211), .C(n_216), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_232), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_285), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_237), .Y(n_323) );
AOI21x1_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_173), .B(n_174), .Y(n_324) );
BUFx6f_ASAP7_75t_SL g325 ( .A(n_267), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_226), .B(n_215), .Y(n_326) );
AND2x6_ASAP7_75t_L g327 ( .A(n_252), .B(n_173), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_241), .A2(n_184), .B1(n_274), .B2(n_256), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_248), .B(n_184), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_285), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_230), .A2(n_166), .B1(n_185), .B2(n_174), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_229), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_251), .B(n_112), .C(n_115), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_267), .B(n_166), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_286), .A2(n_166), .B1(n_185), .B2(n_207), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_245), .B(n_166), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_305), .B(n_254), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_323), .A2(n_286), .B1(n_235), .B2(n_266), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_311), .B(n_277), .Y(n_341) );
INVx6_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_311), .B(n_282), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_326), .B(n_259), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_293), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_328), .B(n_259), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_333), .A2(n_266), .B1(n_228), .B2(n_278), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_305), .B(n_271), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_300), .A2(n_228), .B1(n_233), .B2(n_246), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_295), .A2(n_233), .B1(n_249), .B2(n_240), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_290), .B(n_270), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_328), .B(n_280), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_298), .A2(n_251), .B1(n_257), .B2(n_243), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_297), .B(n_291), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_297), .B(n_243), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_302), .A2(n_166), .B1(n_265), .B2(n_272), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_297), .B(n_261), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_316), .B(n_255), .Y(n_362) );
INVx5_ASAP7_75t_L g363 ( .A(n_297), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_327), .A2(n_263), .B1(n_247), .B2(n_166), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_336), .A2(n_275), .B(n_287), .Y(n_366) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_302), .A2(n_130), .B1(n_133), .B2(n_150), .C1(n_216), .C2(n_281), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_320), .B(n_273), .Y(n_368) );
OAI33xp33_ASAP7_75t_L g369 ( .A1(n_341), .A2(n_130), .A3(n_133), .B1(n_309), .B2(n_115), .B3(n_301), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_356), .A2(n_289), .B(n_318), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_367), .B(n_322), .Y(n_372) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_363), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_367), .B(n_332), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_363), .B(n_291), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_364), .B(n_330), .Y(n_376) );
AOI221x1_ASAP7_75t_L g377 ( .A1(n_347), .A2(n_292), .B1(n_309), .B2(n_148), .C(n_147), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_339), .B(n_273), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_365), .A2(n_319), .B(n_292), .C(n_331), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_365), .B(n_148), .C(n_147), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_364), .B(n_330), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_362), .B(n_294), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_351), .B(n_327), .Y(n_384) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_348), .B(n_147), .C(n_148), .D(n_145), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_366), .A2(n_324), .B(n_329), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_335), .B(n_308), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_363), .B(n_317), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_344), .A2(n_317), .B1(n_310), .B2(n_299), .C(n_296), .Y(n_393) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_368), .A2(n_279), .B(n_188), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_345), .A2(n_307), .B1(n_314), .B2(n_334), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_370), .B(n_351), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_350), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_373), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_338), .B1(n_350), .B2(n_355), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_374), .A2(n_362), .B1(n_338), .B2(n_363), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_377), .B(n_352), .C(n_354), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_390), .Y(n_403) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_373), .B(n_343), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_388), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_170), .B(n_187), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_391), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_381), .B(n_327), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_381), .B(n_327), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_390), .B(n_327), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_394), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_394), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_369), .A2(n_355), .B1(n_353), .B2(n_340), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_394), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_371), .A2(n_299), .B1(n_310), .B2(n_325), .C(n_207), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_391), .Y(n_421) );
NAND4xp25_ASAP7_75t_SL g422 ( .A(n_393), .B(n_360), .C(n_361), .D(n_353), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_373), .B(n_343), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_376), .A2(n_343), .B1(n_307), .B2(n_337), .C(n_342), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_382), .A2(n_343), .B1(n_337), .B2(n_342), .C(n_361), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_383), .B(n_358), .Y(n_426) );
NOR4xp25_ASAP7_75t_SL g427 ( .A(n_392), .B(n_342), .C(n_325), .D(n_8), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_385), .A2(n_358), .B1(n_342), .B2(n_337), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_379), .A2(n_395), .A3(n_383), .B(n_375), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_396), .B(n_395), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_385), .B1(n_358), .B2(n_380), .Y(n_432) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_427), .B(n_373), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_398), .B(n_386), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_398), .B(n_386), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_405), .A2(n_380), .B1(n_389), .B2(n_212), .C(n_217), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_396), .B(n_386), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_415), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_403), .B(n_386), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
OAI33xp33_ASAP7_75t_L g448 ( .A1(n_401), .A2(n_4), .A3(n_5), .B1(n_9), .B2(n_10), .B3(n_12), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_418), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_414), .A2(n_375), .B1(n_386), .B2(n_225), .C(n_217), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_401), .A2(n_212), .B1(n_225), .B2(n_358), .C(n_188), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_399), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_399), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_375), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_416), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_397), .B(n_387), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_419), .A2(n_201), .B(n_170), .C(n_187), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_397), .B(n_387), .Y(n_462) );
NAND2xp67_ASAP7_75t_L g463 ( .A(n_409), .B(n_4), .Y(n_463) );
NOR2xp33_ASAP7_75t_R g464 ( .A(n_422), .B(n_10), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_430), .B(n_387), .Y(n_465) );
OR2x6_ASAP7_75t_SL g466 ( .A(n_421), .B(n_13), .Y(n_466) );
AOI33xp33_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_191), .A3(n_201), .B1(n_202), .B2(n_16), .B3(n_18), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_13), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_417), .B(n_14), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_421), .B(n_359), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_422), .A2(n_359), .A3(n_334), .B(n_191), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_14), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_429), .A2(n_202), .B1(n_334), .B2(n_359), .C(n_276), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_15), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_429), .B(n_359), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_409), .B(n_18), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_447), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_462), .B(n_410), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_438), .B(n_410), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_479), .B(n_411), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_466), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_460), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_479), .B(n_426), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_468), .B(n_426), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_441), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_459), .B(n_406), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_442), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_465), .B(n_423), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_445), .B(n_404), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_442), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_447), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_446), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_473), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_459), .B(n_406), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_473), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_477), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_476), .B(n_404), .Y(n_508) );
NAND2xp33_ASAP7_75t_SL g509 ( .A(n_464), .B(n_427), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_434), .B(n_406), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_477), .B(n_428), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_431), .B(n_423), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_476), .B(n_423), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_446), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_434), .B(n_406), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_456), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_441), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_443), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_435), .B(n_399), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_443), .B(n_399), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_435), .B(n_399), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_465), .B(n_399), .Y(n_522) );
NOR4xp25_ASAP7_75t_SL g523 ( .A(n_433), .B(n_425), .C(n_424), .D(n_402), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_444), .B(n_402), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_469), .B(n_19), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_444), .B(n_19), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_465), .B(n_68), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_465), .B(n_20), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_432), .B(n_21), .C(n_276), .D(n_260), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_437), .B(n_166), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_458), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_458), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_454), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_470), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_480), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_517), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_490), .A2(n_466), .B1(n_432), .B2(n_478), .Y(n_539) );
AOI32xp33_ASAP7_75t_L g540 ( .A1(n_509), .A2(n_470), .A3(n_450), .B1(n_456), .B2(n_451), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_480), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g542 ( .A1(n_509), .A2(n_531), .B1(n_525), .B2(n_471), .C(n_506), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_504), .B(n_463), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g544 ( .A1(n_530), .A2(n_489), .B(n_463), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_527), .A2(n_475), .B1(n_472), .B2(n_454), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_487), .A2(n_436), .B1(n_474), .B2(n_472), .C(n_475), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_536), .B(n_452), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_511), .A2(n_452), .B1(n_455), .B2(n_453), .C(n_461), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_483), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_523), .A2(n_453), .B(n_455), .C(n_448), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_507), .B(n_467), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_484), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_485), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_516), .A2(n_470), .B1(n_453), .B2(n_312), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_495), .Y(n_557) );
AOI31xp33_ASAP7_75t_L g558 ( .A1(n_530), .A2(n_22), .A3(n_26), .B(n_27), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_518), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_524), .B(n_262), .C(n_288), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_527), .A2(n_243), .B(n_265), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_526), .B(n_31), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_512), .B(n_32), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_519), .B(n_34), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_502), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_529), .A2(n_265), .B(n_272), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_502), .A2(n_260), .B1(n_239), .B2(n_244), .C(n_258), .Y(n_568) );
INVxp33_ASAP7_75t_L g569 ( .A(n_484), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_494), .A2(n_312), .B1(n_315), .B2(n_321), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_528), .A2(n_239), .B1(n_244), .B2(n_250), .C(n_258), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_491), .B(n_39), .Y(n_572) );
O2A1O1Ixp33_ASAP7_75t_SL g573 ( .A1(n_500), .A2(n_41), .B(n_42), .C(n_47), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_493), .B(n_48), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_486), .B(n_49), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_500), .Y(n_576) );
OAI22xp33_ASAP7_75t_SL g577 ( .A1(n_482), .A2(n_272), .B1(n_265), .B2(n_243), .Y(n_577) );
AOI311xp33_ASAP7_75t_L g578 ( .A1(n_497), .A2(n_50), .A3(n_53), .B(n_55), .C(n_57), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_534), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_498), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_482), .B(n_272), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_492), .A2(n_250), .B1(n_288), .B2(n_262), .C(n_312), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_529), .A2(n_321), .B(n_315), .C(n_304), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_519), .B(n_60), .Y(n_584) );
AOI22x1_ASAP7_75t_L g585 ( .A1(n_529), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_537), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_553), .B(n_522), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_542), .B(n_482), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_576), .B(n_522), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_538), .B(n_521), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_547), .B(n_521), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_580), .B(n_496), .Y(n_594) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_539), .B(n_508), .Y(n_595) );
XNOR2x1_ASAP7_75t_L g596 ( .A(n_575), .B(n_488), .Y(n_596) );
NAND2x1p5_ASAP7_75t_SL g597 ( .A(n_585), .B(n_496), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_548), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_586), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_544), .A2(n_524), .B(n_499), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_557), .B(n_505), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_581), .B(n_520), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
XOR2x2_ASAP7_75t_L g605 ( .A(n_565), .B(n_499), .Y(n_605) );
AOI211x1_ASAP7_75t_L g606 ( .A1(n_558), .A2(n_513), .B(n_505), .C(n_510), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_550), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_569), .A2(n_499), .B(n_508), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_573), .A2(n_520), .B(n_514), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_567), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_540), .A2(n_510), .B(n_515), .C(n_535), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_543), .B(n_535), .Y(n_613) );
NAND2xp33_ASAP7_75t_R g614 ( .A(n_564), .B(n_515), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_579), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_551), .A2(n_532), .B(n_514), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_545), .B(n_503), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_552), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_545), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_555), .B(n_503), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_560), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_609), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_549), .B(n_573), .C(n_546), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_615), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_595), .B(n_583), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_612), .A2(n_583), .B(n_574), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_600), .A2(n_563), .B(n_574), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_619), .A2(n_563), .B1(n_551), .B2(n_584), .C1(n_572), .C2(n_561), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_614), .A2(n_570), .B1(n_562), .B2(n_581), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_618), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_605), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_601), .B(n_501), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_617), .B(n_566), .Y(n_633) );
OA211x2_ASAP7_75t_L g634 ( .A1(n_608), .A2(n_578), .B(n_582), .C(n_571), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_590), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_610), .A2(n_568), .B(n_501), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_619), .A2(n_577), .A3(n_304), .B1(n_71), .B2(n_72), .C1(n_73), .C2(n_74), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_613), .B(n_65), .Y(n_638) );
AOI211xp5_ASAP7_75t_SL g639 ( .A1(n_616), .A2(n_304), .B(n_76), .C(n_70), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_615), .B(n_262), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_621), .A2(n_597), .B(n_603), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_606), .B(n_597), .C(n_620), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_625), .A2(n_596), .B(n_603), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_634), .A2(n_596), .B1(n_605), .B2(n_607), .Y(n_644) );
NOR4xp75_ASAP7_75t_L g645 ( .A(n_631), .B(n_626), .C(n_627), .D(n_638), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_641), .B(n_621), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_623), .A2(n_598), .B(n_611), .C(n_602), .Y(n_647) );
AOI31xp33_ASAP7_75t_L g648 ( .A1(n_633), .A2(n_603), .A3(n_592), .B(n_593), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_629), .A2(n_591), .B(n_602), .C(n_587), .Y(n_649) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_630), .A2(n_587), .B1(n_591), .B2(n_604), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_622), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_636), .B(n_604), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_635), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_592), .B1(n_588), .B2(n_594), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_639), .A2(n_599), .B(n_588), .Y(n_655) );
OA22x2_ASAP7_75t_L g656 ( .A1(n_624), .A2(n_593), .B1(n_599), .B2(n_218), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_632), .Y(n_657) );
AO22x1_ASAP7_75t_L g658 ( .A1(n_637), .A2(n_272), .B1(n_288), .B2(n_640), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_644), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_651), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_644), .B(n_647), .Y(n_662) );
XOR2xp5_ASAP7_75t_L g663 ( .A(n_657), .B(n_656), .Y(n_663) );
OAI222xp33_ASAP7_75t_L g664 ( .A1(n_660), .A2(n_646), .B1(n_652), .B2(n_654), .C1(n_645), .C2(n_655), .Y(n_664) );
OA22x2_ASAP7_75t_L g665 ( .A1(n_660), .A2(n_643), .B1(n_642), .B2(n_649), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_661), .B(n_653), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_666), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_665), .Y(n_668) );
A2O1A1O1Ixp25_ASAP7_75t_L g669 ( .A1(n_667), .A2(n_662), .B(n_664), .C(n_648), .D(n_659), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_668), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_670), .B(n_667), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_669), .B1(n_663), .B2(n_658), .C(n_650), .Y(n_672) );
endmodule