module real_jpeg_33030_n_21 (n_17, n_8, n_0, n_157, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_147, n_6, n_153, n_151, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_150, n_1, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_155, n_21);

input n_17;
input n_8;
input n_0;
input n_157;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_147;
input n_6;
input n_153;
input n_151;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_21;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_0),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_2),
.B(n_111),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_12),
.B1(n_82),
.B2(n_86),
.C(n_90),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_3),
.B(n_82),
.C(n_86),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_5),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_5),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_71),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_8),
.B(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_11),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_40),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_14),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_84),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_24),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_19),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_19),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_20),
.A2(n_55),
.A3(n_57),
.B1(n_61),
.B2(n_122),
.C1(n_124),
.C2(n_157),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_140),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_139),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_27),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_130),
.B(n_136),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_37),
.B(n_128),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_32),
.B(n_36),
.Y(n_129)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_45),
.B(n_127),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI31xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_74),
.A3(n_109),
.B(n_117),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_60),
.C(n_70),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_48),
.A2(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_70),
.C(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_148),
.Y(n_57)
);

OA21x2_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_104),
.C(n_105),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_94),
.B(n_103),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_153),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_147),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_149),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_150),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_151),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_152),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_154),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_155),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_156),
.Y(n_112)
);


endmodule