module fake_jpeg_2929_n_199 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_22),
.A2(n_20),
.B1(n_32),
.B2(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_43),
.A2(n_63),
.B1(n_69),
.B2(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

NAND2x1_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_54),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_33),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_3),
.C(n_4),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_19),
.B(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_26),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_15),
.B(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_31),
.A2(n_13),
.B(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_17),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_35),
.B1(n_24),
.B2(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_35),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_103),
.B1(n_75),
.B2(n_88),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_24),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_89),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_38),
.A2(n_56),
.B1(n_39),
.B2(n_49),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_115),
.Y(n_145)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_63),
.B1(n_90),
.B2(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_117),
.B1(n_127),
.B2(n_77),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_94),
.B1(n_75),
.B2(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_129),
.B1(n_104),
.B2(n_102),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_76),
.B1(n_97),
.B2(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_125),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_106),
.B1(n_104),
.B2(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_79),
.B1(n_85),
.B2(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_109),
.B1(n_112),
.B2(n_106),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_141),
.B1(n_127),
.B2(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_117),
.B1(n_113),
.B2(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_140),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_84),
.B(n_77),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_142),
.C(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_159),
.B(n_160),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_122),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_162),
.C(n_136),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_140),
.B1(n_145),
.B2(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_161),
.A3(n_124),
.B1(n_142),
.B2(n_85),
.C1(n_132),
.C2(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_122),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_111),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_139),
.B(n_154),
.Y(n_164)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_137),
.B(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_162),
.Y(n_177)
);

OAI322xp33_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_146),
.A3(n_159),
.B1(n_143),
.B2(n_130),
.C1(n_147),
.C2(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_178),
.B1(n_168),
.B2(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_177),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_161),
.B1(n_151),
.B2(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_180),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_118),
.B1(n_125),
.B2(n_79),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_166),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_187),
.B(n_189),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_164),
.B(n_174),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_171),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_185),
.B1(n_176),
.B2(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_172),
.C(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_172),
.C(n_171),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_195),
.C(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_173),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.Y(n_199)
);


endmodule