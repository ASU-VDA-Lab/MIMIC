module fake_netlist_1_837_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_7;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_4), .Y(n_7) );
INVx3_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
INVx3_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_6), .B(n_2), .Y(n_12) );
AOI221x1_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_3), .C(n_4), .Y(n_13) );
OAI21xp5_ASAP7_75t_L g14 ( .A1(n_8), .A2(n_1), .B(n_5), .Y(n_14) );
AOI21xp5_ASAP7_75t_SL g15 ( .A1(n_12), .A2(n_10), .B(n_11), .Y(n_15) );
O2A1O1Ixp5_ASAP7_75t_L g16 ( .A1(n_8), .A2(n_9), .B(n_10), .C(n_11), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_8), .A2(n_9), .B(n_10), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_15), .B(n_9), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_15), .B(n_9), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_14), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_7), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B(n_18), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_20), .B1(n_19), .B2(n_8), .Y(n_24) );
NAND3x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_13), .C(n_16), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_13), .B(n_8), .Y(n_28) );
OAI21xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B(n_27), .Y(n_29) );
endmodule