module fake_jpeg_2093_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_63),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_41),
.C(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_47),
.B1(n_54),
.B2(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_59),
.B1(n_47),
.B2(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_87),
.B1(n_69),
.B2(n_75),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_83),
.B1(n_86),
.B2(n_67),
.Y(n_93)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_55),
.B1(n_46),
.B2(n_44),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_46),
.B1(n_44),
.B2(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_69),
.B1(n_75),
.B2(n_7),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_51),
.B1(n_52),
.B2(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_52),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_37),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_52),
.B(n_3),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_104),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_75),
.B1(n_34),
.B2(n_32),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_85),
.B1(n_19),
.B2(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_76),
.C(n_85),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_25),
.C(n_24),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_78),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_113),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_17),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_23),
.C(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_104),
.B1(n_95),
.B2(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_96),
.B(n_98),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_139),
.B(n_140),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_17),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_135),
.B(n_138),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_18),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_18),
.B(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_132),
.B1(n_145),
.B2(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_150),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_147),
.A2(n_139),
.B1(n_112),
.B2(n_137),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_127),
.B(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_116),
.Y(n_153)
);

AOI321xp33_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_141),
.A3(n_136),
.B1(n_140),
.B2(n_109),
.C(n_111),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_153),
.C(n_151),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_154),
.CI(n_148),
.CON(n_157),
.SN(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_157),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_157),
.Y(n_162)
);


endmodule