module fake_netlist_6_615_n_1775 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1775);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1775;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_46),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_36),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_107),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_11),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_20),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_103),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_28),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_47),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_76),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_95),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_111),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_96),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

BUFx8_ASAP7_75t_SL g198 ( 
.A(n_66),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_126),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_29),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_59),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_45),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_59),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_90),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_99),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_77),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_53),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_19),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_108),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_132),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_131),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_33),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_44),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_93),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_66),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_105),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_106),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_47),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_163),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_67),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_32),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_153),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_33),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_148),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_117),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_118),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_123),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_78),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_46),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_166),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_114),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_71),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_128),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_8),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_53),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_109),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_98),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_161),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_97),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_88),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_115),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_171),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_73),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_167),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_63),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_6),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_79),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_50),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_11),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_152),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_51),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_116),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_113),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_102),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_15),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_34),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_23),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_130),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_127),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_7),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_104),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_129),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_60),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_145),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_120),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_135),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_138),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_159),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_162),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_87),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_15),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_61),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_18),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_62),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_158),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_42),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_7),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_38),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_1),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_94),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_142),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_150),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_51),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_19),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_125),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_64),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_151),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_92),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_62),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_58),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_58),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_49),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_146),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_30),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_140),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_227),
.B(n_0),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_205),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_198),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_178),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_190),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_212),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_184),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_263),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_184),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_2),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_179),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_276),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_180),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_279),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_190),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_182),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_246),
.B(n_2),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_236),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_236),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_236),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_185),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_236),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_236),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_331),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_315),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_196),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_309),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_199),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_241),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_241),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_241),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_203),
.B(n_134),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_241),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_207),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_241),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_208),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_209),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_193),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_193),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_221),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_224),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_270),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_225),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_230),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_232),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_175),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_234),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_176),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_239),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_215),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_189),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_219),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_247),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_215),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_250),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_254),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_255),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_256),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_258),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_189),
.Y(n_426)
);

INVxp33_ASAP7_75t_SL g427 ( 
.A(n_188),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_269),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_R g430 ( 
.A(n_257),
.B(n_5),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_177),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_257),
.B(n_5),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_204),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_357),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_352),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_365),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_350),
.B(n_216),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_368),
.B(n_278),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_432),
.B(n_244),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_372),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_360),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_367),
.A2(n_351),
.B(n_349),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_382),
.B(n_280),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_370),
.B(n_259),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_380),
.B(n_259),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_353),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_384),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_387),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_362),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_388),
.B(n_177),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_366),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_369),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_363),
.A2(n_181),
.B1(n_272),
.B2(n_303),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_378),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_367),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_367),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_385),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_394),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_349),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_364),
.A2(n_183),
.B(n_174),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_354),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_390),
.B(n_192),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_359),
.B(n_201),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_354),
.A2(n_358),
.B(n_356),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_356),
.A2(n_183),
.B(n_174),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_392),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_398),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_399),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_400),
.B(n_201),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_358),
.Y(n_500)
);

NAND2x1_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_242),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_363),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_402),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_371),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_371),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_412),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_381),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_393),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_403),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_442),
.A2(n_401),
.B1(n_348),
.B2(n_197),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_453),
.A2(n_373),
.B1(n_271),
.B2(n_327),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_192),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_479),
.A2(n_442),
.B1(n_453),
.B2(n_271),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_383),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_457),
.B(n_408),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_191),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_457),
.B(n_410),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_427),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_482),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_476),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_478),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_435),
.B(n_383),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_485),
.B(n_191),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_485),
.B(n_213),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_405),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_499),
.B(n_406),
.Y(n_541)
);

NOR2x1p5_ASAP7_75t_L g542 ( 
.A(n_436),
.B(n_355),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_441),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_444),
.B(n_407),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_497),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_486),
.A2(n_246),
.B1(n_327),
.B2(n_343),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g549 ( 
.A1(n_465),
.A2(n_433),
.B1(n_220),
.B2(n_251),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_497),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_477),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_490),
.B(n_197),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_438),
.B(n_386),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_455),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_506),
.B(n_200),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_464),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_448),
.B(n_418),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_497),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_420),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_452),
.B(n_421),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_455),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_446),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_506),
.B(n_412),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_466),
.B(n_425),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_494),
.B(n_200),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_501),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_494),
.A2(n_242),
.B1(n_202),
.B2(n_291),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_501),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_465),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_439),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_439),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_467),
.B(n_397),
.Y(n_588)
);

AND2x2_ASAP7_75t_SL g589 ( 
.A(n_494),
.B(n_213),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_452),
.B(n_409),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_481),
.B(n_411),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_443),
.B(n_416),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_508),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_473),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_445),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_496),
.B(n_391),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_502),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_445),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_447),
.B(n_431),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_447),
.B(n_434),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_454),
.B(n_434),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_509),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_498),
.A2(n_302),
.B1(n_295),
.B2(n_293),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_503),
.A2(n_265),
.B1(n_321),
.B2(n_287),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_473),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_509),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_459),
.B(n_416),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_440),
.B(n_415),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_469),
.A2(n_222),
.B(n_206),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_461),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_451),
.B(n_229),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_461),
.B(n_431),
.Y(n_621)
);

BUFx8_ASAP7_75t_SL g622 ( 
.A(n_437),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_458),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_462),
.B(n_431),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_458),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_469),
.A2(n_202),
.B1(n_249),
.B2(n_291),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_462),
.B(n_419),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_458),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_463),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_463),
.B(n_417),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_471),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_471),
.B(n_206),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_483),
.B(n_431),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_483),
.A2(n_249),
.B1(n_204),
.B2(n_294),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_484),
.B(n_429),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_484),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_458),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_487),
.B(n_194),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_487),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_492),
.A2(n_336),
.B1(n_286),
.B2(n_313),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_458),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_495),
.B(n_284),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_513),
.B(n_270),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_513),
.B(n_270),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_529),
.B(n_253),
.C(n_413),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_524),
.A2(n_424),
.B1(n_186),
.B2(n_288),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_559),
.B(n_187),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_573),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_573),
.Y(n_652)
);

OAI22x1_ASAP7_75t_L g653 ( 
.A1(n_641),
.A2(n_285),
.B1(n_217),
.B2(n_346),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_474),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_518),
.B(n_474),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_600),
.B(n_426),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_513),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_524),
.A2(n_312),
.B1(n_282),
.B2(n_283),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_614),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_526),
.B(n_474),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_526),
.B(n_474),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_524),
.B(n_474),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_566),
.B(n_331),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_524),
.A2(n_316),
.B1(n_296),
.B2(n_298),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_520),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_614),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_589),
.A2(n_304),
.B1(n_297),
.B2(n_294),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_512),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_589),
.A2(n_335),
.B1(n_297),
.B2(n_290),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_566),
.B(n_331),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_524),
.B(n_451),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_524),
.B(n_451),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_520),
.B(n_223),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_539),
.B(n_228),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_543),
.B(n_541),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_331),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_519),
.A2(n_318),
.B1(n_299),
.B2(n_301),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_623),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_523),
.B(n_233),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_456),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_544),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_600),
.B(n_210),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_543),
.B(n_305),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_525),
.B(n_243),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_594),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_512),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_566),
.B(n_331),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_623),
.Y(n_689)
);

INVx8_ASAP7_75t_L g690 ( 
.A(n_632),
.Y(n_690)
);

NAND2x1_ASAP7_75t_L g691 ( 
.A(n_577),
.B(n_460),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_569),
.B(n_331),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_540),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_604),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_511),
.B(n_306),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_585),
.B(n_460),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_587),
.B(n_226),
.Y(n_699)
);

INVxp33_ASAP7_75t_SL g700 ( 
.A(n_555),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_511),
.A2(n_248),
.B(n_210),
.C(n_211),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_563),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_535),
.B(n_260),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_569),
.B(n_229),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_623),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_519),
.A2(n_320),
.B1(n_308),
.B2(n_319),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_587),
.B(n_226),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_544),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_540),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_532),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_553),
.A2(n_240),
.B1(n_238),
.B2(n_237),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_616),
.B(n_330),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_607),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_548),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_627),
.B(n_261),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_576),
.A2(n_240),
.B(n_218),
.C(n_237),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_475),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_553),
.A2(n_311),
.B(n_292),
.C(n_275),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_590),
.B(n_231),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_535),
.B(n_262),
.Y(n_722)
);

AO22x1_ASAP7_75t_L g723 ( 
.A1(n_596),
.A2(n_211),
.B1(n_218),
.B2(n_238),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_590),
.B(n_267),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_622),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_615),
.Y(n_726)
);

OAI221xp5_ASAP7_75t_L g727 ( 
.A1(n_515),
.A2(n_634),
.B1(n_626),
.B2(n_641),
.C(n_579),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_597),
.B(n_267),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_519),
.A2(n_292),
.B1(n_311),
.B2(n_273),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_519),
.A2(n_337),
.B1(n_333),
.B2(n_345),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_615),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_597),
.B(n_273),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_601),
.B(n_275),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_SL g734 ( 
.A(n_567),
.B(n_480),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_582),
.B(n_437),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_548),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_625),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_630),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_576),
.A2(n_304),
.B(n_290),
.C(n_326),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_611),
.B(n_245),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_625),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_608),
.B(n_317),
.Y(n_742)
);

OAI221xp5_ASAP7_75t_L g743 ( 
.A1(n_638),
.A2(n_326),
.B1(n_344),
.B2(n_341),
.C(n_322),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_553),
.A2(n_317),
.B(n_339),
.C(n_340),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_635),
.B(n_264),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_643),
.A2(n_335),
.B1(n_322),
.B2(n_344),
.C(n_341),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_266),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_571),
.B(n_274),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_281),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_606),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_530),
.B(n_347),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_636),
.B(n_347),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_619),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_629),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_530),
.B(n_245),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_613),
.A2(n_334),
.B1(n_248),
.B2(n_268),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_546),
.B(n_245),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_557),
.A2(n_328),
.B1(n_268),
.B2(n_289),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_629),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_576),
.A2(n_328),
.B(n_334),
.C(n_289),
.Y(n_762)
);

OAI22x1_ASAP7_75t_SL g763 ( 
.A1(n_618),
.A2(n_329),
.B1(n_307),
.B2(n_310),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_567),
.B(n_472),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_606),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_578),
.A2(n_245),
.B1(n_300),
.B2(n_468),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_546),
.B(n_300),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_560),
.B(n_575),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_562),
.B(n_342),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_521),
.B(n_324),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_551),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_533),
.B(n_314),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_603),
.B(n_300),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_625),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_567),
.B(n_472),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_533),
.B(n_428),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_546),
.B(n_300),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_556),
.A2(n_423),
.B(n_422),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_551),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_556),
.A2(n_422),
.B(n_468),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_580),
.A2(n_516),
.B1(n_554),
.B2(n_564),
.Y(n_781)
);

AO22x1_ASAP7_75t_L g782 ( 
.A1(n_554),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_675),
.A2(n_580),
.B1(n_554),
.B2(n_592),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_663),
.A2(n_514),
.B(n_517),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_727),
.A2(n_517),
.B(n_557),
.C(n_554),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_768),
.B(n_552),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_768),
.B(n_593),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_681),
.A2(n_552),
.B(n_591),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_668),
.A2(n_552),
.B(n_558),
.C(n_588),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_668),
.A2(n_617),
.B1(n_632),
.B2(n_538),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_657),
.A2(n_591),
.B(n_605),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_675),
.B(n_670),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_705),
.A2(n_621),
.B(n_633),
.C(n_624),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_657),
.A2(n_565),
.B(n_605),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_670),
.B(n_545),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_705),
.A2(n_568),
.B(n_581),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_781),
.B(n_545),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_754),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_689),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_689),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_755),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_689),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_752),
.A2(n_632),
.B1(n_577),
.B2(n_561),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_756),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_761),
.Y(n_806)
);

INVx6_ASAP7_75t_L g807 ( 
.A(n_737),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_682),
.B(n_709),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_750),
.B(n_567),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_713),
.A2(n_516),
.B(n_644),
.C(n_640),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_680),
.A2(n_598),
.B1(n_516),
.B2(n_632),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_693),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_713),
.A2(n_617),
.B1(n_632),
.B2(n_538),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_666),
.B(n_549),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_650),
.B(n_522),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_646),
.A2(n_637),
.B(n_550),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_650),
.B(n_522),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_647),
.A2(n_637),
.B(n_550),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_729),
.A2(n_639),
.B(n_631),
.C(n_617),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_669),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_693),
.B(n_542),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_703),
.B(n_631),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_710),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_747),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_L g825 ( 
.A1(n_680),
.A2(n_449),
.B(n_470),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_685),
.B(n_550),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_698),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_716),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_685),
.B(n_599),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_651),
.B(n_599),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_676),
.B(n_674),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_750),
.B(n_542),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_751),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_736),
.B(n_449),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_672),
.A2(n_537),
.B(n_584),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_673),
.A2(n_537),
.B(n_584),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_652),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_737),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_664),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_662),
.A2(n_534),
.B(n_528),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_686),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_752),
.A2(n_534),
.B(n_528),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_691),
.A2(n_671),
.B(n_663),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_769),
.A2(n_628),
.B1(n_574),
.B2(n_531),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_671),
.A2(n_692),
.B(n_688),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_688),
.A2(n_574),
.B(n_531),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_749),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_694),
.B(n_628),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_757),
.A2(n_581),
.B(n_568),
.C(n_609),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_760),
.B(n_642),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_695),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_760),
.A2(n_628),
.B(n_586),
.C(n_609),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_776),
.A2(n_572),
.B(n_570),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_696),
.B(n_583),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_649),
.B(n_642),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_715),
.B(n_726),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_731),
.B(n_583),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_738),
.B(n_595),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_648),
.B(n_470),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_735),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_748),
.B(n_602),
.C(n_620),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_737),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_R g863 ( 
.A(n_725),
.B(n_136),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_687),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_764),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_741),
.Y(n_867)
);

NOR2x1p5_ASAP7_75t_SL g868 ( 
.A(n_645),
.B(n_620),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_702),
.A2(n_12),
.B(n_14),
.C(n_16),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_741),
.B(n_538),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_701),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_749),
.B(n_17),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_690),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_656),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_770),
.A2(n_536),
.B(n_620),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_772),
.A2(n_679),
.B(n_706),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_654),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_780),
.B(n_160),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_719),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_679),
.A2(n_536),
.B(n_620),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_536),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_704),
.B(n_17),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_774),
.B(n_620),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_655),
.A2(n_137),
.B(n_121),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_720),
.A2(n_744),
.B(n_767),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_660),
.A2(n_112),
.B(n_100),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_661),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_SL g889 ( 
.A1(n_759),
.A2(n_21),
.B(n_22),
.C(n_24),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_659),
.A2(n_84),
.B(n_82),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_667),
.B(n_81),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_699),
.B(n_21),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_677),
.A2(n_758),
.B1(n_777),
.B2(n_767),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_656),
.B(n_22),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_777),
.A2(n_70),
.B(n_25),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_722),
.B(n_24),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_711),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_717),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_712),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_SL g900 ( 
.A(n_700),
.B(n_734),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_708),
.B(n_26),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_684),
.B(n_29),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_678),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_697),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_656),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_717),
.B(n_41),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_771),
.A2(n_41),
.B(n_42),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_779),
.A2(n_43),
.B(n_44),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_745),
.B(n_43),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_721),
.A2(n_48),
.B(n_49),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_707),
.B(n_50),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_L g912 ( 
.A(n_745),
.B(n_52),
.C(n_54),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_714),
.A2(n_55),
.B(n_56),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_730),
.A2(n_55),
.B(n_57),
.C(n_60),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_718),
.A2(n_57),
.B(n_64),
.C(n_68),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_724),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_683),
.B(n_68),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_690),
.A2(n_69),
.B(n_753),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_728),
.B(n_69),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_683),
.B(n_775),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_739),
.A2(n_762),
.B(n_740),
.C(n_733),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_732),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_742),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_690),
.A2(n_778),
.B(n_773),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_658),
.A2(n_665),
.B(n_723),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_758),
.A2(n_746),
.B(n_743),
.C(n_683),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_766),
.B(n_782),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_797),
.A2(n_653),
.B(n_763),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_786),
.B(n_923),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_899),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_798),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_797),
.A2(n_784),
.B(n_855),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_809),
.B(n_787),
.Y(n_934)
);

OA22x2_ASAP7_75t_L g935 ( 
.A1(n_847),
.A2(n_911),
.B1(n_903),
.B2(n_927),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_812),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_899),
.Y(n_937)
);

AO31x2_ASAP7_75t_L g938 ( 
.A1(n_789),
.A2(n_906),
.A3(n_810),
.B(n_921),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_798),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_880),
.B(n_875),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_798),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_911),
.A2(n_873),
.B1(n_909),
.B2(n_893),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_785),
.A2(n_789),
.B(n_845),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_905),
.B(n_834),
.Y(n_944)
);

NAND2x1_ASAP7_75t_L g945 ( 
.A(n_801),
.B(n_807),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_860),
.Y(n_946)
);

AO31x2_ASAP7_75t_L g947 ( 
.A1(n_810),
.A2(n_852),
.A3(n_915),
.B(n_804),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_863),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_840),
.A2(n_836),
.B(n_835),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_863),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_783),
.A2(n_831),
.B(n_847),
.C(n_814),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_798),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_831),
.B(n_900),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_814),
.A2(n_925),
.B(n_893),
.C(n_811),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_837),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_850),
.A2(n_795),
.B1(n_790),
.B2(n_813),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_916),
.B(n_922),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_799),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_821),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_827),
.B(n_822),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_822),
.B(n_839),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_841),
.B(n_851),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_853),
.A2(n_876),
.B(n_842),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_874),
.B(n_832),
.Y(n_964)
);

OAI21xp33_ASAP7_75t_L g965 ( 
.A1(n_856),
.A2(n_825),
.B(n_896),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_926),
.A2(n_895),
.B(n_793),
.C(n_886),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_838),
.Y(n_967)
);

AO31x2_ASAP7_75t_L g968 ( 
.A1(n_852),
.A2(n_915),
.A3(n_829),
.B(n_826),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_878),
.B(n_888),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_874),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_833),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_864),
.B(n_823),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_823),
.B(n_828),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_816),
.A2(n_818),
.B(n_796),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_866),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_788),
.A2(n_879),
.B(n_904),
.C(n_913),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_874),
.B(n_801),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_828),
.B(n_808),
.Y(n_978)
);

AND2x6_ASAP7_75t_L g979 ( 
.A(n_838),
.B(n_867),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_815),
.B(n_817),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_874),
.B(n_838),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_912),
.B(n_914),
.C(n_919),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_SL g983 ( 
.A1(n_819),
.A2(n_872),
.B(n_867),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_850),
.A2(n_882),
.B(n_884),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_830),
.B(n_848),
.Y(n_985)
);

NAND2x1_ASAP7_75t_L g986 ( 
.A(n_807),
.B(n_872),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_920),
.B(n_894),
.Y(n_987)
);

NAND2x1_ASAP7_75t_L g988 ( 
.A(n_807),
.B(n_867),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_SL g989 ( 
.A1(n_914),
.A2(n_917),
.B(n_898),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_881),
.A2(n_849),
.B(n_870),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_790),
.A2(n_918),
.B(n_924),
.C(n_861),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_813),
.A2(n_861),
.B(n_844),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_802),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_902),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_859),
.Y(n_995)
);

AO31x2_ASAP7_75t_L g996 ( 
.A1(n_869),
.A2(n_892),
.A3(n_901),
.B(n_908),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_854),
.B(n_857),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_808),
.B(n_805),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_858),
.B(n_806),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_800),
.A2(n_803),
.B(n_862),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_820),
.A2(n_865),
.B1(n_897),
.B2(n_871),
.Y(n_1001)
);

AO31x2_ASAP7_75t_L g1002 ( 
.A1(n_869),
.A2(n_887),
.A3(n_885),
.B(n_890),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_872),
.B(n_907),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_868),
.B(n_891),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_889),
.A2(n_910),
.B(n_883),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_SL g1006 ( 
.A1(n_889),
.A2(n_792),
.B(n_786),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_792),
.B(n_786),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_812),
.B(n_520),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_792),
.B(n_786),
.Y(n_1009)
);

AO31x2_ASAP7_75t_L g1010 ( 
.A1(n_789),
.A2(n_906),
.A3(n_720),
.B(n_729),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_874),
.B(n_657),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_809),
.B(n_479),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_791),
.A2(n_657),
.B(n_794),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_792),
.B(n_786),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_792),
.A2(n_906),
.B(n_787),
.C(n_675),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_899),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_798),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_877),
.A2(n_846),
.B(n_843),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_789),
.A2(n_906),
.A3(n_720),
.B(n_729),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_791),
.A2(n_657),
.B(n_794),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_809),
.B(n_479),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_798),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_792),
.B(n_786),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_787),
.A2(n_768),
.B1(n_906),
.B2(n_792),
.Y(n_1024)
);

OAI22x1_ASAP7_75t_L g1025 ( 
.A1(n_787),
.A2(n_766),
.B1(n_768),
.B2(n_906),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_877),
.A2(n_846),
.B(n_843),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_792),
.B(n_786),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_877),
.A2(n_846),
.B(n_843),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_906),
.B(n_787),
.C(n_685),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_785),
.A2(n_789),
.B(n_792),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_877),
.A2(n_846),
.B(n_843),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_SL g1032 ( 
.A1(n_895),
.A2(n_785),
.B(n_886),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_792),
.B(n_786),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_809),
.B(n_479),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_792),
.B(n_786),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_785),
.A2(n_789),
.B(n_792),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_785),
.A2(n_789),
.B(n_792),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_792),
.B(n_786),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_812),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_787),
.B(n_847),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_792),
.A2(n_670),
.B1(n_668),
.B2(n_713),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_812),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_812),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_792),
.B(n_786),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_809),
.B(n_479),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_809),
.B(n_479),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_792),
.B(n_786),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_785),
.A2(n_789),
.B(n_792),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_792),
.A2(n_906),
.B(n_787),
.C(n_675),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_824),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_789),
.A2(n_906),
.A3(n_720),
.B(n_729),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_877),
.A2(n_846),
.B(n_843),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_791),
.A2(n_657),
.B(n_794),
.Y(n_1053)
);

AND2x6_ASAP7_75t_L g1054 ( 
.A(n_811),
.B(n_792),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_798),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_SL g1056 ( 
.A1(n_792),
.A2(n_906),
.B1(n_729),
.B2(n_668),
.C(n_670),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_880),
.B(n_690),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_789),
.A2(n_906),
.A3(n_720),
.B(n_729),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_787),
.B(n_768),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_931),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1042),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_1043),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_971),
.Y(n_1064)
);

OR2x6_ASAP7_75t_L g1065 ( 
.A(n_1057),
.B(n_944),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_934),
.B(n_1029),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1025),
.A2(n_953),
.B1(n_995),
.B2(n_965),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_929),
.B(n_960),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_929),
.B(n_969),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_1057),
.B(n_944),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_971),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_936),
.Y(n_1073)
);

CKINVDCx6p67_ASAP7_75t_R g1074 ( 
.A(n_946),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_954),
.A2(n_951),
.B(n_942),
.C(n_982),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_966),
.B(n_989),
.C(n_1041),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1034),
.B(n_1045),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_939),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_956),
.A2(n_1041),
.A3(n_1006),
.B1(n_935),
.B2(n_1037),
.Y(n_1080)
);

AOI222xp33_ASAP7_75t_L g1081 ( 
.A1(n_1040),
.A2(n_956),
.B1(n_989),
.B2(n_1046),
.C1(n_961),
.C2(n_959),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_970),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_979),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_944),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_987),
.A2(n_935),
.B1(n_1054),
.B2(n_978),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1050),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_959),
.B(n_1008),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1039),
.B(n_972),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_975),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_940),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1007),
.B(n_1009),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_L g1092 ( 
.A(n_948),
.B(n_950),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_994),
.B(n_957),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_940),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_979),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_958),
.B(n_993),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_962),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_940),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_964),
.B(n_1057),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_998),
.A2(n_973),
.B(n_999),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_930),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_991),
.A2(n_976),
.B(n_980),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_939),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_SL g1107 ( 
.A1(n_1030),
.A2(n_1036),
.B(n_1037),
.C(n_1048),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_964),
.B(n_928),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_939),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_937),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_979),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_952),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1054),
.A2(n_1056),
.B1(n_1033),
.B2(n_1035),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_980),
.A2(n_983),
.B(n_1027),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1016),
.B(n_970),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_999),
.B(n_1027),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_945),
.B(n_952),
.Y(n_1117)
);

INVx8_ASAP7_75t_L g1118 ( 
.A(n_979),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1033),
.B(n_1035),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1054),
.A2(n_1032),
.B1(n_992),
.B2(n_1036),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1001),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_952),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_1005),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_932),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_981),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_943),
.A2(n_992),
.B(n_1047),
.C(n_984),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1017),
.Y(n_1128)
);

NAND2x1p5_ASAP7_75t_L g1129 ( 
.A(n_1017),
.B(n_1055),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_1004),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_932),
.B(n_941),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_981),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_986),
.A2(n_988),
.B1(n_967),
.B2(n_977),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_997),
.B(n_1004),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1017),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_1055),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1022),
.B(n_996),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1013),
.A2(n_1020),
.B(n_1053),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1003),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1055),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_985),
.B(n_933),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_SL g1142 ( 
.A(n_1011),
.B(n_977),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1000),
.B(n_938),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_990),
.A2(n_974),
.B(n_949),
.C(n_1052),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1011),
.B(n_938),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_996),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1018),
.A2(n_1026),
.B(n_1031),
.C(n_1028),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_968),
.B(n_947),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_947),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_947),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_968),
.B(n_1058),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_968),
.B(n_1010),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1010),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1002),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_963),
.B(n_1010),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_1002),
.A2(n_1019),
.B(n_1051),
.C(n_1058),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_931),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1059),
.B(n_520),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_971),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_931),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1024),
.A2(n_906),
.B(n_792),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_964),
.B(n_1057),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1029),
.A2(n_787),
.B1(n_768),
.B2(n_700),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1059),
.A2(n_1024),
.B1(n_668),
.B2(n_670),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1059),
.B(n_520),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1029),
.A2(n_1049),
.B(n_1015),
.C(n_1024),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_971),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_939),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_964),
.B(n_1057),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1042),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_931),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_939),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1043),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_931),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_943),
.A2(n_1036),
.B(n_1030),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_1039),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_931),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1057),
.B(n_944),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_939),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1059),
.B(n_1024),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1029),
.B(n_787),
.C(n_768),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_931),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_939),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_971),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_939),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1086),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1067),
.B(n_1158),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1112),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1072),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1167),
.A2(n_1192),
.B1(n_1070),
.B2(n_1069),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1149),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1083),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1163),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1064),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1083),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1087),
.A2(n_1100),
.B1(n_1187),
.B2(n_1171),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1064),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1118),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1070),
.B(n_1066),
.Y(n_1212)
);

AO21x2_ASAP7_75t_L g1213 ( 
.A1(n_1147),
.A2(n_1138),
.B(n_1144),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1168),
.A2(n_1180),
.B1(n_1186),
.B2(n_1178),
.Y(n_1214)
);

BUFx4f_ASAP7_75t_SL g1215 ( 
.A(n_1073),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1137),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1172),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1105),
.A2(n_1114),
.B(n_1170),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1078),
.B(n_1157),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1068),
.A2(n_1182),
.B1(n_1160),
.B2(n_1195),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1108),
.A2(n_1159),
.B1(n_1180),
.B2(n_1178),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1222)
);

CKINVDCx6p67_ASAP7_75t_R g1223 ( 
.A(n_1135),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1081),
.A2(n_1120),
.B1(n_1165),
.B2(n_1191),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1077),
.A2(n_1148),
.B(n_1146),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1116),
.B(n_1130),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1118),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_SL g1228 ( 
.A1(n_1148),
.A2(n_1085),
.B(n_1153),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1083),
.B(n_1096),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_1127),
.A2(n_1107),
.B(n_1156),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1184),
.A2(n_1084),
.B1(n_1099),
.B2(n_1069),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1151),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1172),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1080),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1162),
.B(n_1169),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1083),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1074),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1176),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1061),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1096),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1081),
.A2(n_1089),
.B1(n_1103),
.B2(n_1175),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1196),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1096),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1076),
.A2(n_1088),
.B1(n_1134),
.B2(n_1196),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1080),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1062),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1177),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1183),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1094),
.B(n_1185),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1188),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1060),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1184),
.A2(n_1095),
.B1(n_1090),
.B2(n_1145),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1155),
.A2(n_1143),
.B(n_1152),
.Y(n_1254)
);

BUFx4f_ASAP7_75t_SL g1255 ( 
.A(n_1174),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_1122),
.B1(n_1121),
.B2(n_1075),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1155),
.A2(n_1143),
.B(n_1119),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1145),
.A2(n_1098),
.B1(n_1102),
.B2(n_1075),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1093),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1091),
.B(n_1102),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1161),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1101),
.A2(n_1166),
.B1(n_1175),
.B2(n_1065),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1080),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1091),
.B(n_1119),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1098),
.B(n_1121),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1124),
.A2(n_1141),
.B(n_1113),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1139),
.A2(n_1082),
.B(n_1117),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1096),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1104),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1082),
.A2(n_1117),
.B(n_1125),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1111),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1097),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1164),
.B(n_1193),
.Y(n_1273)
);

INVx6_ASAP7_75t_L g1274 ( 
.A(n_1111),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1065),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1111),
.A2(n_1166),
.B1(n_1101),
.B2(n_1065),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVx5_ASAP7_75t_L g1278 ( 
.A(n_1111),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_SL g1279 ( 
.A(n_1123),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1110),
.A2(n_1115),
.B(n_1142),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1071),
.A2(n_1189),
.B1(n_1118),
.B2(n_1142),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1071),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1140),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1131),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1131),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1129),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1136),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1092),
.B(n_1071),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1106),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1106),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1079),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1189),
.A2(n_1132),
.B1(n_1126),
.B2(n_1133),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1189),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1126),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1132),
.A2(n_1079),
.B(n_1109),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1173),
.A2(n_1197),
.B1(n_1109),
.B2(n_1179),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1173),
.A2(n_1197),
.B(n_1109),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1079),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1194),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1179),
.A2(n_734),
.B1(n_787),
.B2(n_768),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1190),
.A2(n_1029),
.B1(n_787),
.B2(n_906),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1190),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1194),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1194),
.B(n_1067),
.Y(n_1304)
);

INVx8_ASAP7_75t_L g1305 ( 
.A(n_1118),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1072),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1072),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1072),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1167),
.A2(n_1059),
.B1(n_1024),
.B2(n_1029),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1067),
.B(n_1158),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1067),
.B(n_1158),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1150),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1088),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1150),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1072),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1072),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1112),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1167),
.A2(n_1059),
.B1(n_1024),
.B2(n_1029),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1067),
.B(n_1158),
.Y(n_1319)
);

AO21x1_ASAP7_75t_L g1320 ( 
.A1(n_1063),
.A2(n_956),
.B(n_906),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1083),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1201),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1266),
.B(n_1257),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1217),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1233),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1318),
.A2(n_1309),
.B1(n_1224),
.B2(n_1202),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1254),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1216),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1201),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1266),
.B(n_1257),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1312),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1295),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1216),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1275),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1314),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1308),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1199),
.B(n_1310),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1254),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1199),
.B(n_1310),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1236),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1308),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1311),
.B(n_1319),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1203),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1232),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1311),
.A2(n_1319),
.B1(n_1320),
.B2(n_1214),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1210),
.B(n_1225),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1225),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1225),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1234),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1210),
.B(n_1264),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1264),
.B(n_1265),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1245),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1265),
.B(n_1304),
.Y(n_1353)
);

INVxp33_ASAP7_75t_L g1354 ( 
.A(n_1250),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1226),
.B(n_1263),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1263),
.B(n_1230),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1239),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1221),
.B(n_1222),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1269),
.Y(n_1359)
);

XNOR2xp5_ASAP7_75t_L g1360 ( 
.A(n_1208),
.B(n_1239),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1278),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1275),
.B(n_1282),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.B(n_1230),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1213),
.A2(n_1230),
.B(n_1228),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1315),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1228),
.A2(n_1256),
.B(n_1301),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1218),
.B(n_1273),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1270),
.A2(n_1267),
.B(n_1229),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1300),
.A2(n_1241),
.B(n_1220),
.Y(n_1369)
);

INVxp33_ASAP7_75t_L g1370 ( 
.A(n_1219),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1218),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1282),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1260),
.B(n_1212),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1218),
.B(n_1273),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1235),
.B(n_1272),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1293),
.B(n_1280),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1293),
.B(n_1229),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1315),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1316),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1316),
.B(n_1205),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1206),
.B(n_1209),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1252),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1259),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1258),
.A2(n_1231),
.B(n_1270),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1261),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1278),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1267),
.A2(n_1229),
.B(n_1243),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1305),
.B(n_1274),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1278),
.B(n_1271),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1238),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1246),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1305),
.B(n_1274),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1242),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1285),
.B(n_1198),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1295),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1247),
.Y(n_1397)
);

NAND2x1_ASAP7_75t_L g1398 ( 
.A(n_1204),
.B(n_1274),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1248),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1346),
.B(n_1253),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1322),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1354),
.B(n_1200),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1326),
.A2(n_1313),
.B1(n_1281),
.B2(n_1317),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1346),
.B(n_1251),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1368),
.B(n_1367),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1329),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1374),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1389),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1336),
.Y(n_1409)
);

NOR4xp25_ASAP7_75t_SL g1410 ( 
.A(n_1396),
.B(n_1302),
.C(n_1283),
.D(n_1286),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1374),
.B(n_1289),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1331),
.B(n_1268),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1350),
.B(n_1313),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1358),
.B(n_1290),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1350),
.B(n_1313),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1363),
.B(n_1288),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1398),
.Y(n_1418)
);

OAI222xp33_ASAP7_75t_L g1419 ( 
.A1(n_1345),
.A2(n_1276),
.B1(n_1262),
.B2(n_1292),
.C1(n_1294),
.C2(n_1284),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1337),
.B(n_1295),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1387),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1341),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1338),
.Y(n_1423)
);

AOI211xp5_ASAP7_75t_L g1424 ( 
.A1(n_1369),
.A2(n_1249),
.B(n_1317),
.C(n_1200),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_SL g1425 ( 
.A(n_1323),
.B(n_1321),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1358),
.B(n_1277),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1339),
.B(n_1295),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1339),
.B(n_1294),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1335),
.B(n_1243),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1365),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1398),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1360),
.A2(n_1223),
.B1(n_1274),
.B2(n_1204),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1387),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1342),
.B(n_1271),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_1287),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1357),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1327),
.B(n_1271),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1356),
.B(n_1303),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_1351),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1351),
.B(n_1353),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1353),
.B(n_1240),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1355),
.B(n_1240),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1344),
.B(n_1240),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1383),
.B(n_1243),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1356),
.B(n_1207),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1370),
.A2(n_1223),
.B1(n_1238),
.B2(n_1237),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1378),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1347),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1426),
.B(n_1359),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1426),
.B(n_1380),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1424),
.B(n_1384),
.C(n_1373),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1424),
.B(n_1392),
.C(n_1325),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1403),
.B(n_1417),
.C(n_1435),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1417),
.A2(n_1376),
.B1(n_1362),
.B2(n_1366),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1407),
.B(n_1332),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1407),
.B(n_1332),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1432),
.B(n_1376),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1414),
.B(n_1380),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1419),
.A2(n_1360),
.B(n_1376),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1435),
.B(n_1414),
.C(n_1402),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1401),
.B(n_1324),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1407),
.B(n_1364),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1409),
.B(n_1388),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1420),
.B(n_1364),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1422),
.B(n_1388),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1447),
.B(n_1379),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1394),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1432),
.A2(n_1376),
.B1(n_1362),
.B2(n_1366),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1446),
.A2(n_1375),
.B1(n_1389),
.B2(n_1393),
.Y(n_1469)
);

NAND4xp25_ASAP7_75t_SL g1470 ( 
.A(n_1400),
.B(n_1381),
.C(n_1296),
.D(n_1382),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1418),
.B(n_1362),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1427),
.B(n_1364),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1427),
.B(n_1327),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1406),
.A2(n_1389),
.B1(n_1393),
.B2(n_1377),
.Y(n_1474)
);

AOI21xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1400),
.A2(n_1366),
.B(n_1323),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1430),
.B(n_1366),
.C(n_1372),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1415),
.Y(n_1478)
);

OAI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1430),
.A2(n_1323),
.B(n_1330),
.Y(n_1479)
);

NAND4xp25_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1372),
.C(n_1385),
.D(n_1382),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1418),
.A2(n_1330),
.B1(n_1323),
.B2(n_1377),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1413),
.A2(n_1362),
.B1(n_1323),
.B2(n_1330),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1405),
.B(n_1327),
.Y(n_1484)
);

NAND3xp33_ASAP7_75t_L g1485 ( 
.A(n_1410),
.B(n_1399),
.C(n_1397),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1405),
.B(n_1348),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1405),
.B(n_1348),
.Y(n_1487)
);

NOR3xp33_ASAP7_75t_L g1488 ( 
.A(n_1419),
.B(n_1386),
.C(n_1361),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1434),
.B(n_1328),
.Y(n_1489)
);

OAI21xp33_ASAP7_75t_L g1490 ( 
.A1(n_1434),
.A2(n_1330),
.B(n_1428),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1410),
.B(n_1395),
.C(n_1330),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1328),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1437),
.A2(n_1390),
.B(n_1395),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1411),
.A2(n_1377),
.B1(n_1237),
.B2(n_1333),
.C(n_1389),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1439),
.B(n_1333),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1416),
.B(n_1411),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1443),
.B(n_1399),
.C(n_1397),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1438),
.B(n_1348),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1436),
.A2(n_1389),
.B1(n_1393),
.B2(n_1377),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1438),
.B(n_1349),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1416),
.B(n_1349),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1442),
.B(n_1352),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1444),
.B(n_1334),
.C(n_1343),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_L g1505 ( 
.A(n_1444),
.B(n_1385),
.C(n_1383),
.D(n_1343),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1404),
.B(n_1334),
.C(n_1371),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1442),
.B(n_1352),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1391),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1478),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1478),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1484),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1499),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1484),
.Y(n_1513)
);

AND2x4_ASAP7_75t_SL g1514 ( 
.A(n_1488),
.B(n_1408),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_1404),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_1476),
.B(n_1421),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1463),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1493),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1458),
.B(n_1449),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1486),
.B(n_1425),
.Y(n_1521)
);

NAND2x1_ASAP7_75t_L g1522 ( 
.A(n_1498),
.B(n_1408),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1486),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1450),
.B(n_1418),
.Y(n_1524)
);

NAND2x1_ASAP7_75t_SL g1525 ( 
.A(n_1462),
.B(n_1421),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1464),
.B(n_1448),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1499),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1423),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1487),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1465),
.B(n_1431),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1467),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1487),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1455),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1457),
.B(n_1408),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1462),
.B(n_1425),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1464),
.B(n_1448),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1461),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1500),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1473),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1489),
.B(n_1441),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1481),
.B(n_1423),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1456),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1472),
.B(n_1497),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1448),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_1441),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1515),
.B(n_1503),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1546),
.B(n_1466),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1509),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1516),
.B(n_1451),
.C(n_1452),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1529),
.B(n_1475),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1520),
.B(n_1503),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1531),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1531),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1517),
.B(n_1518),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1475),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1563)
);

NAND4xp75_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1471),
.C(n_1483),
.D(n_1437),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1543),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1507),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1532),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1543),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1512),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_SL g1570 ( 
.A(n_1539),
.B(n_1452),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1523),
.Y(n_1571)
);

NAND4xp75_ASAP7_75t_L g1572 ( 
.A(n_1508),
.B(n_1483),
.C(n_1459),
.D(n_1227),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1453),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1538),
.B(n_1502),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1523),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1512),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1527),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1523),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1520),
.B(n_1502),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1522),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1526),
.B(n_1480),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1520),
.B(n_1490),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1520),
.B(n_1454),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1526),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1537),
.B(n_1485),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1525),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1537),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1551),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1570),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1561),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1570),
.A2(n_1553),
.B1(n_1572),
.B2(n_1539),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1552),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1577),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1573),
.B(n_1522),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1551),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1542),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1584),
.B(n_1536),
.Y(n_1601)
);

AND2x4_ASAP7_75t_SL g1602 ( 
.A(n_1584),
.B(n_1580),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1556),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1587),
.B(n_1542),
.Y(n_1609)
);

INVx3_ASAP7_75t_SL g1610 ( 
.A(n_1588),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1553),
.B(n_1534),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1587),
.B(n_1527),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1552),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1561),
.B(n_1534),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1582),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1552),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1549),
.B(n_1534),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1564),
.B(n_1470),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1572),
.A2(n_1479),
.B1(n_1514),
.B2(n_1535),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1577),
.B(n_1548),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1559),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1549),
.B(n_1535),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1583),
.Y(n_1625)
);

CKINVDCx16_ASAP7_75t_R g1626 ( 
.A(n_1585),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1566),
.B(n_1541),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1581),
.B(n_1536),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1582),
.B(n_1521),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1566),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1585),
.A2(n_1469),
.B(n_1535),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1550),
.B(n_1540),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1618),
.A2(n_1479),
.B1(n_1514),
.B2(n_1468),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1626),
.B(n_1555),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1588),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1590),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1592),
.B(n_1574),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1593),
.A2(n_1514),
.B1(n_1408),
.B2(n_1555),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1555),
.Y(n_1639)
);

AOI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1623),
.A2(n_1562),
.B1(n_1574),
.B2(n_1589),
.C1(n_1586),
.C2(n_1504),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.B(n_1562),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1600),
.B(n_1621),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1602),
.B(n_1588),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1586),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1601),
.B(n_1562),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1610),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1595),
.B(n_1597),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1586),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1615),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1610),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1629),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1598),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1611),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1215),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1630),
.B(n_1624),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1624),
.B(n_1550),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1604),
.B(n_1589),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1627),
.B(n_1557),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1599),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1603),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1631),
.A2(n_1482),
.B1(n_1474),
.B2(n_1431),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1620),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1605),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1606),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1622),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1557),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1650),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1662),
.A2(n_1596),
.B(n_1614),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1607),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1612),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1653),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1664),
.A2(n_1633),
.B1(n_1663),
.B2(n_1638),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1653),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1628),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1628),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1652),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1660),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1656),
.A2(n_1609),
.B1(n_1613),
.B2(n_1612),
.C(n_1617),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1639),
.B(n_1609),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1634),
.B(n_1589),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1661),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.B(n_1632),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1640),
.A2(n_1632),
.B1(n_1494),
.B2(n_1525),
.C(n_1616),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1652),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1655),
.B(n_1255),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1634),
.B(n_1559),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1560),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1635),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1687),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1694),
.B(n_1635),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1676),
.A2(n_1637),
.B1(n_1666),
.B2(n_1665),
.C(n_1667),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1683),
.B(n_1643),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1680),
.B(n_1649),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1674),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1675),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1677),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1670),
.B(n_1672),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1684),
.B(n_1635),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1689),
.B(n_1644),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1681),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1659),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1691),
.B(n_1657),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1644),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1684),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1678),
.B(n_1644),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1696),
.B(n_1692),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1698),
.A2(n_1688),
.B(n_1671),
.Y(n_1716)
);

OAI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1712),
.A2(n_1682),
.B(n_1686),
.C(n_1690),
.Y(n_1717)
);

AOI222xp33_ASAP7_75t_L g1718 ( 
.A1(n_1695),
.A2(n_1705),
.B1(n_1699),
.B2(n_1702),
.C1(n_1710),
.C2(n_1713),
.Y(n_1718)
);

AOI222xp33_ASAP7_75t_L g1719 ( 
.A1(n_1705),
.A2(n_1692),
.B1(n_1673),
.B2(n_1693),
.C1(n_1649),
.C2(n_1665),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1699),
.A2(n_1666),
.B(n_1636),
.Y(n_1720)
);

O2A1O1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1701),
.A2(n_1693),
.B(n_1691),
.C(n_1645),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1700),
.A2(n_1645),
.B1(n_1642),
.B2(n_1646),
.C(n_1668),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1710),
.A2(n_1649),
.B(n_1658),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1707),
.A2(n_1646),
.B1(n_1642),
.B2(n_1594),
.C(n_1616),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1697),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1697),
.A2(n_1658),
.B(n_1594),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1707),
.A2(n_1619),
.B1(n_1431),
.B2(n_1569),
.C(n_1576),
.Y(n_1727)
);

OA22x2_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1697),
.B1(n_1696),
.B2(n_1706),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1721),
.B(n_1696),
.C(n_1703),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1725),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1715),
.B(n_1714),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1720),
.B(n_1704),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1723),
.B(n_1708),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1718),
.B(n_1709),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1719),
.B(n_1722),
.C(n_1717),
.D(n_1724),
.Y(n_1735)
);

XNOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1727),
.B(n_1711),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1720),
.B(n_1726),
.Y(n_1737)
);

NAND4xp25_ASAP7_75t_L g1738 ( 
.A(n_1718),
.B(n_1658),
.C(n_1619),
.D(n_1491),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1718),
.B(n_1485),
.C(n_1298),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1716),
.A2(n_1580),
.B(n_1558),
.C(n_1576),
.Y(n_1740)
);

NOR3xp33_ASAP7_75t_L g1741 ( 
.A(n_1734),
.B(n_1735),
.C(n_1730),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_SL g1742 ( 
.A(n_1740),
.B(n_1279),
.C(n_1506),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1731),
.B(n_1571),
.Y(n_1743)
);

NAND4xp25_ASAP7_75t_L g1744 ( 
.A(n_1729),
.B(n_1521),
.C(n_1558),
.D(n_1498),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1738),
.A2(n_1482),
.B1(n_1565),
.B2(n_1568),
.C(n_1560),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1737),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1733),
.B(n_1521),
.C(n_1563),
.D(n_1578),
.Y(n_1747)
);

OAI22x1_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1732),
.B1(n_1736),
.B2(n_1739),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1741),
.A2(n_1728),
.B1(n_1521),
.B2(n_1579),
.Y(n_1749)
);

NOR2x1_ASAP7_75t_L g1750 ( 
.A(n_1747),
.B(n_1571),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1579),
.B1(n_1575),
.B2(n_1568),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1743),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1742),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1745),
.A2(n_1579),
.B1(n_1575),
.B2(n_1565),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1748),
.A2(n_1227),
.B(n_1211),
.Y(n_1755)
);

NAND2x1_ASAP7_75t_L g1756 ( 
.A(n_1750),
.B(n_1575),
.Y(n_1756)
);

NAND4xp75_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1211),
.C(n_1578),
.D(n_1569),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1749),
.Y(n_1758)
);

NOR2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1759)
);

AND3x4_ASAP7_75t_L g1760 ( 
.A(n_1751),
.B(n_1429),
.C(n_1412),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1759),
.Y(n_1761)
);

XNOR2xp5_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1757),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1755),
.Y(n_1763)
);

XOR2x2_ASAP7_75t_L g1764 ( 
.A(n_1762),
.B(n_1760),
.Y(n_1764)
);

AOI222xp33_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1761),
.B1(n_1763),
.B2(n_1756),
.C1(n_1563),
.C2(n_1545),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1511),
.B1(n_1513),
.B2(n_1545),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1765),
.A2(n_1563),
.B(n_1297),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1513),
.B1(n_1511),
.B2(n_1533),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1767),
.A2(n_1297),
.B(n_1291),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_1299),
.B1(n_1302),
.B2(n_1421),
.Y(n_1770)
);

AOI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1544),
.B(n_1528),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1770),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1771),
.B1(n_1421),
.B2(n_1433),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1544),
.B1(n_1528),
.B2(n_1533),
.C(n_1236),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1236),
.B(n_1321),
.C(n_1340),
.Y(n_1775)
);


endmodule