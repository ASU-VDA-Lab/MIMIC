module fake_jpeg_26425_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_47),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_0),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_52),
.B1(n_63),
.B2(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_19),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_20),
.B1(n_28),
.B2(n_32),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_59),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_28),
.B1(n_33),
.B2(n_21),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_35),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_29),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_74),
.B(n_80),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_83),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_46),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_58),
.B(n_6),
.C(n_5),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_49),
.C(n_67),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_50),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_82),
.B(n_85),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_9),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_1),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_8),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_12),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_117),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_112),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_76),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_81),
.Y(n_127)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_95),
.B1(n_86),
.B2(n_90),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_99),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_99),
.B(n_72),
.C(n_87),
.D(n_79),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_149),
.B1(n_106),
.B2(n_104),
.C(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_99),
.C(n_91),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_58),
.B1(n_84),
.B2(n_96),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_107),
.B1(n_104),
.B2(n_93),
.Y(n_161)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_152),
.Y(n_172)
);

XOR2x2_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_112),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_117),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_105),
.B1(n_119),
.B2(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_164),
.B1(n_143),
.B2(n_127),
.Y(n_181)
);

OAI22x1_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_124),
.B1(n_119),
.B2(n_125),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_133),
.C(n_147),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_182),
.C(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_177),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_154),
.B1(n_159),
.B2(n_162),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_145),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_128),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_188),
.C(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_159),
.C(n_157),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_171),
.C(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_154),
.B1(n_172),
.B2(n_175),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_180),
.B(n_174),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_205),
.B(n_187),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_189),
.B1(n_161),
.B2(n_150),
.Y(n_209)
);

AOI221xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_179),
.B1(n_175),
.B2(n_180),
.C(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_211),
.C(n_200),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_179),
.B1(n_186),
.B2(n_188),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_126),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_207),
.C(n_206),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_13),
.B(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.C(n_97),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_214),
.B1(n_220),
.B2(n_217),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_223),
.B(n_5),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_15),
.B(n_6),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_5),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_97),
.Y(n_227)
);


endmodule