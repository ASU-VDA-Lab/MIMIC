module fake_jpeg_13659_n_561 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_561);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_61),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_7),
.C(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_18),
.B(n_7),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_76),
.Y(n_132)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_79),
.B(n_118),
.Y(n_198)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_15),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_106),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_96),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_20),
.B(n_6),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_112),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_117),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_121),
.Y(n_149)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_48),
.B(n_0),
.CON(n_117),
.SN(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_24),
.B(n_5),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_8),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g122 ( 
.A(n_48),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g193 ( 
.A(n_122),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_64),
.A2(n_44),
.B1(n_51),
.B2(n_49),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_125),
.A2(n_128),
.B1(n_134),
.B2(n_147),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_60),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_127),
.A2(n_137),
.B1(n_148),
.B2(n_179),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_65),
.A2(n_44),
.B1(n_51),
.B2(n_54),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_44),
.B1(n_51),
.B2(n_49),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_91),
.A2(n_56),
.B1(n_46),
.B2(n_45),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_77),
.A2(n_34),
.B1(n_43),
.B2(n_39),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_75),
.A2(n_56),
.B1(n_46),
.B2(n_45),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_153),
.A2(n_166),
.B1(n_180),
.B2(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_31),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_154),
.B(n_169),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_33),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_168),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_75),
.A2(n_56),
.B1(n_40),
.B2(n_41),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_103),
.B(n_43),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_39),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_105),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_107),
.A2(n_56),
.B1(n_59),
.B2(n_37),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_61),
.A2(n_83),
.B1(n_94),
.B2(n_88),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_189),
.B1(n_116),
.B2(n_121),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_87),
.B(n_59),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_190),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_72),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_195),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_117),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_66),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_3),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_97),
.B(n_3),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_78),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_196),
.B1(n_67),
.B2(n_123),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_114),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_204),
.B(n_207),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_205),
.Y(n_300)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_209),
.A2(n_185),
.B1(n_194),
.B2(n_171),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_99),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_210),
.B(n_218),
.Y(n_295)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_230),
.B(n_239),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_115),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_162),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_222),
.A2(n_240),
.B1(n_264),
.B2(n_157),
.Y(n_291)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_226),
.B(n_231),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_0),
.B1(n_14),
.B2(n_132),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_0),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_232),
.Y(n_315)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_175),
.B(n_0),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_234),
.A2(n_265),
.B(n_272),
.Y(n_288)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_158),
.B(n_144),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_181),
.A2(n_142),
.B1(n_149),
.B2(n_135),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_172),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_248),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_255),
.Y(n_283)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_259),
.Y(n_289)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_174),
.B(n_173),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_252),
.B(n_253),
.C(n_271),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_173),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_258),
.B(n_262),
.Y(n_323)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_261),
.Y(n_305)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_139),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_139),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_187),
.A2(n_127),
.B(n_180),
.C(n_166),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_266),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_128),
.A2(n_147),
.B1(n_200),
.B2(n_146),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_151),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_151),
.B(n_167),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_269),
.B(n_234),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_167),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_161),
.C(n_195),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_130),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_132),
.B1(n_152),
.B2(n_141),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_286),
.A2(n_243),
.B(n_241),
.Y(n_342)
);

AO21x2_ASAP7_75t_L g287 ( 
.A1(n_220),
.A2(n_200),
.B(n_146),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_287),
.A2(n_205),
.B1(n_254),
.B2(n_211),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_290),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_291),
.A2(n_308),
.B1(n_316),
.B2(n_229),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_218),
.A2(n_157),
.B1(n_183),
.B2(n_185),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_296),
.B1(n_301),
.B2(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_225),
.B1(n_240),
.B2(n_212),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_267),
.A2(n_141),
.B1(n_171),
.B2(n_194),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_222),
.A2(n_126),
.B1(n_264),
.B2(n_263),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_210),
.A2(n_215),
.B1(n_268),
.B2(n_239),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_320),
.B1(n_236),
.B2(n_237),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_285),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_230),
.A2(n_252),
.B1(n_253),
.B2(n_239),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_252),
.C(n_253),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_322),
.C(n_310),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_245),
.A2(n_248),
.B1(n_256),
.B2(n_249),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_238),
.B(n_223),
.C(n_265),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_261),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_327),
.B(n_351),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_224),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_347),
.Y(n_370)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_262),
.B(n_242),
.C(n_233),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_330),
.A2(n_342),
.B(n_337),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_331),
.B(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_333),
.A2(n_335),
.B1(n_344),
.B2(n_367),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_295),
.B(n_259),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_302),
.A2(n_257),
.B(n_251),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_337),
.A2(n_342),
.B(n_363),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_216),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_338),
.B(n_343),
.Y(n_379)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_341),
.A2(n_362),
.B1(n_364),
.B2(n_274),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_289),
.B(n_314),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_291),
.A2(n_308),
.B1(n_287),
.B2(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_310),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_346),
.B(n_303),
.Y(n_372)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_349),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_289),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_294),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_352),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_277),
.B(n_280),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_355),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_283),
.B(n_324),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g391 ( 
.A1(n_354),
.A2(n_298),
.B(n_327),
.Y(n_391)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g369 ( 
.A1(n_356),
.A2(n_360),
.B(n_365),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_273),
.C(n_284),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_283),
.B(n_317),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_346),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_359),
.Y(n_375)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_361),
.B(n_363),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_304),
.A2(n_293),
.B1(n_287),
.B2(n_275),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_292),
.B(n_286),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_287),
.A2(n_275),
.B1(n_299),
.B2(n_320),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_299),
.A2(n_287),
.B1(n_286),
.B2(n_290),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_366),
.A2(n_273),
.B(n_284),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_282),
.A2(n_319),
.B1(n_274),
.B2(n_297),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_368),
.A2(n_374),
.B1(n_382),
.B2(n_388),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_372),
.B(n_383),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_312),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_373),
.B(n_380),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_328),
.A2(n_297),
.B1(n_307),
.B2(n_326),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_307),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_381),
.A2(n_384),
.B(n_398),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_334),
.A2(n_326),
.B1(n_300),
.B2(n_276),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_349),
.A2(n_276),
.B(n_313),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_313),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_386),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_278),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_334),
.A2(n_300),
.B1(n_298),
.B2(n_278),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_391),
.B(n_392),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_336),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_394),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_348),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_350),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_399),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_340),
.C(n_345),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_401),
.B(n_339),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_366),
.B(n_364),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_404),
.A2(n_427),
.B(n_394),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_376),
.A2(n_362),
.B1(n_329),
.B2(n_332),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_405),
.A2(n_393),
.B1(n_374),
.B2(n_380),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_398),
.A2(n_352),
.B(n_353),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_371),
.B(n_333),
.Y(n_410)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_410),
.Y(n_457)
);

AOI22x1_ASAP7_75t_SL g411 ( 
.A1(n_382),
.A2(n_344),
.B1(n_388),
.B2(n_390),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_411),
.A2(n_372),
.B(n_384),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_377),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_413),
.Y(n_434)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_417),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_378),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_416),
.B(n_419),
.Y(n_455)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_389),
.B(n_355),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_421),
.Y(n_440)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_389),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_397),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_375),
.A2(n_367),
.B1(n_335),
.B2(n_341),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_423),
.A2(n_376),
.B1(n_375),
.B2(n_397),
.Y(n_436)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_430),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_381),
.A2(n_330),
.B(n_356),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_386),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_347),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_432),
.Y(n_454)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_433),
.B(n_408),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_436),
.A2(n_453),
.B1(n_427),
.B2(n_431),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_438),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_379),
.B1(n_402),
.B2(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_443),
.A2(n_459),
.B1(n_404),
.B2(n_425),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_430),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_444),
.B(n_420),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_385),
.C(n_383),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_448),
.C(n_452),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_392),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_447),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_373),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_390),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_403),
.Y(n_469)
);

XOR2x1_ASAP7_75t_SL g482 ( 
.A(n_450),
.B(n_451),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_408),
.B(n_369),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_360),
.C(n_365),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_404),
.A2(n_335),
.B1(n_423),
.B2(n_410),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_335),
.Y(n_456)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_412),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_432),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_405),
.A2(n_335),
.B1(n_416),
.B2(n_419),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_434),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_473),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_467),
.Y(n_485)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_463),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_451),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_417),
.B1(n_415),
.B2(n_418),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

OA21x2_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_425),
.B(n_418),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_429),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_475),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_469),
.B(n_411),
.Y(n_489)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_440),
.Y(n_470)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_477),
.B1(n_481),
.B2(n_458),
.Y(n_495)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g476 ( 
.A(n_435),
.B(n_427),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_476),
.A2(n_411),
.B(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_424),
.C(n_407),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.C(n_447),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_424),
.C(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_SL g505 ( 
.A(n_487),
.B(n_472),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_433),
.C(n_443),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_490),
.C(n_497),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_494),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_435),
.C(n_446),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_455),
.Y(n_491)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_491),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_464),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_448),
.Y(n_494)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_450),
.C(n_449),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_476),
.B(n_474),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_439),
.Y(n_499)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_454),
.C(n_437),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_488),
.C(n_490),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_511),
.B(n_503),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_486),
.A2(n_483),
.B1(n_465),
.B2(n_453),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_507),
.A2(n_460),
.B1(n_457),
.B2(n_481),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_516),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_461),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_513),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_510),
.A2(n_498),
.B(n_484),
.Y(n_523)
);

AOI31xp33_ASAP7_75t_L g511 ( 
.A1(n_496),
.A2(n_470),
.A3(n_463),
.B(n_473),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_462),
.C(n_469),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_517),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_469),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_467),
.C(n_475),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_515),
.A2(n_497),
.B1(n_485),
.B2(n_500),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_520),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_502),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_514),
.Y(n_522)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_522),
.Y(n_532)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_524),
.A2(n_530),
.B(n_437),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_492),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_526),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_484),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_529),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_421),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_516),
.B(n_504),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_506),
.C(n_507),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_535),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_494),
.C(n_504),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_454),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_538),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_477),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_540),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_518),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_543),
.B(n_544),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_523),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_521),
.C(n_525),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_546),
.B(n_547),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_489),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g548 ( 
.A(n_541),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_542),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_545),
.A2(n_539),
.B(n_536),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_549),
.A2(n_551),
.B(n_547),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_545),
.A2(n_537),
.B(n_532),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_553),
.A2(n_456),
.B(n_426),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_552),
.B(n_550),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_554),
.B(n_555),
.C(n_460),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_557),
.B(n_409),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_558),
.A2(n_413),
.B(n_482),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_482),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_415),
.B(n_524),
.Y(n_561)
);


endmodule