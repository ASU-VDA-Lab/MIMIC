module fake_ariane_1556_n_113 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_25, n_113);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_113;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_106;
wire n_111;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_100;
wire n_62;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_82;
wire n_57;
wire n_70;
wire n_85;
wire n_94;
wire n_101;
wire n_58;
wire n_65;
wire n_112;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_81;
wire n_87;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_54;

INVx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_26),
.B1(n_33),
.B2(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_10),
.A2(n_14),
.B(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_21),
.B(n_9),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_37),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_4),
.B1(n_24),
.B2(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

OAI21x1_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_53),
.B(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_6),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_22),
.A2(n_1),
.B1(n_8),
.B2(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_2),
.B(n_5),
.C(n_12),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_19),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_41),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_74),
.B(n_56),
.C(n_61),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_70),
.B(n_57),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_67),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_60),
.B(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

AO21x2_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_85),
.B(n_83),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_89),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_66),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_96),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_58),
.A3(n_86),
.B1(n_103),
.B2(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_104),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_108),
.B(n_45),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_42),
.B(n_47),
.Y(n_113)
);


endmodule