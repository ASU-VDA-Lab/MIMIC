module fake_jpeg_28270_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx10_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_22),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_24),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_60),
.B1(n_27),
.B2(n_36),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_27),
.B1(n_35),
.B2(n_13),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

OR2x4_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_40),
.Y(n_62)
);

NOR2x1_ASAP7_75t_R g84 ( 
.A(n_62),
.B(n_31),
.Y(n_84)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_36),
.B1(n_34),
.B2(n_27),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_32),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_21),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_13),
.B1(n_63),
.B2(n_19),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_45),
.B1(n_35),
.B2(n_36),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_59),
.B1(n_47),
.B2(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_106),
.B1(n_95),
.B2(n_97),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_52),
.B1(n_79),
.B2(n_81),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_18),
.B1(n_19),
.B2(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_105),
.B1(n_34),
.B2(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_31),
.B(n_37),
.C(n_33),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_84),
.B1(n_86),
.B2(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_115),
.B1(n_122),
.B2(n_106),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_107),
.B1(n_123),
.B2(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_86),
.B1(n_87),
.B2(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_70),
.B1(n_18),
.B2(n_80),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_38),
.B1(n_47),
.B2(n_80),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_129),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_107),
.B1(n_99),
.B2(n_100),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_56),
.B(n_31),
.C(n_55),
.Y(n_170)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_135),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_106),
.B(n_104),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_137),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_138),
.B1(n_78),
.B2(n_82),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_125),
.B(n_111),
.Y(n_137)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_144),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_89),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_143),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_148),
.B1(n_37),
.B2(n_28),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_104),
.B(n_35),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_104),
.B1(n_77),
.B2(n_78),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_104),
.B(n_77),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_104),
.B1(n_78),
.B2(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_77),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_149),
.B(n_153),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_116),
.C(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_142),
.C(n_151),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_175),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_34),
.B1(n_94),
.B2(n_37),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_37),
.B1(n_55),
.B2(n_51),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_176),
.Y(n_179)
);

OAI22x1_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_139),
.B1(n_146),
.B2(n_42),
.Y(n_189)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_30),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_174),
.B1(n_16),
.B2(n_12),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_12),
.B1(n_46),
.B2(n_64),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_61),
.B1(n_12),
.B2(n_16),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_170),
.Y(n_206)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_185),
.B(n_188),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_148),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_23),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_30),
.C(n_22),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_170),
.C(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_155),
.B(n_15),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_15),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_199),
.B1(n_20),
.B2(n_9),
.Y(n_208)
);

AOI22x1_ASAP7_75t_SL g195 ( 
.A1(n_157),
.A2(n_173),
.B1(n_168),
.B2(n_160),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_25),
.B1(n_20),
.B2(n_9),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_25),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_172),
.C(n_167),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_165),
.C(n_162),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_165),
.C(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_205),
.C(n_215),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_170),
.C(n_175),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_218),
.B1(n_0),
.B2(n_1),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_23),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_30),
.C(n_22),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_192),
.C(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_204),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_180),
.B1(n_189),
.B2(n_184),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_228),
.B1(n_231),
.B2(n_2),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_198),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_190),
.B(n_182),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_234),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_23),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_215),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_217),
.B1(n_201),
.B2(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_22),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_233),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_214),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_236),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_210),
.C(n_30),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_236),
.C(n_242),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_22),
.C(n_33),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_42),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_22),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_230),
.B(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_256),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_232),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_219),
.C(n_227),
.Y(n_253)
);

XOR2x2_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_231),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_258),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_247),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_265),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_250),
.B(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_3),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_266),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_264),
.C(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

AOI221xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_268),
.B(n_259),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_271),
.B(n_6),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_277),
.C(n_33),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_5),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_6),
.B(n_7),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_8),
.Y(n_284)
);

A2O1A1O1Ixp25_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_8),
.B(n_33),
.C(n_198),
.D(n_278),
.Y(n_285)
);


endmodule