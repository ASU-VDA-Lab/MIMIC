module fake_jpeg_20146_n_50 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_50);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_50;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_8),
.B1(n_16),
.B2(n_13),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_25),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_39),
.B1(n_23),
.B2(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_27),
.C(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_3),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_3),
.B(n_5),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_40),
.C(n_38),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B(n_41),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_43),
.B(n_27),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_21),
.B(n_9),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);


endmodule