module fake_netlist_1_8535_n_733 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_733);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_733;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g81 ( .A(n_1), .Y(n_81) );
INVx3_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
NOR2xp67_ASAP7_75t_L g84 ( .A(n_10), .B(n_9), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_29), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_75), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_55), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_9), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_79), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_49), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_70), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_73), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_32), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
OR2x2_ASAP7_75t_L g99 ( .A(n_74), .B(n_62), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_31), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_20), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_0), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_40), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_65), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_51), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_35), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_52), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_25), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_60), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_69), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_22), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_50), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_6), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_77), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_71), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_14), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_67), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_38), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_23), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_13), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_58), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_96), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_96), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
BUFx8_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_116), .B(n_1), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_100), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_104), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_103), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_92), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_90), .B(n_2), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_112), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_115), .A2(n_34), .B(n_76), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
BUFx8_ASAP7_75t_L g158 ( .A(n_99), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g160 ( .A1(n_89), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_95), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_83), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_102), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_106), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_102), .B(n_8), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_113), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_120), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_121), .A2(n_8), .B1(n_11), .B2(n_12), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_105), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_101), .B(n_39), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_85), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_141), .B(n_107), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx5_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_141), .B(n_128), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_132), .B(n_118), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_175), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_152), .B(n_128), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_175), .B(n_121), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g188 ( .A(n_136), .B(n_94), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_131), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_175), .B(n_124), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_132), .A2(n_133), .B1(n_171), .B2(n_168), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_175), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_133), .B(n_127), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_154), .B(n_139), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_137), .B(n_127), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
BUFx10_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_173), .B(n_86), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_174), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_167), .B(n_84), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_175), .B(n_124), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_167), .B(n_119), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_173), .B(n_81), .Y(n_208) );
INVxp67_ASAP7_75t_L g209 ( .A(n_139), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_131), .Y(n_211) );
BUFx10_ASAP7_75t_L g212 ( .A(n_154), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_151), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_131), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_175), .B(n_111), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_138), .B(n_81), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_136), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_138), .B(n_122), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_174), .Y(n_222) );
BUFx4f_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_174), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_136), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_154), .B(n_122), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_140), .B(n_119), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_148), .Y(n_229) );
INVxp33_ASAP7_75t_SL g230 ( .A(n_136), .Y(n_230) );
AND2x6_ASAP7_75t_L g231 ( .A(n_142), .B(n_117), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_140), .B(n_118), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_174), .B(n_111), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_143), .B(n_93), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_164), .B(n_93), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_174), .Y(n_238) );
INVx5_ASAP7_75t_L g239 ( .A(n_144), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_158), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_210), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_196), .A2(n_157), .B1(n_150), .B2(n_153), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_229), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_225), .B(n_169), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_214), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_213), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_233), .B(n_158), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_196), .A2(n_153), .B1(n_150), .B2(n_157), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_240), .B(n_158), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_203), .B(n_158), .Y(n_253) );
NOR2x1p5_ASAP7_75t_L g254 ( .A(n_217), .B(n_171), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_196), .A2(n_145), .B1(n_159), .B2(n_155), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_209), .A2(n_160), .B(n_172), .C(n_170), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_176), .B(n_171), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_209), .B(n_171), .Y(n_259) );
NAND3xp33_ASAP7_75t_SL g260 ( .A(n_186), .B(n_88), .C(n_143), .Y(n_260) );
NOR2xp33_ASAP7_75t_SL g261 ( .A(n_230), .B(n_88), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_220), .B(n_159), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_177), .A2(n_155), .B(n_145), .C(n_161), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_178), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_223), .A2(n_156), .B(n_163), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_237), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_203), .B(n_162), .Y(n_268) );
OAI22xp5_ASAP7_75t_SL g269 ( .A1(n_235), .A2(n_156), .B1(n_170), .B2(n_166), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_235), .B(n_170), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_185), .A2(n_161), .B(n_162), .C(n_163), .Y(n_271) );
AO22x1_ASAP7_75t_L g272 ( .A1(n_231), .A2(n_166), .B1(n_134), .B2(n_135), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_196), .A2(n_149), .B1(n_168), .B2(n_157), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_208), .A2(n_149), .B1(n_153), .B2(n_150), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_208), .A2(n_166), .B1(n_142), .B2(n_148), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
NOR2xp67_ASAP7_75t_L g278 ( .A(n_200), .B(n_142), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_216), .A2(n_144), .B1(n_147), .B2(n_146), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_226), .B(n_146), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_220), .B(n_144), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_216), .A2(n_144), .B1(n_147), .B2(n_146), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_232), .B(n_146), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_232), .B(n_135), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_226), .B(n_134), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_221), .B(n_147), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_180), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_199), .Y(n_288) );
OAI22xp5_ASAP7_75t_SL g289 ( .A1(n_235), .A2(n_156), .B1(n_13), .B2(n_14), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_182), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_200), .A2(n_156), .B1(n_15), .B2(n_16), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_206), .B(n_42), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_191), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_219), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_181), .B(n_11), .Y(n_295) );
NAND2x1p5_ASAP7_75t_L g296 ( .A(n_181), .B(n_15), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_231), .Y(n_297) );
AO22x1_ASAP7_75t_L g298 ( .A1(n_231), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_193), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_191), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_231), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_193), .A2(n_19), .B1(n_24), .B2(n_26), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_199), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_192), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_212), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_212), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_204), .A2(n_27), .B1(n_28), .B2(n_30), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_195), .B(n_234), .Y(n_308) );
AND2x6_ASAP7_75t_SL g309 ( .A(n_204), .B(n_36), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_257), .B(n_234), .Y(n_310) );
NOR2xp33_ASAP7_75t_R g311 ( .A(n_249), .B(n_188), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_266), .A2(n_269), .B(n_281), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_261), .A2(n_231), .B1(n_195), .B2(n_227), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_288), .B(n_222), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_245), .B(n_227), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_256), .A2(n_223), .B(n_187), .C(n_205), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_270), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_287), .B(n_190), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_263), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_256), .A2(n_197), .B(n_238), .C(n_215), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_267), .Y(n_324) );
OA22x2_ASAP7_75t_L g325 ( .A1(n_270), .A2(n_197), .B1(n_221), .B2(n_224), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_287), .A2(n_224), .B1(n_222), .B2(n_194), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
NOR2xp33_ASAP7_75t_R g328 ( .A(n_260), .B(n_288), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g329 ( .A(n_260), .B(n_179), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_245), .B(n_184), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_241), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_265), .B(n_239), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_299), .A2(n_238), .B1(n_239), .B2(n_179), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_262), .A2(n_238), .B(n_192), .C(n_236), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_286), .A2(n_238), .B(n_239), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_308), .A2(n_239), .B(n_236), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_265), .B(n_179), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_285), .B(n_179), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_299), .A2(n_207), .B1(n_201), .B2(n_198), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_246), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_278), .A2(n_207), .B(n_201), .C(n_198), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_284), .A2(n_183), .B(n_202), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_275), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_277), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_264), .A2(n_183), .B(n_218), .C(n_202), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_246), .B(n_183), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_283), .A2(n_183), .B(n_202), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g351 ( .A1(n_289), .A2(n_218), .B1(n_202), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_271), .A2(n_218), .B(n_43), .C(n_53), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_268), .A2(n_218), .B(n_54), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_253), .A2(n_37), .B(n_56), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_241), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_276), .A2(n_57), .B1(n_59), .B2(n_61), .C(n_63), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_243), .B(n_66), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_243), .B(n_80), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_303), .B(n_306), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_254), .B(n_251), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_255), .A2(n_251), .B1(n_273), .B2(n_279), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_274), .B(n_305), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_291), .B(n_292), .C(n_297), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_247), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_351), .A2(n_307), .B(n_282), .C(n_252), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_362), .B(n_272), .Y(n_366) );
AOI21xp5_ASAP7_75t_SL g367 ( .A1(n_317), .A2(n_250), .B(n_242), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_320), .B(n_295), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_312), .A2(n_248), .B(n_297), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_296), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_312), .A2(n_301), .B(n_241), .Y(n_373) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_344), .A2(n_293), .A3(n_304), .B(n_258), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_360), .A2(n_296), .B1(n_301), .B2(n_302), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_316), .B(n_309), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_346), .A2(n_302), .B1(n_242), .B2(n_241), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_242), .B(n_290), .Y(n_378) );
BUFx10_ASAP7_75t_L g379 ( .A(n_359), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_313), .B(n_242), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_337), .B(n_298), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_318), .A2(n_300), .B1(n_361), .B2(n_345), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_336), .B(n_310), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_331), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_350), .A2(n_323), .B(n_338), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_350), .A2(n_348), .B(n_338), .Y(n_386) );
INVx8_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_341), .A2(n_334), .B(n_343), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_319), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_347), .B(n_363), .C(n_352), .Y(n_390) );
INVx6_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_330), .B(n_314), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_332), .A2(n_333), .B(n_353), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
AO31x2_ASAP7_75t_L g395 ( .A1(n_357), .A2(n_358), .A3(n_353), .B(n_354), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_328), .B(n_364), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_356), .A2(n_321), .B(n_329), .C(n_326), .Y(n_397) );
BUFx10_ASAP7_75t_L g398 ( .A(n_340), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_372), .B(n_380), .Y(n_401) );
BUFx2_ASAP7_75t_R g402 ( .A(n_366), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_387), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_325), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_376), .A2(n_311), .B1(n_342), .B2(n_325), .C(n_335), .Y(n_407) );
OAI322xp33_ASAP7_75t_L g408 ( .A1(n_376), .A2(n_315), .A3(n_349), .B1(n_355), .B2(n_368), .C1(n_381), .C2(n_383), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_394), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_389), .B(n_379), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_394), .A2(n_375), .B1(n_377), .B2(n_397), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_393), .B(n_390), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_373), .B(n_370), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_379), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_387), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_374), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_392), .B(n_390), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_380), .B(n_371), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
OA21x2_ASAP7_75t_L g421 ( .A1(n_397), .A2(n_378), .B(n_377), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_367), .A2(n_382), .B(n_365), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_381), .A2(n_396), .B1(n_375), .B2(n_398), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_384), .B(n_399), .Y(n_424) );
OAI21x1_ASAP7_75t_L g425 ( .A1(n_384), .A2(n_399), .B(n_395), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_395), .A2(n_387), .B(n_391), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_391), .B1(n_395), .B2(n_256), .C(n_208), .Y(n_427) );
OAI21x1_ASAP7_75t_SL g428 ( .A1(n_391), .A2(n_393), .B(n_370), .Y(n_428) );
AO21x2_ASAP7_75t_L g429 ( .A1(n_422), .A2(n_395), .B(n_428), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_426), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_422), .A2(n_428), .B(n_417), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_411), .A2(n_423), .B1(n_427), .B2(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_408), .B(n_400), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_426), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_427), .A2(n_411), .B(n_417), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_406), .B(n_401), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_416), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
OR2x6_ASAP7_75t_L g441 ( .A(n_416), .B(n_420), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_409), .B(n_406), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_401), .B(n_404), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_419), .B(n_420), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_418), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_401), .B(n_404), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_418), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_413), .A2(n_425), .B(n_420), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_410), .B(n_419), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_419), .B(n_401), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_421), .B(n_413), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_425), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_419), .B(n_401), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_405), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_413), .A2(n_412), .B(n_424), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_419), .B(n_414), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_412), .B(n_426), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_412), .A2(n_424), .B(n_421), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_441), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_443), .B(n_412), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_433), .Y(n_468) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_433), .B(n_426), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_436), .B(n_405), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_444), .B(n_426), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_436), .B(n_405), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_439), .B(n_408), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_442), .B(n_415), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_445), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_445), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_444), .B(n_407), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_448), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_440), .B(n_405), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_440), .B(n_405), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_447), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_441), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_458), .B(n_424), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_443), .B(n_421), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_447), .Y(n_487) );
INVxp33_ASAP7_75t_L g488 ( .A(n_459), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_448), .B(n_421), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_448), .B(n_407), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_462), .B(n_421), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_432), .B(n_403), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_432), .B(n_403), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_454), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_462), .B(n_402), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_462), .B(n_402), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_458), .B(n_403), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_446), .B(n_415), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_446), .B(n_415), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_438), .B(n_464), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_438), .B(n_464), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_456), .B(n_437), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_454), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_458), .B(n_435), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_456), .B(n_442), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_449), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_430), .B(n_435), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_430), .B(n_431), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_485), .B(n_431), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_499), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_513), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_467), .B(n_431), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_467), .B(n_429), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_468), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_471), .B(n_452), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_499), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_471), .B(n_429), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_513), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_486), .B(n_429), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_469), .B(n_434), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_513), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_486), .B(n_449), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_503), .B(n_450), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_508), .B(n_449), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_449), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_503), .B(n_451), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_509), .B(n_434), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_509), .B(n_457), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_510), .B(n_457), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_510), .B(n_457), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_510), .B(n_461), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_478), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_485), .B(n_461), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_505), .B(n_461), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_504), .B(n_451), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_514), .B(n_463), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_505), .B(n_463), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_514), .B(n_463), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_469), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_474), .B(n_455), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_488), .B(n_455), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_514), .B(n_504), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_491), .B(n_515), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_483), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_485), .B(n_465), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_515), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_512), .B(n_492), .Y(n_559) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_496), .B(n_466), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_512), .B(n_492), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_487), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_491), .B(n_515), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_487), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_493), .B(n_502), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_493), .B(n_502), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_501), .B(n_475), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_470), .B(n_482), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_470), .B(n_482), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_494), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_470), .B(n_482), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_472), .B(n_481), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_479), .A2(n_474), .B1(n_490), .B2(n_501), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_466), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_521), .Y(n_576) );
NAND2x1_ASAP7_75t_SL g577 ( .A(n_574), .B(n_497), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_555), .B(n_489), .Y(n_578) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_560), .B(n_496), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_521), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_531), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_553), .B(n_490), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_551), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_553), .B(n_479), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_552), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_555), .B(n_558), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_568), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_532), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_550), .B(n_498), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_558), .B(n_500), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_563), .B(n_489), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_563), .B(n_480), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_538), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_568), .B(n_489), .Y(n_598) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_528), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_569), .B(n_472), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_574), .B(n_498), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_569), .B(n_472), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_522), .B(n_500), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_541), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_571), .B(n_481), .Y(n_606) );
NOR2xp33_ASAP7_75t_R g607 ( .A(n_560), .B(n_465), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_559), .B(n_494), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_567), .A2(n_498), .B1(n_497), .B2(n_484), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_527), .B(n_497), .C(n_506), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_571), .B(n_481), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_572), .B(n_465), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_561), .B(n_506), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_530), .B(n_480), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_572), .B(n_465), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_565), .B(n_473), .Y(n_618) );
AND3x2_ASAP7_75t_L g619 ( .A(n_575), .B(n_473), .C(n_476), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_566), .B(n_535), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_518), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_535), .B(n_473), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_520), .B(n_484), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_534), .B(n_476), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_529), .B(n_476), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_543), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_545), .B(n_477), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_529), .B(n_477), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_556), .B(n_477), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_581), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_584), .B(n_520), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_582), .B(n_526), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_589), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_588), .B(n_522), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_579), .A2(n_560), .B1(n_547), .B2(n_554), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_601), .A2(n_526), .B1(n_523), .B2(n_517), .C1(n_519), .C2(n_516), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_590), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_591), .B(n_524), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_579), .A2(n_547), .B1(n_550), .B2(n_524), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_596), .B(n_546), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_600), .B(n_557), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_621), .B(n_519), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_600), .B(n_557), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_586), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_601), .B(n_516), .C(n_547), .D(n_557), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_587), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_602), .B(n_547), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_611), .Y(n_652) );
NOR2xp67_ASAP7_75t_L g653 ( .A(n_612), .B(n_528), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_625), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_609), .B(n_532), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_602), .B(n_540), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_583), .B(n_562), .C(n_556), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_628), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_615), .B(n_595), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_578), .B(n_544), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_597), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_626), .B(n_546), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_604), .Y(n_664) );
AOI321xp33_ASAP7_75t_L g665 ( .A1(n_592), .A2(n_516), .A3(n_557), .B1(n_544), .B2(n_548), .C(n_540), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_611), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_605), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_585), .B(n_564), .Y(n_668) );
AOI31xp33_ASAP7_75t_L g669 ( .A1(n_592), .A2(n_516), .A3(n_564), .B(n_562), .Y(n_669) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_637), .A2(n_610), .B(n_603), .C(n_618), .Y(n_670) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_657), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g672 ( .A1(n_634), .A2(n_578), .A3(n_595), .B1(n_606), .B2(n_613), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_651), .B(n_606), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_631), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_651), .B(n_613), .Y(n_675) );
OAI22xp33_ASAP7_75t_SL g676 ( .A1(n_652), .A2(n_593), .B1(n_603), .B2(n_577), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_638), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_665), .A2(n_593), .B(n_599), .C(n_624), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_663), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_663), .B(n_598), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_666), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_669), .A2(n_608), .B(n_627), .Y(n_683) );
AOI221x1_ASAP7_75t_SL g684 ( .A1(n_668), .A2(n_616), .B1(n_620), .B2(n_623), .C(n_570), .Y(n_684) );
AO22x1_ASAP7_75t_L g685 ( .A1(n_640), .A2(n_607), .B1(n_614), .B2(n_617), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_635), .Y(n_686) );
INVx1_ASAP7_75t_SL g687 ( .A(n_654), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_639), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_666), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_658), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_636), .A2(n_630), .B(n_594), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_668), .A2(n_570), .B(n_624), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_649), .A2(n_619), .B(n_617), .Y(n_693) );
AOI211xp5_ASAP7_75t_SL g694 ( .A1(n_676), .A2(n_652), .B(n_653), .C(n_657), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_655), .B1(n_633), .B2(n_632), .C(n_659), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_679), .B(n_607), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_679), .A2(n_644), .B(n_660), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_672), .A2(n_643), .B(n_646), .C(n_656), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_693), .A2(n_656), .B(n_642), .C(n_662), .Y(n_699) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_687), .B(n_667), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_680), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_671), .A2(n_664), .B1(n_647), .B2(n_661), .C(n_650), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_671), .B(n_648), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_682), .B(n_645), .C(n_641), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_683), .A2(n_484), .B1(n_598), .B2(n_614), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_686), .B(n_622), .Y(n_706) );
AOI322xp5_ASAP7_75t_L g707 ( .A1(n_690), .A2(n_548), .A3(n_539), .B1(n_537), .B2(n_549), .C1(n_622), .C2(n_542), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_670), .A2(n_692), .B1(n_689), .B2(n_682), .C(n_677), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_696), .B(n_685), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_700), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_708), .B(n_699), .C(n_702), .Y(n_711) );
XOR2xp5_ASAP7_75t_L g712 ( .A(n_703), .B(n_674), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_697), .A2(n_689), .B1(n_691), .B2(n_688), .C(n_681), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_701), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_694), .A2(n_678), .B(n_675), .C(n_673), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_L g716 ( .A1(n_698), .A2(n_528), .B(n_525), .C(n_518), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g717 ( .A1(n_707), .A2(n_695), .B(n_704), .C(n_706), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_711), .B(n_705), .C(n_528), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_710), .Y(n_719) );
AOI211xp5_ASAP7_75t_SL g720 ( .A1(n_717), .A2(n_484), .B(n_536), .C(n_542), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_715), .B(n_525), .C(n_536), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_712), .B(n_542), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_720), .A2(n_713), .B(n_716), .C(n_714), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_719), .B(n_709), .C(n_525), .Y(n_724) );
NAND5xp2_ASAP7_75t_L g725 ( .A(n_718), .B(n_537), .C(n_539), .D(n_549), .E(n_542), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_723), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_725), .B(n_721), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_726), .B(n_722), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_728), .Y(n_729) );
AO21x1_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_727), .B(n_724), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_730), .B(n_573), .C(n_495), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_731), .A2(n_573), .B1(n_495), .B2(n_507), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_732), .A2(n_573), .B1(n_480), .B2(n_511), .Y(n_733) );
endmodule