module fake_jpeg_15904_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_74),
.Y(n_107)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_46),
.Y(n_104)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_42),
.B1(n_60),
.B2(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_58),
.B1(n_59),
.B2(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_55),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_1),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_73),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_3),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_51),
.B1(n_56),
.B2(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_82),
.B1(n_54),
.B2(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_69),
.B1(n_41),
.B2(n_53),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_121)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_49),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_2),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_98),
.B1(n_97),
.B2(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_121),
.B(n_92),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_123),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_4),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_107),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_131),
.B(n_109),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_112),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_114),
.B1(n_90),
.B2(n_106),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_101),
.B1(n_115),
.B2(n_117),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_121),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_125),
.C(n_113),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_140),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_125),
.B1(n_91),
.B2(n_49),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_125),
.B1(n_54),
.B2(n_7),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_139),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_144),
.B1(n_143),
.B2(n_141),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_147),
.B1(n_135),
.B2(n_19),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_18),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_151),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_16),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_20),
.B(n_36),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_15),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_14),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_22),
.B(n_30),
.C(n_29),
.D(n_28),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_113),
.C(n_13),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_11),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_10),
.Y(n_161)
);


endmodule