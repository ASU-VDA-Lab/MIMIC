module fake_jpeg_13816_n_434 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_434);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_434;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_18),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_63),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_84),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_88),
.Y(n_115)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_1),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_76),
.B(n_26),
.Y(n_96)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_24),
.A2(n_1),
.B(n_3),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_85),
.B(n_90),
.Y(n_130)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_87),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_36),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_92),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_95),
.A2(n_97),
.B1(n_108),
.B2(n_121),
.Y(n_157)
);

OR2x2_ASAP7_75t_SL g183 ( 
.A(n_96),
.B(n_11),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_39),
.B1(n_37),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_127),
.B1(n_66),
.B2(n_56),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_37),
.B1(n_43),
.B2(n_32),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_49),
.A2(n_46),
.B1(n_45),
.B2(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_123),
.B1(n_13),
.B2(n_11),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_43),
.B1(n_37),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_32),
.B1(n_42),
.B2(n_24),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_30),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_28),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_77),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_72),
.A2(n_44),
.B1(n_28),
.B2(n_26),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_61),
.A3(n_69),
.B1(n_82),
.B2(n_85),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_44),
.B1(n_35),
.B2(n_34),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_12),
.B1(n_95),
.B2(n_97),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_50),
.B(n_35),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_11),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_145),
.B(n_147),
.Y(n_214)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_65),
.B1(n_78),
.B2(n_23),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_148),
.A2(n_182),
.B(n_119),
.Y(n_230)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_150),
.A2(n_114),
.B1(n_134),
.B2(n_110),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_151),
.A2(n_155),
.B1(n_193),
.B2(n_103),
.Y(n_232)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_61),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_105),
.C(n_144),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_47),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_177),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_87),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_169),
.Y(n_203)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_87),
.B1(n_4),
.B2(n_5),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_117),
.B1(n_133),
.B2(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_168),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_3),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_171),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_130),
.B1(n_103),
.B2(n_114),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_6),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_173),
.B(n_175),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_178),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_117),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_101),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_10),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

OR2x4_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_10),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_12),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_164),
.B1(n_172),
.B2(n_176),
.Y(n_197)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_190),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_11),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_197),
.A2(n_201),
.B1(n_196),
.B2(n_194),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_224),
.B1(n_232),
.B2(n_157),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_202),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_154),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_169),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_180),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_135),
.B1(n_109),
.B2(n_113),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_135),
.B1(n_113),
.B2(n_111),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_216),
.A2(n_198),
.B(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_126),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_231),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_233),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_162),
.B(n_185),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_126),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_183),
.B(n_110),
.CI(n_134),
.CON(n_233),
.SN(n_233)
);

O2A1O1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_12),
.B(n_101),
.C(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_151),
.B1(n_167),
.B2(n_148),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_236),
.A2(n_251),
.B1(n_252),
.B2(n_262),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_249),
.B1(n_256),
.B2(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_203),
.B(n_160),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_239),
.B(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_241),
.B(n_226),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_154),
.C(n_171),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_245),
.C(n_269),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_209),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_158),
.C(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_193),
.B1(n_150),
.B2(n_147),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_258),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_152),
.B1(n_166),
.B2(n_190),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_184),
.B1(n_165),
.B2(n_161),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_189),
.B(n_181),
.C(n_146),
.D(n_188),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_253),
.A2(n_220),
.B(n_229),
.Y(n_291)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_187),
.B1(n_163),
.B2(n_179),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_163),
.B1(n_192),
.B2(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_203),
.B(n_208),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_214),
.B(n_207),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_224),
.A2(n_221),
.B1(n_196),
.B2(n_210),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_236),
.B1(n_262),
.B2(n_251),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_207),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_267),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_200),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_223),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_210),
.A2(n_227),
.B(n_235),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_272),
.B(n_209),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_227),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_235),
.B1(n_233),
.B2(n_215),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_233),
.B1(n_225),
.B2(n_217),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_278),
.B1(n_272),
.B2(n_254),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_238),
.A2(n_217),
.B1(n_218),
.B2(n_226),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_296),
.C(n_304),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_280),
.A2(n_282),
.B(n_287),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_223),
.B(n_234),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_299),
.B(n_241),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_260),
.Y(n_288)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_303),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_220),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_293),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_218),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_295),
.B(n_300),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_242),
.C(n_245),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_273),
.A2(n_249),
.B(n_264),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_247),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_302),
.A2(n_257),
.B1(n_256),
.B2(n_246),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_268),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_248),
.C(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_240),
.B(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_252),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_266),
.C(n_263),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_320),
.C(n_321),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_312),
.A2(n_319),
.B1(n_333),
.B2(n_286),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_284),
.B1(n_290),
.B2(n_281),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_274),
.A2(n_246),
.B1(n_253),
.B2(n_271),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_255),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_270),
.C(n_279),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_323),
.B(n_330),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_280),
.A2(n_299),
.B(n_291),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_331),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_305),
.C(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_329),
.C(n_284),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_277),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_282),
.A2(n_277),
.B(n_302),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_276),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_332),
.B(n_334),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_274),
.A2(n_278),
.B1(n_275),
.B2(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_290),
.A2(n_306),
.B(n_293),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_283),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_343),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_338),
.A2(n_345),
.B1(n_312),
.B2(n_328),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_343),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_333),
.A2(n_295),
.B1(n_276),
.B2(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_349),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_297),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_303),
.B1(n_298),
.B2(n_301),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_298),
.C(n_301),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_354),
.C(n_308),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_292),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_356),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_319),
.A2(n_286),
.B1(n_324),
.B2(n_311),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_316),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_358),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_286),
.C(n_327),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_330),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_316),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_357),
.B(n_331),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_344),
.C(n_339),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_363),
.C(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_323),
.C(n_318),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_325),
.C(n_328),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_366),
.B(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_372),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_350),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_371),
.B(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_345),
.A2(n_334),
.B1(n_310),
.B2(n_315),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_374),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_342),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_356),
.Y(n_384)
);

AND3x1_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_322),
.C(n_326),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_378),
.A2(n_340),
.B(n_341),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_367),
.A2(n_340),
.B(n_336),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_388),
.B(n_367),
.Y(n_402)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_377),
.B(n_348),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_386),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_335),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_346),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_370),
.C(n_354),
.Y(n_405)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_392),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_379),
.B(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_399),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_397),
.A2(n_403),
.B(n_380),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_379),
.B(n_373),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_387),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_386),
.B(n_364),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_344),
.Y(n_400)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_400),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_405),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_375),
.B(n_376),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_407),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_381),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_397),
.A2(n_375),
.B1(n_361),
.B2(n_352),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_409),
.A2(n_411),
.B(n_388),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_395),
.B(n_385),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_395),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_404),
.A2(n_390),
.B(n_382),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_414),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_362),
.B1(n_365),
.B2(n_374),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_400),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_421),
.B(n_391),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_390),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_419),
.B(n_420),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_403),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_410),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_423),
.A2(n_426),
.B(n_394),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_424),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_SL g426 ( 
.A1(n_416),
.A2(n_394),
.B(n_389),
.C(n_372),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_425),
.B(n_417),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_429),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_428),
.B1(n_418),
.B2(n_407),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_431),
.B(n_405),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_422),
.C(n_370),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_368),
.C(n_322),
.Y(n_434)
);


endmodule