module real_jpeg_16096_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_41),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_0),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_108),
.Y(n_107)
);

NAND2x1_ASAP7_75t_SL g128 ( 
.A(n_0),
.B(n_129),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_41),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_84),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_6),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_6),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_6),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_7),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_8),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_11),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_183),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_145),
.B(n_182),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_117),
.B(n_144),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_89),
.B(n_116),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_18),
.B(n_52),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.C(n_46),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_19)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_20),
.A2(n_35),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

O2A1O1Ixp5_ASAP7_75t_L g152 ( 
.A1(n_20),
.A2(n_98),
.B(n_107),
.C(n_135),
.Y(n_152)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_26),
.A2(n_27),
.B1(n_123),
.B2(n_130),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_31),
.C(n_35),
.Y(n_88)
);

OR2x4_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_44),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_30),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_32),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_37),
.A2(n_38),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_42),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_42),
.A2(n_43),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_57),
.B(n_68),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_49),
.B(n_95),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_71),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_72),
.C(n_88),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_62),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_104),
.B(n_109),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_55),
.A2(n_63),
.B(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_92),
.B(n_94),
.C(n_98),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_92),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_69),
.B1(n_92),
.B2(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_68),
.B(n_123),
.C(n_128),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_87),
.B2(n_88),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_86),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_79),
.C(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_82),
.B(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_102),
.B(n_115),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_106),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_107),
.C(n_166),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_92),
.A2(n_113),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_95),
.A2(n_96),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_95),
.B(n_141),
.C(n_157),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_111),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_110),
.B(n_114),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_106),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_107),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_119),
.Y(n_144)
);

XOR2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_131),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_131),
.C(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_139),
.C(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_147),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_149),
.B(n_150),
.C(n_161),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_155),
.C(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_181),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_169),
.C(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_175),
.B(n_180),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_175),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_220),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_219),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_219),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_202),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_200),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_218),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);


endmodule