module real_jpeg_2731_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_41),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_1),
.B(n_26),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_3),
.B(n_44),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_3),
.B(n_35),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_32),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_3),
.B(n_78),
.Y(n_281)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_26),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_51),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_4),
.B(n_41),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_4),
.B(n_44),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_4),
.B(n_32),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_5),
.B(n_51),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_35),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_32),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_78),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_63),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_6),
.B(n_35),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_8),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_8),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_26),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_8),
.B(n_41),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_8),
.B(n_44),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_8),
.B(n_32),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_8),
.B(n_35),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_8),
.B(n_78),
.Y(n_294)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_13),
.B(n_51),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_13),
.B(n_26),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_41),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_44),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_32),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_41),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_14),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_14),
.B(n_78),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_19),
.B(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_81),
.C(n_92),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_81),
.CI(n_92),
.CON(n_149),
.SN(n_149)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_21),
.B(n_61),
.C(n_72),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.C(n_47),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_22),
.A2(n_23),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_24),
.B(n_33),
.C(n_38),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_31),
.A2(n_38),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_31),
.B(n_213),
.C(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_31),
.A2(n_38),
.B1(n_213),
.B2(n_219),
.Y(n_218)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_33),
.A2(n_34),
.B1(n_77),
.B2(n_101),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_33),
.A2(n_34),
.B1(n_174),
.B2(n_252),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_75),
.C(n_77),
.Y(n_74)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_36),
.B(n_171),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_38),
.B(n_85),
.C(n_86),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_39),
.B(n_47),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_40),
.B(n_43),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_41),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_42),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_42),
.A2(n_84),
.B1(n_85),
.B2(n_95),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_42),
.B(n_85),
.C(n_193),
.Y(n_232)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_57),
.C(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_57),
.A2(n_58),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_58),
.B(n_139),
.C(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_67),
.C(n_69),
.Y(n_132)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_115),
.C(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_67),
.A2(n_68),
.B1(n_115),
.B2(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.C(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_74),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_100),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_77),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_77),
.A2(n_101),
.B1(n_269),
.B2(n_270),
.Y(n_282)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_78),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_114),
.C(n_120),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_111),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_80),
.A2(n_111),
.B1(n_120),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_85),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.C(n_113),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_93),
.B(n_108),
.CI(n_113),
.CON(n_151),
.SN(n_151)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_104),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_94),
.B(n_98),
.Y(n_358)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_99),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_99),
.A2(n_100),
.B1(n_209),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_101),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_102),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_103),
.A2(n_185),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_104),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_116),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_119),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_119),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_143),
.B2(n_144),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_133),
.B2(n_142),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_138),
.A2(n_139),
.B1(n_161),
.B2(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_177),
.B(n_372),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_149),
.B(n_150),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_149),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.C(n_155),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_151),
.B(n_152),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_151),
.Y(n_373)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_155),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.C(n_167),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_156),
.A2(n_157),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_158),
.B(n_160),
.CI(n_162),
.CON(n_334),
.SN(n_334)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_165),
.B(n_167),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.C(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_168),
.A2(n_169),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_173),
.A2(n_174),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_173),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_174),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_175),
.A2(n_176),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_176),
.Y(n_346)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI31xp33_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_348),
.A3(n_361),
.B(n_366),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_328),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_253),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_226),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_182),
.B(n_226),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.C(n_216),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_183),
.B(n_325),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_183),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.CI(n_192),
.CON(n_183),
.SN(n_183)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_188),
.C(n_192),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_187),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_186),
.B(n_187),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_191),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_194),
.B(n_210),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_194),
.B(n_237),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_196),
.B(n_216),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_206),
.B2(n_215),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_207),
.C(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_203),
.C(n_205),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_202),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_224),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_217),
.B(n_220),
.CI(n_224),
.CON(n_315),
.SN(n_315)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_221),
.B(n_223),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_264),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_226),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_243),
.CI(n_244),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_227),
.B(n_243),
.C(n_244),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_228),
.B(n_231),
.C(n_238),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_238),
.B2(n_239),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_232),
.B(n_234),
.C(n_236),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_246),
.B(n_247),
.C(n_249),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_323),
.B(n_327),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_311),
.B(n_322),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_283),
.B(n_310),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_274),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_261),
.CI(n_262),
.CON(n_275),
.SN(n_275)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_272),
.C(n_273),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.C(n_282),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_307),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_275),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_277),
.B1(n_282),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_304),
.B(n_309),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_295),
.B(n_303),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.B(n_302),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_318),
.C(n_319),
.Y(n_326)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_315),
.Y(n_376)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_347),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_347),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_333),
.C(n_336),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_334),
.Y(n_380)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_341),
.C(n_342),
.Y(n_355)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_362),
.B(n_367),
.C(n_370),
.D(n_371),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_359),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_359),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.C(n_356),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_352),
.B1(n_356),
.B2(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_365),
.Y(n_370)
);


endmodule