module real_jpeg_11358_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_41),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_26),
.B1(n_30),
.B2(n_41),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_32),
.B(n_37),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_32),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_4),
.A2(n_75),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_22),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g55 ( 
.A1(n_12),
.A2(n_21),
.B(n_22),
.C(n_56),
.D(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_70),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_30),
.B(n_47),
.C(n_83),
.D(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_12),
.B(n_57),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_38),
.B(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_86),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_85),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_61),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_42),
.C(n_55),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_18),
.A2(n_19),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_31),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_48),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_33),
.A2(n_50),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_36),
.B(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_36),
.B(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_37),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_38),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_39),
.A2(n_112),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_39),
.B(n_119),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_42),
.A2(n_43),
.B1(n_55),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_54),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_52),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_54),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_79),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_78),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_129),
.B(n_135),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_108),
.B(n_128),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_92),
.B1(n_93),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_101),
.C(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_116),
.B(n_127),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_114),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_122),
.B(n_126),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);


endmodule