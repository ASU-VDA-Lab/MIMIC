module real_aes_3542_n_5 (n_4, n_0, n_3, n_2, n_1, n_5);
input n_4;
input n_0;
input n_3;
input n_2;
input n_1;
output n_5;
wire n_16;
wire n_13;
wire n_15;
wire n_7;
wire n_8;
wire n_6;
wire n_12;
wire n_9;
wire n_14;
wire n_10;
wire n_11;
BUFx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
OAI21xp5_ASAP7_75t_SL g6 ( .A1(n_1), .A2(n_4), .B(n_7), .Y(n_6) );
AND3x1_ASAP7_75t_L g16 ( .A(n_1), .B(n_10), .C(n_14), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g5 ( .A1(n_2), .A2(n_6), .B1(n_15), .B2(n_16), .Y(n_5) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_11), .Y(n_14) );
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_4), .A2(n_13), .B(n_14), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_11), .B(n_12), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
BUFx8_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
endmodule