module fake_jpeg_25619_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_6),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_5),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_62),
.B1(n_9),
.B2(n_11),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_35),
.B1(n_40),
.B2(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_62),
.B1(n_60),
.B2(n_55),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_55),
.Y(n_65)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_61),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_69),
.B(n_67),
.Y(n_74)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_66),
.CI(n_63),
.CON(n_73),
.SN(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_13),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_14),
.B(n_16),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_18),
.C(n_19),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_30),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_73),
.Y(n_83)
);


endmodule