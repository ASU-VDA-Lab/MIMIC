module fake_jpeg_1102_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_20),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_13),
.C(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_13),
.A2(n_17),
.B1(n_26),
.B2(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_24),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_26),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_23),
.B1(n_14),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_65),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22x1_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_22),
.B1(n_18),
.B2(n_7),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_45),
.B(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_8),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_74),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_41),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_62),
.C(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_64),
.C(n_68),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_71),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_75),
.C(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_75),
.B1(n_77),
.B2(n_60),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_48),
.C(n_52),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_81),
.B(n_82),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_94),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_89),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_48),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_18),
.C(n_22),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_97),
.A3(n_10),
.B1(n_11),
.B2(n_9),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_11),
.B(n_55),
.Y(n_101)
);


endmodule