module fake_jpeg_19445_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_21),
.B1(n_17),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_40),
.B1(n_13),
.B2(n_16),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_13),
.B1(n_18),
.B2(n_16),
.Y(n_40)
);

OR2x4_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_23),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_14),
.B(n_23),
.C(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_32),
.B1(n_29),
.B2(n_15),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_43),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_54),
.Y(n_57)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_12),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_25),
.C(n_27),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_53),
.C(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_66),
.B1(n_55),
.B2(n_53),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_63),
.B(n_31),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_43),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_14),
.C(n_10),
.Y(n_67)
);

BUFx12f_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_37),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_47),
.B1(n_25),
.B2(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_61),
.B(n_60),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_0),
.B(n_1),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_65),
.C(n_64),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_0),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_65),
.B1(n_62),
.B2(n_31),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_62),
.B1(n_74),
.B2(n_72),
.Y(n_88)
);

OA21x2_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_72),
.B(n_7),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_8),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_10),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_8),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_79),
.B1(n_80),
.B2(n_85),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_91),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_96),
.B(n_89),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_100),
.B(n_95),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_9),
.Y(n_106)
);


endmodule