module fake_netlist_6_1305_n_1084 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_265, n_113, n_39, n_63, n_223, n_270, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1084);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_270;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1084;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_683;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_138),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_134),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_191),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_101),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_116),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_209),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_240),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_185),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_157),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_243),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_100),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_180),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_192),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_73),
.Y(n_300)
);

HB1xp67_ASAP7_75t_SL g301 ( 
.A(n_172),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_215),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_85),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_171),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_14),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_122),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_127),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_228),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_210),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_137),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_41),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_187),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_107),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_235),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_245),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_259),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_57),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_217),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_129),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_125),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_238),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_130),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_184),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_67),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_244),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_41),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_31),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_119),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_136),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_36),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_86),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_275),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_283),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_330),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_277),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_277),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_278),
.B(n_0),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_280),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_276),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_282),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_278),
.B(n_314),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_287),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_288),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_280),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_292),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_281),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_304),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_301),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_293),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_378),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_328),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_361),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_337),
.A2(n_317),
.B1(n_306),
.B2(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_368),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_311),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_342),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_324),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_347),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_371),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_369),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_371),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_350),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_362),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_328),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_373),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_340),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_309),
.B(n_308),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_340),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_341),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_312),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_343),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_343),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_344),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_336),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_345),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_345),
.B(n_306),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_428),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_356),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_425),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_356),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_381),
.A2(n_365),
.B1(n_351),
.B2(n_406),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_425),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_317),
.B1(n_353),
.B2(n_336),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_359),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_381),
.B(n_375),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

NAND3xp33_ASAP7_75t_SL g448 ( 
.A(n_385),
.B(n_390),
.C(n_388),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_391),
.B(n_274),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

BUFx4f_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_354),
.C(n_349),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_381),
.B(n_327),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_394),
.B(n_303),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_349),
.C(n_348),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_303),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_384),
.B(n_333),
.Y(n_463)
);

INVx4_ASAP7_75t_SL g464 ( 
.A(n_382),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_400),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_426),
.B(n_284),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_285),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_392),
.B(n_409),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_389),
.B(n_396),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_426),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

INVxp33_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_407),
.B(n_352),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_426),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_409),
.B(n_411),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_382),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_414),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_395),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_409),
.B(n_286),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_390),
.B(n_289),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_424),
.B(n_291),
.C(n_290),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_420),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_412),
.B(n_294),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_463),
.B(n_419),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_432),
.B(n_419),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_431),
.B(n_422),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_434),
.B(n_422),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_469),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_432),
.B(n_421),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_444),
.A2(n_399),
.B1(n_427),
.B2(n_299),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_481),
.A2(n_399),
.B(n_427),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_298),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

AO22x1_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_310),
.B1(n_313),
.B2(n_305),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_318),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_433),
.B(n_319),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_480),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_475),
.B(n_320),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_479),
.B(n_321),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_472),
.B(n_323),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_443),
.B(n_325),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_429),
.B(n_326),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_446),
.B(n_329),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_459),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_430),
.B(n_316),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_454),
.B(n_458),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_488),
.B(n_48),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_488),
.B(n_49),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_457),
.A2(n_52),
.B1(n_53),
.B2(n_51),
.Y(n_524)
);

O2A1O1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_459),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_470),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_470),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_54),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_492),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_494),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_56),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_455),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_469),
.B(n_58),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_489),
.B(n_59),
.Y(n_535)
);

AND3x1_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_4),
.C(n_5),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_6),
.C(n_7),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_487),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_430),
.B(n_8),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_489),
.B(n_8),
.C(n_9),
.Y(n_541)
);

A2O1A1Ixp33_ASAP7_75t_L g542 ( 
.A1(n_456),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_455),
.B(n_10),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_477),
.B(n_60),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_61),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_487),
.B(n_62),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_471),
.B(n_63),
.Y(n_547)
);

AND2x6_ASAP7_75t_SL g548 ( 
.A(n_465),
.B(n_11),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_435),
.B(n_64),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_495),
.B(n_453),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_471),
.B(n_65),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_442),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_490),
.B(n_12),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_437),
.B(n_12),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_482),
.B(n_13),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_66),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_SL g561 ( 
.A(n_483),
.B(n_461),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_468),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_495),
.A2(n_467),
.B1(n_466),
.B2(n_463),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_473),
.B(n_68),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_492),
.B(n_69),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_482),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_491),
.B(n_13),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_553),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_511),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_550),
.A2(n_448),
.B1(n_466),
.B2(n_463),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_463),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_500),
.B(n_463),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_565),
.A2(n_492),
.B1(n_474),
.B2(n_448),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_540),
.A2(n_462),
.B(n_445),
.C(n_440),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_501),
.B(n_445),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_534),
.A2(n_523),
.B(n_522),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_506),
.Y(n_578)
);

INVx8_ASAP7_75t_L g579 ( 
.A(n_529),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_L g580 ( 
.A1(n_540),
.A2(n_486),
.B(n_484),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_518),
.A2(n_491),
.B1(n_494),
.B2(n_483),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_508),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_550),
.A2(n_491),
.B1(n_441),
.B2(n_449),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_563),
.A2(n_483),
.B1(n_494),
.B2(n_461),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_522),
.A2(n_461),
.B(n_494),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_510),
.A2(n_461),
.B1(n_441),
.B2(n_449),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_523),
.A2(n_464),
.B(n_71),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_521),
.A2(n_464),
.B(n_72),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_504),
.B(n_436),
.C(n_15),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_532),
.A2(n_464),
.B(n_74),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_516),
.B(n_16),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_526),
.B(n_70),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_565),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_559),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_527),
.B(n_75),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_547),
.A2(n_77),
.B(n_76),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_506),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_SL g601 ( 
.A1(n_535),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_551),
.A2(n_79),
.B(n_78),
.Y(n_602)
);

AOI21x1_ASAP7_75t_L g603 ( 
.A1(n_539),
.A2(n_81),
.B(n_80),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_533),
.B(n_82),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_497),
.B(n_17),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_567),
.A2(n_84),
.B(n_83),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_505),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_514),
.A2(n_88),
.B(n_87),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_513),
.A2(n_90),
.B(n_89),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_556),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_SL g611 ( 
.A1(n_549),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_557),
.A2(n_92),
.B(n_91),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_498),
.B(n_22),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_528),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_517),
.A2(n_94),
.B(n_93),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_552),
.A2(n_97),
.B(n_96),
.Y(n_616)
);

INVx11_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_542),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_546),
.A2(n_99),
.B(n_98),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_566),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_23),
.Y(n_622)
);

BUFx12f_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_560),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_544),
.A2(n_103),
.B(n_102),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_558),
.Y(n_626)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_104),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_507),
.B(n_24),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_499),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_503),
.B(n_105),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_604),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_621),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_629),
.B(n_559),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_586),
.A2(n_545),
.B(n_538),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_597),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_577),
.A2(n_525),
.B(n_554),
.Y(n_636)
);

AOI21xp33_ASAP7_75t_L g637 ( 
.A1(n_605),
.A2(n_496),
.B(n_541),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_576),
.B(n_530),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_583),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_620),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_578),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_572),
.A2(n_564),
.B(n_549),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_573),
.A2(n_524),
.A3(n_562),
.B(n_531),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_L g644 ( 
.A(n_584),
.B(n_520),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_585),
.A2(n_564),
.B(n_561),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_588),
.A2(n_531),
.B(n_512),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_592),
.A2(n_515),
.B(n_543),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_593),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_594),
.B(n_536),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_600),
.A2(n_530),
.B(n_529),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_630),
.A2(n_529),
.B(n_568),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_575),
.A2(n_568),
.B(n_537),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_612),
.A2(n_537),
.B(n_108),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_595),
.A2(n_109),
.B(n_106),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_624),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_571),
.A2(n_548),
.B(n_111),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_25),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_574),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_590),
.A2(n_603),
.B(n_616),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_619),
.A2(n_112),
.B(n_110),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_591),
.A2(n_606),
.B(n_613),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_596),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_604),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_579),
.A2(n_114),
.B(n_113),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_626),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_622),
.B(n_574),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_589),
.B(n_26),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_598),
.B(n_115),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_579),
.A2(n_118),
.B(n_117),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_627),
.B(n_120),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_620),
.Y(n_674)
);

NAND2x1_ASAP7_75t_L g675 ( 
.A(n_609),
.B(n_121),
.Y(n_675)
);

AOI221x1_ASAP7_75t_L g676 ( 
.A1(n_628),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_599),
.A2(n_124),
.B(n_123),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_587),
.B(n_29),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_607),
.B(n_126),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_610),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_611),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_624),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_579),
.B(n_581),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_617),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_602),
.B(n_128),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_608),
.A2(n_189),
.B(n_271),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_569),
.B(n_615),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_582),
.A2(n_625),
.B(n_569),
.C(n_601),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_623),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_610),
.A2(n_193),
.B(n_270),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_642),
.A2(n_190),
.B(n_269),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_684),
.B(n_131),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_646),
.A2(n_188),
.B(n_267),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_668),
.B(n_33),
.Y(n_694)
);

OAI321xp33_ASAP7_75t_L g695 ( 
.A1(n_689),
.A2(n_33),
.A3(n_34),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_632),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_639),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_658),
.A2(n_659),
.B1(n_649),
.B2(n_663),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_631),
.B(n_132),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_667),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_657),
.A2(n_665),
.B1(n_663),
.B2(n_689),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_648),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_650),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_635),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_633),
.B(n_657),
.Y(n_705)
);

O2A1O1Ixp5_ASAP7_75t_SL g706 ( 
.A1(n_637),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_631),
.B(n_272),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_638),
.B(n_38),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_679),
.B(n_133),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_659),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_631),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_648),
.B(n_42),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_660),
.B(n_669),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_651),
.A2(n_198),
.B(n_264),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_641),
.Y(n_716)
);

INVx3_ASAP7_75t_SL g717 ( 
.A(n_656),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_638),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_665),
.B(n_43),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_641),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_685),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_654),
.A2(n_200),
.B(n_263),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_682),
.B(n_640),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_652),
.A2(n_199),
.B(n_262),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_678),
.B(n_46),
.Y(n_726)
);

INVx3_ASAP7_75t_SL g727 ( 
.A(n_685),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_637),
.B(n_47),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_675),
.A2(n_135),
.B(n_139),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_683),
.A2(n_140),
.B(n_141),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_681),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_683),
.A2(n_143),
.B(n_144),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_664),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_SL g736 ( 
.A(n_666),
.B(n_149),
.Y(n_736)
);

NOR2x1_ASAP7_75t_SL g737 ( 
.A(n_673),
.B(n_150),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_644),
.B(n_266),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_670),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_690),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_653),
.B(n_151),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_697),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_704),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_716),
.B(n_720),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_705),
.A2(n_636),
.B1(n_671),
.B2(n_670),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_727),
.A2(n_688),
.B1(n_687),
.B2(n_673),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_720),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_721),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_698),
.B(n_687),
.Y(n_749)
);

NOR2x1_ASAP7_75t_R g750 ( 
.A(n_696),
.B(n_680),
.Y(n_750)
);

CKINVDCx11_ASAP7_75t_R g751 ( 
.A(n_717),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_719),
.A2(n_676),
.B1(n_647),
.B2(n_686),
.Y(n_752)
);

OAI21x1_ASAP7_75t_SL g753 ( 
.A1(n_737),
.A2(n_723),
.B(n_722),
.Y(n_753)
);

BUFx8_ASAP7_75t_L g754 ( 
.A(n_732),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_701),
.A2(n_686),
.B1(n_677),
.B2(n_662),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_696),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_703),
.Y(n_757)
);

NAND2x1p5_ASAP7_75t_L g758 ( 
.A(n_736),
.B(n_655),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_704),
.B(n_153),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_694),
.B(n_643),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_731),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_698),
.A2(n_645),
.B1(n_643),
.B2(n_661),
.Y(n_762)
);

AO21x1_ASAP7_75t_SL g763 ( 
.A1(n_722),
.A2(n_643),
.B(n_634),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_728),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_718),
.A2(n_261),
.B1(n_159),
.B2(n_160),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_720),
.Y(n_766)
);

CKINVDCx6p67_ASAP7_75t_R g767 ( 
.A(n_692),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_733),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_700),
.Y(n_769)
);

CKINVDCx11_ASAP7_75t_R g770 ( 
.A(n_721),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_715),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_709),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_713),
.B(n_163),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_714),
.A2(n_164),
.B(n_165),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_707),
.B(n_166),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_739),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_719),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_708),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_693),
.A2(n_173),
.B(n_174),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_692),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_709),
.A2(n_710),
.B1(n_711),
.B2(n_726),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_707),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_709),
.B(n_175),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_176),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_709),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_738),
.B(n_260),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_741),
.A2(n_181),
.B(n_182),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_740),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_699),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_695),
.A2(n_183),
.B1(n_186),
.B2(n_194),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_735),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_724),
.B(n_201),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_735),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_730),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_734),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_725),
.A2(n_208),
.B(n_211),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_691),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_729),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_706),
.Y(n_800)
);

NAND2x1_ASAP7_75t_L g801 ( 
.A(n_736),
.B(n_212),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_782),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_761),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_760),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_777),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_768),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_757),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_762),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_742),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_749),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_769),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_789),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_753),
.A2(n_257),
.B(n_219),
.Y(n_813)
);

AO21x2_ASAP7_75t_L g814 ( 
.A1(n_798),
.A2(n_255),
.B(n_220),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_796),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_779),
.Y(n_816)
);

AO21x2_ASAP7_75t_L g817 ( 
.A1(n_798),
.A2(n_253),
.B(n_221),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_800),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_789),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_789),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_797),
.A2(n_218),
.B(n_222),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_789),
.B(n_223),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_758),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_746),
.B(n_224),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_773),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_763),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_747),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_799),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_799),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_747),
.B(n_252),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_771),
.Y(n_831)
);

AO21x2_ASAP7_75t_L g832 ( 
.A1(n_788),
.A2(n_225),
.B(n_226),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_752),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_744),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_752),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_744),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_783),
.B(n_227),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_745),
.B(n_229),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_758),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_775),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_230),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_755),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_748),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_784),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_766),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_815),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_804),
.B(n_782),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_815),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_823),
.B(n_776),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_810),
.B(n_743),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_804),
.B(n_774),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_827),
.Y(n_855)
);

AO31x2_ASAP7_75t_L g856 ( 
.A1(n_808),
.A2(n_833),
.A3(n_835),
.B(n_843),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_803),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_804),
.B(n_767),
.Y(n_858)
);

AO21x2_ASAP7_75t_L g859 ( 
.A1(n_841),
.A2(n_794),
.B(n_792),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_803),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_828),
.B(n_781),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_SL g862 ( 
.A(n_842),
.B(n_756),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_824),
.A2(n_791),
.B1(n_778),
.B2(n_764),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_828),
.B(n_759),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_833),
.B(n_772),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_823),
.B(n_776),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

BUFx2_ASAP7_75t_SL g868 ( 
.A(n_812),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_835),
.B(n_786),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_790),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_802),
.A2(n_791),
.B1(n_772),
.B2(n_786),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_808),
.A2(n_765),
.B(n_795),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_810),
.B(n_764),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_807),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_829),
.Y(n_875)
);

AOI33xp33_ASAP7_75t_L g876 ( 
.A1(n_816),
.A2(n_778),
.A3(n_765),
.B1(n_795),
.B2(n_785),
.B3(n_793),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_808),
.B(n_843),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_812),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_812),
.B(n_751),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_806),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_829),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_844),
.B(n_787),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_823),
.B(n_801),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_827),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_844),
.B(n_770),
.Y(n_885)
);

INVx2_ASAP7_75t_R g886 ( 
.A(n_839),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_809),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_R g888 ( 
.A(n_834),
.B(n_750),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_805),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_824),
.A2(n_754),
.B1(n_232),
.B2(n_233),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_805),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_824),
.A2(n_754),
.B1(n_234),
.B2(n_236),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_823),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_826),
.B(n_231),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_826),
.B(n_237),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_853),
.B(n_847),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_SL g897 ( 
.A1(n_890),
.A2(n_842),
.B(n_838),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_867),
.B(n_826),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_863),
.B(n_847),
.C(n_838),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_SL g900 ( 
.A1(n_876),
.A2(n_824),
.B(n_816),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_892),
.B(n_822),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_871),
.B(n_824),
.C(n_839),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_861),
.A2(n_822),
.B1(n_826),
.B2(n_837),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_864),
.B(n_825),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_864),
.B(n_825),
.Y(n_905)
);

OA21x2_ASAP7_75t_L g906 ( 
.A1(n_849),
.A2(n_841),
.B(n_840),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_861),
.A2(n_822),
.B1(n_826),
.B2(n_837),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_850),
.B(n_825),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_850),
.B(n_805),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_885),
.B(n_834),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_862),
.B(n_846),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_855),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_SL g913 ( 
.A1(n_865),
.A2(n_822),
.B(n_837),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_882),
.B(n_811),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_882),
.B(n_811),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_867),
.B(n_826),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_865),
.A2(n_837),
.B1(n_836),
.B2(n_819),
.Y(n_917)
);

AND2x2_ASAP7_75t_SL g918 ( 
.A(n_872),
.B(n_830),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_874),
.B(n_819),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_869),
.A2(n_820),
.B1(n_848),
.B2(n_812),
.Y(n_920)
);

OA21x2_ASAP7_75t_L g921 ( 
.A1(n_849),
.A2(n_840),
.B(n_818),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_858),
.B(n_848),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_854),
.B(n_846),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_SL g924 ( 
.A1(n_869),
.A2(n_832),
.B1(n_813),
.B2(n_817),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_854),
.B(n_846),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_874),
.B(n_820),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_914),
.B(n_915),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_921),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_921),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_921),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_908),
.B(n_904),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_886),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_910),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_906),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_919),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_919),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_918),
.B(n_886),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_898),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_918),
.B(n_886),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_906),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_898),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_906),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_916),
.B(n_884),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_916),
.B(n_856),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_926),
.B(n_856),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_926),
.B(n_856),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_899),
.B(n_858),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_905),
.B(n_856),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_922),
.B(n_856),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_923),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_925),
.B(n_893),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_947),
.B(n_922),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_930),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_927),
.B(n_949),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_935),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_937),
.B(n_901),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_927),
.B(n_909),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_931),
.B(n_896),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_932),
.B(n_937),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_936),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_933),
.B(n_920),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_948),
.A2(n_900),
.B(n_902),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_931),
.B(n_897),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_933),
.B(n_893),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_932),
.B(n_924),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_948),
.B(n_880),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_953),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_956),
.B(n_944),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_956),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_953),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_964),
.Y(n_971)
);

NOR2x2_ASAP7_75t_L g972 ( 
.A(n_963),
.B(n_879),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_962),
.A2(n_911),
.B(n_813),
.C(n_832),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_958),
.B(n_949),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_957),
.B(n_950),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_963),
.B(n_945),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_954),
.B(n_950),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_955),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_960),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_969),
.A2(n_952),
.B1(n_965),
.B2(n_961),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_967),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_971),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_968),
.B(n_959),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_972),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_973),
.B(n_911),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_981),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_985),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_984),
.Y(n_989)
);

OAI222xp33_ASAP7_75t_L g990 ( 
.A1(n_986),
.A2(n_973),
.B1(n_976),
.B2(n_965),
.C1(n_978),
.C2(n_979),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_986),
.A2(n_976),
.B(n_939),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_988),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_987),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_987),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_988),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_989),
.Y(n_996)
);

NOR4xp75_ASAP7_75t_L g997 ( 
.A(n_995),
.B(n_991),
.C(n_980),
.D(n_985),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_996),
.B(n_989),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_995),
.B(n_985),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_992),
.B(n_983),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_993),
.A2(n_990),
.B(n_982),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_994),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_995),
.A2(n_939),
.B(n_975),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_959),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_1001),
.B(n_888),
.C(n_895),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_1000),
.B(n_894),
.C(n_895),
.Y(n_1007)
);

NOR3x1_ASAP7_75t_L g1008 ( 
.A(n_1003),
.B(n_1002),
.C(n_997),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_998),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_1006),
.B(n_894),
.C(n_974),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1004),
.B(n_977),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1009),
.B(n_966),
.Y(n_1012)
);

NAND4xp75_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_830),
.C(n_944),
.D(n_938),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_SL g1014 ( 
.A(n_1005),
.B(n_913),
.C(n_907),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_SL g1015 ( 
.A1(n_1007),
.A2(n_938),
.B(n_941),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_SL g1016 ( 
.A(n_1004),
.B(n_868),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1004),
.B(n_946),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1015),
.Y(n_1018)
);

OAI211xp5_ASAP7_75t_L g1019 ( 
.A1(n_1011),
.A2(n_930),
.B(n_872),
.C(n_845),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_1013),
.A2(n_813),
.B1(n_941),
.B2(n_903),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1012),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1017),
.A2(n_934),
.B1(n_940),
.B2(n_942),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1010),
.A2(n_813),
.B1(n_946),
.B2(n_945),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1016),
.A2(n_832),
.B1(n_951),
.B2(n_943),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1014),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_1011),
.A2(n_934),
.B1(n_942),
.B2(n_940),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1011),
.B(n_845),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1013),
.A2(n_832),
.B1(n_951),
.B2(n_943),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1013),
.A2(n_929),
.B1(n_928),
.B2(n_951),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_1011),
.Y(n_1030)
);

AND3x1_ASAP7_75t_L g1031 ( 
.A(n_1011),
.B(n_845),
.C(n_929),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_1011),
.B(n_951),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1013),
.A2(n_859),
.B1(n_928),
.B2(n_883),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_SL g1034 ( 
.A(n_1025),
.B(n_917),
.C(n_870),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1030),
.B(n_881),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_1021),
.B(n_821),
.C(n_883),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_1027),
.B(n_818),
.C(n_242),
.Y(n_1037)
);

NAND4xp75_ASAP7_75t_L g1038 ( 
.A(n_1018),
.B(n_872),
.C(n_873),
.D(n_877),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_1032),
.B(n_883),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_1028),
.B(n_873),
.C(n_817),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1041)
);

NAND4xp25_ASAP7_75t_L g1042 ( 
.A(n_1020),
.B(n_852),
.C(n_866),
.D(n_877),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1031),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1033),
.A2(n_875),
.B(n_881),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1023),
.B(n_875),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1029),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_SL g1047 ( 
.A(n_1024),
.B(n_817),
.C(n_814),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_1022),
.B(n_878),
.C(n_831),
.Y(n_1048)
);

OAI31xp33_ASAP7_75t_L g1049 ( 
.A1(n_1025),
.A2(n_866),
.A3(n_852),
.B(n_817),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_1018),
.B(n_239),
.Y(n_1050)
);

NAND4xp75_ASAP7_75t_L g1051 ( 
.A(n_1025),
.B(n_872),
.C(n_814),
.D(n_851),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1046),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1043),
.Y(n_1053)
);

AND3x4_ASAP7_75t_L g1054 ( 
.A(n_1050),
.B(n_866),
.C(n_852),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_1041),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1035),
.Y(n_1056)
);

AO22x2_ASAP7_75t_L g1057 ( 
.A1(n_1038),
.A2(n_868),
.B1(n_893),
.B2(n_814),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1034),
.B(n_860),
.Y(n_1058)
);

XOR2xp5_ASAP7_75t_L g1059 ( 
.A(n_1042),
.B(n_246),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1044),
.A2(n_821),
.B(n_831),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_1045),
.Y(n_1061)
);

NAND4xp75_ASAP7_75t_L g1062 ( 
.A(n_1049),
.B(n_814),
.C(n_248),
.D(n_250),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_1052),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1055),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1053),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_1059),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1054),
.A2(n_1037),
.B1(n_1039),
.B2(n_1048),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1061),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1064),
.B(n_1056),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_1062),
.C(n_1040),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1063),
.A2(n_1047),
.B(n_1058),
.C(n_1036),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1065),
.B(n_1060),
.C(n_1057),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_1069),
.A2(n_1066),
.B(n_1067),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_1051),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1074),
.A2(n_1071),
.B(n_1072),
.C(n_1073),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_247),
.B(n_251),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_878),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1075),
.A2(n_840),
.B(n_859),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_859),
.B(n_831),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_1076),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1079),
.A2(n_878),
.B(n_851),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1080),
.A2(n_878),
.B1(n_887),
.B2(n_889),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_R g1083 ( 
.A1(n_1082),
.A2(n_1081),
.B1(n_878),
.B2(n_891),
.C(n_857),
.Y(n_1083)
);

AOI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_887),
.B(n_889),
.C(n_860),
.Y(n_1084)
);


endmodule