module fake_jpeg_18651_n_284 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_51),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_39),
.C(n_42),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_42),
.C(n_41),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_18),
.Y(n_58)
);

NAND2x1p5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_21),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_44),
.B1(n_36),
.B2(n_40),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_38),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_70),
.C(n_75),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_22),
.B(n_40),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_39),
.B1(n_35),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_71),
.B1(n_87),
.B2(n_96),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_38),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_28),
.B1(n_34),
.B2(n_25),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_44),
.B1(n_40),
.B2(n_36),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_101),
.B1(n_42),
.B2(n_41),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.B(n_35),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_84),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_27),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_35),
.B1(n_33),
.B2(n_36),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_23),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_99),
.B1(n_42),
.B2(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_18),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_36),
.B1(n_44),
.B2(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_44),
.B1(n_27),
.B2(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_60),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_44),
.B1(n_29),
.B2(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_95),
.B1(n_71),
.B2(n_91),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_114),
.B(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_21),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_64),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_41),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_86),
.B(n_80),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_137),
.B(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_135),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_79),
.B1(n_86),
.B2(n_66),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_143),
.B1(n_145),
.B2(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_89),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_76),
.B1(n_65),
.B2(n_70),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_116),
.B(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_70),
.C(n_67),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_111),
.C(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_105),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_75),
.B1(n_63),
.B2(n_91),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_156),
.B1(n_122),
.B2(n_34),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_75),
.B1(n_83),
.B2(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_167),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_107),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_168),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_116),
.B1(n_88),
.B2(n_121),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_114),
.B1(n_112),
.B2(n_125),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_114),
.C(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_136),
.B1(n_142),
.B2(n_139),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_115),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_112),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_172),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_108),
.B1(n_105),
.B2(n_103),
.Y(n_172)
);

CKINVDCx10_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_180),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_155),
.B1(n_154),
.B2(n_147),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_176),
.B1(n_175),
.B2(n_171),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_28),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_143),
.B1(n_134),
.B2(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_25),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_149),
.B1(n_144),
.B2(n_140),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_151),
.B1(n_133),
.B2(n_32),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_197),
.B1(n_205),
.B2(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_196),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_16),
.B1(n_1),
.B2(n_4),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_176),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_19),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_157),
.C(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_220),
.C(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_197),
.B1(n_192),
.B2(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_160),
.B1(n_159),
.B2(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_221),
.B1(n_189),
.B2(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_159),
.C(n_165),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_32),
.B1(n_19),
.B2(n_24),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_32),
.C(n_24),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_206),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_32),
.B1(n_17),
.B2(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_24),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_214),
.A2(n_201),
.B1(n_196),
.B2(n_195),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_215),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_185),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_214),
.A2(n_217),
.B1(n_190),
.B2(n_202),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_244),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_226),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_224),
.B(n_219),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_230),
.B(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_217),
.B1(n_222),
.B2(n_223),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_188),
.B(n_209),
.C(n_207),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_232),
.B(n_6),
.C(n_9),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_4),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_237),
.C(n_234),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_249),
.B(n_10),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_249),
.B1(n_6),
.B2(n_10),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_17),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_248),
.C(n_247),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_264),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_247),
.C(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_249),
.CI(n_6),
.CON(n_267),
.SN(n_267)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_258),
.B(n_11),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_258),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_273),
.Y(n_276)
);

AOI31xp67_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_274),
.A3(n_268),
.B(n_267),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_263),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_267),
.Y(n_277)
);

NAND4xp25_ASAP7_75t_SL g278 ( 
.A(n_276),
.B(n_262),
.C(n_266),
.D(n_13),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_5),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_281),
.B(n_12),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_266),
.B(n_17),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_13),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_14),
.C(n_15),
.Y(n_284)
);


endmodule