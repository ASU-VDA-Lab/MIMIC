module fake_netlist_6_2350_n_88 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_88);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_88;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_86;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

AND2x2_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_9),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_0),
.B(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_5),
.A2(n_17),
.B1(n_14),
.B2(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_4),
.B1(n_2),
.B2(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2x1p5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp67_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_3),
.Y(n_47)
);

NOR2x1p5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_5),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_26),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

OAI21x1_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_31),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_33),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_6),
.B(n_34),
.C(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI21x1_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_34),
.B(n_43),
.Y(n_57)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.Y(n_58)
);

AO21x2_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_43),
.B(n_40),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_39),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_38),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_44),
.A3(n_53),
.B1(n_65),
.B2(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_61),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_51),
.B(n_40),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_44),
.B(n_55),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_53),
.C(n_54),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_73),
.C(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_77),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_61),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_86),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_84),
.B(n_85),
.Y(n_88)
);


endmodule