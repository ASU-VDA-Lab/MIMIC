module fake_jpeg_889_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_0),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_64),
.B1(n_60),
.B2(n_72),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_80),
.B1(n_69),
.B2(n_73),
.Y(n_113)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_72),
.B(n_64),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_59),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_62),
.C(n_84),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.C(n_61),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_53),
.B(n_65),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_80),
.B1(n_73),
.B2(n_69),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_93),
.B1(n_70),
.B2(n_55),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_86),
.B1(n_53),
.B2(n_65),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_125),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_90),
.B1(n_89),
.B2(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_67),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_131),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_90),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_63),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_51),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_104),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_148),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_49),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_68),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_54),
.B1(n_68),
.B2(n_75),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_3),
.B(n_5),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_54),
.B(n_75),
.C(n_24),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_155),
.B(n_28),
.C(n_43),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_119),
.B(n_131),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_158),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_1),
.B(n_2),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_159),
.B(n_2),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_1),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_142),
.B1(n_137),
.B2(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.C(n_172),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AO221x1_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_152),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_25),
.C(n_47),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_30),
.B1(n_41),
.B2(n_39),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_27),
.B(n_42),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_172),
.B1(n_168),
.B2(n_177),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_151),
.B1(n_157),
.B2(n_152),
.C(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_181),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_152),
.B(n_156),
.C(n_32),
.D(n_35),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_187),
.B(n_188),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_13),
.B1(n_18),
.B2(n_20),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_178),
.B(n_174),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_163),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_162),
.C(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_173),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_197),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_196),
.B(n_177),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_177),
.B(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_199),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_182),
.B1(n_189),
.B2(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_201),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_194),
.B1(n_191),
.B2(n_37),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_23),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_203),
.A3(n_198),
.B1(n_36),
.B2(n_26),
.C1(n_38),
.C2(n_48),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_208),
.B1(n_205),
.B2(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_21),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_22),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_22),
.B(n_23),
.Y(n_213)
);


endmodule