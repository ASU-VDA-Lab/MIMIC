module fake_jpeg_25844_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_73),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_1),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_52),
.B1(n_47),
.B2(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_86),
.B1(n_48),
.B2(n_65),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_52),
.B1(n_56),
.B2(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_66),
.B(n_68),
.C(n_49),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_3),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_88),
.B1(n_56),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_79),
.B1(n_63),
.B2(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_62),
.B1(n_54),
.B2(n_59),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_48),
.B1(n_65),
.B2(n_63),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_69),
.B1(n_63),
.B2(n_64),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_60),
.B1(n_51),
.B2(n_67),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_60),
.B1(n_51),
.B2(n_67),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_102),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_85),
.B1(n_25),
.B2(n_26),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_20),
.B1(n_44),
.B2(n_43),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_7),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_4),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_92),
.C(n_6),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_97),
.C(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_110),
.B1(n_111),
.B2(n_103),
.Y(n_127)
);

INVxp33_ASAP7_75t_SL g126 ( 
.A(n_124),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_129),
.Y(n_141)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_114),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_110),
.B1(n_99),
.B2(n_93),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_136),
.B1(n_139),
.B2(n_9),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_99),
.B1(n_103),
.B2(n_10),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_138),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_8),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_28),
.C(n_39),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_150),
.C(n_128),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.C(n_146),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_140),
.C(n_137),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_145),
.C(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_159),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_130),
.Y(n_161)
);

OAI311xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_149),
.A3(n_18),
.B1(n_19),
.C1(n_30),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_15),
.B(n_33),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_34),
.Y(n_165)
);


endmodule