module fake_jpeg_5832_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_20),
.CON(n_43),
.SN(n_43)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_50),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_53),
.Y(n_87)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_19),
.B1(n_28),
.B2(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_45),
.B1(n_65),
.B2(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_19),
.B1(n_42),
.B2(n_28),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_83),
.B1(n_42),
.B2(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_39),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_24),
.B(n_26),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_34),
.B1(n_28),
.B2(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_21),
.Y(n_110)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_38),
.B1(n_45),
.B2(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_104),
.B1(n_101),
.B2(n_41),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_34),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_86),
.C(n_21),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_38),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_37),
.C(n_44),
.Y(n_131)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_102),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_110),
.Y(n_133)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_111),
.B1(n_116),
.B2(n_121),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_55),
.B1(n_53),
.B2(n_48),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_115),
.Y(n_147)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_48),
.B1(n_27),
.B2(n_26),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_76),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_29),
.Y(n_126)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_10),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_127),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_74),
.B(n_80),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_38),
.B(n_121),
.Y(n_170)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_137),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_83),
.B(n_37),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_148),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_38),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_127),
.B1(n_148),
.B2(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_146),
.C(n_107),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_93),
.Y(n_139)
);

CKINVDCx10_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_93),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_38),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_86),
.C(n_41),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_23),
.B(n_38),
.C(n_21),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_165),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_114),
.C(n_118),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_155),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_132),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_117),
.B1(n_44),
.B2(n_18),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_162),
.B1(n_167),
.B2(n_135),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_161),
.B(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_44),
.C(n_62),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_117),
.B1(n_17),
.B2(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_146),
.C(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_172),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_134),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_38),
.C(n_103),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_132),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_R g211 ( 
.A1(n_178),
.A2(n_151),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_155),
.C(n_176),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_122),
.B1(n_130),
.B2(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_133),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_103),
.B1(n_115),
.B2(n_106),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_193),
.B1(n_198),
.B2(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_126),
.B1(n_145),
.B2(n_40),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_134),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_119),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_203),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_134),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_124),
.B1(n_40),
.B2(n_25),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_40),
.B1(n_73),
.B2(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_1),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_40),
.B(n_22),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_22),
.B(n_32),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_23),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_224),
.C(n_202),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_160),
.B(n_153),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_218),
.B1(n_181),
.B2(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_211),
.A2(n_221),
.B1(n_191),
.B2(n_200),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_164),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_0),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_223),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_174),
.B1(n_21),
.B2(n_16),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_16),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_222),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_32),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_182),
.C(n_177),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_196),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_91),
.B1(n_73),
.B2(n_58),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_25),
.B1(n_56),
.B2(n_52),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_185),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_237),
.B(n_240),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_193),
.C(n_190),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_199),
.B1(n_198),
.B2(n_192),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_244),
.B1(n_248),
.B2(n_216),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_205),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_1),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_235),
.B(n_228),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_32),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_259),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_221),
.B(n_238),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_205),
.B1(n_226),
.B2(n_207),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_244),
.B1(n_245),
.B2(n_213),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_216),
.B1(n_204),
.B2(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_217),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_227),
.B(n_16),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_206),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_204),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_276),
.B(n_32),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_245),
.B1(n_248),
.B2(n_213),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_282),
.B1(n_257),
.B2(n_258),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_232),
.C(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_22),
.C(n_16),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_257),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_232),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_259),
.Y(n_290)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_73),
.B1(n_91),
.B2(n_52),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_32),
.B1(n_22),
.B2(n_3),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_253),
.B1(n_266),
.B2(n_262),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_289),
.B(n_293),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_275),
.B(n_274),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_279),
.B1(n_273),
.B2(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_296),
.B1(n_274),
.B2(n_8),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_281),
.C(n_2),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_278),
.B(n_8),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_23),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_8),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_302),
.B(n_4),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_16),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_306),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_7),
.Y(n_306)
);

NOR2x1_ASAP7_75t_R g307 ( 
.A(n_298),
.B(n_287),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_308),
.B(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_295),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_291),
.B1(n_284),
.B2(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_4),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_297),
.B(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_318),
.B(n_5),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.C(n_5),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_6),
.B(n_9),
.C(n_12),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_6),
.B(n_12),
.Y(n_324)
);

AOI211xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_6),
.B(n_12),
.C(n_13),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_1),
.Y(n_326)
);


endmodule