module fake_jpeg_30556_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_42),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_1),
.B(n_2),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_45),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_39),
.B(n_37),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_8),
.B(n_9),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_47),
.B1(n_43),
.B2(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_80),
.B1(n_82),
.B2(n_4),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_68),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_7),
.C(n_8),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_6),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_21),
.B1(n_32),
.B2(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_17),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_6),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_7),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_97),
.B1(n_22),
.B2(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_10),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_108),
.B1(n_88),
.B2(n_93),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_107),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_96),
.B1(n_89),
.B2(n_97),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_86),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_103),
.B(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_109),
.Y(n_114)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_113),
.B(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_105),
.C(n_102),
.Y(n_117)
);

AOI221xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_35),
.B1(n_25),
.B2(n_27),
.C(n_28),
.Y(n_118)
);


endmodule