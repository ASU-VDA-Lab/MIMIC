module fake_jpeg_1886_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_71),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_40),
.B2(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_44),
.B1(n_66),
.B2(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_51),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_40),
.B1(n_50),
.B2(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_84),
.B1(n_42),
.B2(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_78),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_50),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_42),
.B(n_47),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_43),
.B(n_36),
.C(n_48),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g80 ( 
.A(n_64),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_85),
.B1(n_79),
.B2(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_90),
.B1(n_103),
.B2(n_38),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_42),
.C(n_41),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_17),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_47),
.B1(n_38),
.B2(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_38),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_4),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_18),
.C(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_4),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_19),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_106),
.B(n_118),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_11),
.Y(n_143)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_121),
.B1(n_11),
.B2(n_10),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_8),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_28),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_133),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_136),
.C(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_129),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_128),
.B1(n_123),
.B2(n_146),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_130),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_124),
.C(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_15),
.C(n_16),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_23),
.Y(n_158)
);


endmodule