module fake_jpeg_6165_n_28 (n_3, n_2, n_1, n_0, n_4, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

AND2x6_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_9),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_13),
.B(n_10),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_21),
.Y(n_24)
);

AOI211xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_25),
.B(n_7),
.C(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

OAI21x1_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_8),
.B(n_12),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_8),
.Y(n_28)
);


endmodule