module fake_jpeg_19495_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_65),
.Y(n_87)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_34),
.B1(n_20),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_52),
.B1(n_56),
.B2(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_19),
.B1(n_20),
.B2(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_26),
.B1(n_16),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_22),
.B1(n_16),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_72),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_88),
.B1(n_97),
.B2(n_48),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_42),
.B1(n_38),
.B2(n_40),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_63),
.B1(n_45),
.B2(n_35),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_46),
.B1(n_42),
.B2(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_82),
.B1(n_103),
.B2(n_45),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_47),
.C(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_40),
.B1(n_38),
.B2(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_89),
.Y(n_127)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_48),
.B1(n_63),
.B2(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_111),
.B1(n_113),
.B2(n_122),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_120),
.B1(n_84),
.B2(n_33),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_45),
.B1(n_35),
.B2(n_43),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_45),
.B1(n_35),
.B2(n_57),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_88),
.B1(n_68),
.B2(n_79),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_18),
.CON(n_118),
.SN(n_118)
);

OAI211xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_91),
.B(n_102),
.C(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_78),
.B1(n_85),
.B2(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_18),
.B1(n_10),
.B2(n_15),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_101),
.B1(n_98),
.B2(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_99),
.B1(n_92),
.B2(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_95),
.B1(n_79),
.B2(n_76),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_139),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_76),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_113),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_141),
.B(n_146),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_83),
.B(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_110),
.B1(n_112),
.B2(n_131),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_12),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_13),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_70),
.B(n_75),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_150),
.B(n_163),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_107),
.A2(n_95),
.B1(n_33),
.B2(n_28),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_84),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_156),
.B1(n_160),
.B2(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_33),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_162),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_111),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_141),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_166),
.B(n_168),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_122),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_180),
.B1(n_185),
.B2(n_154),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_9),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_115),
.C(n_110),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_183),
.C(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_188),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_108),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_192),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_162),
.B1(n_133),
.B2(n_146),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_143),
.B1(n_142),
.B2(n_148),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_115),
.C(n_112),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_108),
.B(n_105),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_2),
.B(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_105),
.B1(n_27),
.B2(n_21),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_151),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_116),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_21),
.C(n_9),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_137),
.A2(n_0),
.B(n_2),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_201),
.B1(n_225),
.B2(n_182),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_163),
.B1(n_150),
.B2(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_161),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_204),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_9),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_15),
.C(n_8),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_218),
.C(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_172),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_187),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_2),
.B(n_4),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_197),
.B(n_181),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_11),
.C(n_14),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_175),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_11),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_15),
.C(n_8),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_165),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_193),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_231),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_248),
.B1(n_249),
.B2(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_197),
.B(n_173),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_222),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_171),
.B1(n_196),
.B2(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_219),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_230),
.B(n_206),
.C(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_205),
.C(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_266),
.C(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_227),
.B1(n_239),
.B2(n_242),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_218),
.B(n_194),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_255),
.B(n_228),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_207),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_186),
.B(n_195),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_210),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_248),
.B(n_205),
.CI(n_208),
.CON(n_262),
.SN(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_208),
.Y(n_264)
);

NOR2x1_ASAP7_75t_R g265 ( 
.A(n_234),
.B(n_190),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_168),
.C(n_212),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_236),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_279),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_268),
.B1(n_261),
.B2(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_237),
.C(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_224),
.C(n_255),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_229),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_229),
.B1(n_240),
.B2(n_231),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_283),
.B1(n_237),
.B2(n_228),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_233),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_256),
.B1(n_253),
.B2(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_288),
.B1(n_267),
.B2(n_245),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_268),
.B1(n_259),
.B2(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_278),
.Y(n_302)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_258),
.Y(n_291)
);

OAI21x1_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_294),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_281),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_277),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_267),
.C(n_238),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_235),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_299),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_269),
.B1(n_271),
.B2(n_170),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_285),
.B1(n_185),
.B2(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_289),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_293),
.C(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_298),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_316),
.B(n_317),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_305),
.C(n_301),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_309),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_314),
.Y(n_321)
);

OAI311xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_319),
.A3(n_300),
.B1(n_310),
.C1(n_274),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_243),
.C(n_10),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_12),
.C(n_13),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_5),
.C(n_6),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_5),
.Y(n_326)
);


endmodule