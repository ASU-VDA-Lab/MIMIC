module fake_jpeg_14291_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_28),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_113),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_20),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_83),
.B(n_108),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_105),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_95),
.Y(n_160)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_97),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_22),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_22),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_26),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_32),
.Y(n_138)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_28),
.B(n_9),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_122),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_19),
.Y(n_124)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_33),
.B1(n_52),
.B2(n_57),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_126),
.A2(n_199),
.B1(n_55),
.B2(n_97),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_65),
.A2(n_52),
.B1(n_19),
.B2(n_42),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_151),
.A2(n_176),
.B1(n_185),
.B2(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_44),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_23),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_161),
.B(n_173),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_83),
.A2(n_49),
.B1(n_19),
.B2(n_42),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_162),
.A2(n_178),
.B1(n_206),
.B2(n_170),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_23),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_107),
.B(n_31),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_52),
.B1(n_42),
.B2(n_43),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_82),
.A2(n_49),
.B1(n_43),
.B2(n_26),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_189),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_112),
.A2(n_43),
.B1(n_58),
.B2(n_57),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_106),
.B(n_25),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_74),
.B(n_58),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_74),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_64),
.B(n_25),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_202),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_62),
.A2(n_49),
.B1(n_55),
.B2(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_119),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_98),
.B(n_24),
.Y(n_202)
);

AO22x2_ASAP7_75t_L g205 ( 
.A1(n_63),
.A2(n_47),
.B1(n_26),
.B2(n_41),
.Y(n_205)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_32),
.B1(n_27),
.B2(n_41),
.Y(n_206)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_209),
.Y(n_316)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_210),
.Y(n_303)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_99),
.B1(n_102),
.B2(n_71),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_212),
.B(n_278),
.Y(n_295)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_213),
.Y(n_306)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_214),
.Y(n_310)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_152),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_217),
.B(n_237),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_178),
.B1(n_162),
.B2(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_218),
.A2(n_208),
.B1(n_220),
.B2(n_245),
.Y(n_291)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_220),
.Y(n_340)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_137),
.A2(n_34),
.B(n_47),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_224),
.B(n_234),
.C(n_251),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_146),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_127),
.Y(n_230)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_170),
.A2(n_34),
.B1(n_124),
.B2(n_67),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_231),
.Y(n_308)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_131),
.B(n_122),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_235),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_128),
.B(n_95),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_134),
.B(n_118),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_129),
.B(n_36),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_242),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_156),
.B(n_110),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_268),
.Y(n_286)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_240),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_133),
.A2(n_56),
.B(n_46),
.C(n_45),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_32),
.B1(n_24),
.B2(n_56),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_244),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_36),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_245),
.B(n_246),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_59),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_135),
.A2(n_87),
.B1(n_104),
.B2(n_103),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_247),
.A2(n_266),
.B1(n_267),
.B2(n_270),
.Y(n_326)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_163),
.Y(n_249)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_110),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_172),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_253),
.B(n_261),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_144),
.A2(n_132),
.B1(n_155),
.B2(n_139),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_254),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_149),
.Y(n_256)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_258),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_262),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_175),
.B(n_0),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_269),
.C(n_3),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_169),
.B(n_31),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_172),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_265),
.B(n_271),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_139),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_93),
.C(n_89),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_145),
.A2(n_84),
.B1(n_81),
.B2(n_77),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_181),
.B(n_40),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_141),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_274),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_154),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_154),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_181),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_143),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_143),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

BUFx6f_ASAP7_75t_SL g296 ( 
.A(n_279),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_141),
.Y(n_280)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_177),
.B(n_9),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_13),
.Y(n_333)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_282),
.Y(n_312)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_171),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_285),
.B(n_300),
.C(n_14),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_291),
.A2(n_307),
.B1(n_329),
.B2(n_255),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_229),
.A2(n_140),
.B1(n_200),
.B2(n_184),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_211),
.B(n_203),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_208),
.A2(n_203),
.B1(n_200),
.B2(n_150),
.Y(n_307)
);

AOI32xp33_ASAP7_75t_L g324 ( 
.A1(n_246),
.A2(n_166),
.A3(n_147),
.B1(n_184),
.B2(n_159),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_324),
.A2(n_224),
.B(n_269),
.C(n_235),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_273),
.A2(n_159),
.B1(n_150),
.B2(n_168),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_256),
.B1(n_240),
.B2(n_279),
.Y(n_347)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_218),
.A2(n_188),
.B1(n_187),
.B2(n_166),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_333),
.B(n_17),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_266),
.A2(n_188),
.B1(n_187),
.B2(n_147),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_235),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_273),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_0),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_338),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_222),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_3),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_238),
.B(n_229),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_260),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_251),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_216),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_359),
.B1(n_362),
.B2(n_372),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_227),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_357),
.C(n_286),
.Y(n_421)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_351),
.B(n_394),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_352),
.A2(n_389),
.B(n_392),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_342),
.Y(n_353)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_308),
.A2(n_210),
.B1(n_215),
.B2(n_268),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_354),
.Y(n_413)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_302),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_358),
.A2(n_361),
.B1(n_366),
.B2(n_368),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_291),
.A2(n_242),
.B1(n_282),
.B2(n_277),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_360),
.B(n_363),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_294),
.A2(n_235),
.B1(n_239),
.B2(n_233),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_283),
.B1(n_232),
.B2(n_230),
.Y(n_362)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_294),
.A2(n_239),
.B1(n_233),
.B2(n_260),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_294),
.A2(n_243),
.B1(n_251),
.B2(n_241),
.Y(n_368)
);

XOR2x2_ASAP7_75t_L g369 ( 
.A(n_293),
.B(n_221),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_340),
.Y(n_399)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_300),
.B(n_214),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_384),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_219),
.B1(n_223),
.B2(n_212),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_373),
.A2(n_374),
.B1(n_376),
.B2(n_297),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_301),
.A2(n_213),
.B1(n_226),
.B2(n_259),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_301),
.A2(n_250),
.B1(n_209),
.B2(n_257),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_385),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_280),
.B1(n_236),
.B2(n_5),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_378),
.A2(n_379),
.B1(n_380),
.B2(n_382),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_236),
.B1(n_14),
.B2(n_5),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_338),
.A2(n_11),
.B1(n_18),
.B2(n_5),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_381),
.B(n_386),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_326),
.A2(n_337),
.B1(n_284),
.B2(n_344),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_287),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_383),
.B(n_315),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_3),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_4),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_388),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_325),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_284),
.B(n_252),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_345),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_390)
);

OA22x2_ASAP7_75t_L g397 ( 
.A1(n_390),
.A2(n_379),
.B1(n_380),
.B2(n_378),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_318),
.B(n_252),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_391),
.B(n_393),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_SL g392 ( 
.A1(n_330),
.A2(n_11),
.B(n_14),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_331),
.B(n_15),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_284),
.B(n_15),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_395),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_304),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_437),
.C(n_421),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_434),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_399),
.B(n_401),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_383),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_414),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_340),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_309),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_402),
.B(n_406),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_374),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_382),
.A2(n_295),
.B1(n_308),
.B2(n_330),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_410),
.A2(n_424),
.B1(n_395),
.B2(n_376),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_364),
.A2(n_295),
.B(n_286),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_411),
.A2(n_428),
.B(n_430),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_389),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_356),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_418),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_365),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_401),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_358),
.A2(n_299),
.B1(n_286),
.B2(n_312),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_425),
.A2(n_317),
.B1(n_290),
.B2(n_296),
.Y(n_468)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_364),
.A2(n_297),
.B(n_314),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_348),
.A2(n_332),
.B(n_320),
.Y(n_430)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_431),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_339),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_389),
.A2(n_303),
.B(n_311),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_430),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_305),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_407),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_439),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_432),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_425),
.A2(n_366),
.B1(n_348),
.B2(n_361),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_441),
.A2(n_442),
.B1(n_448),
.B2(n_468),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_400),
.B1(n_368),
.B2(n_409),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_444),
.C(n_446),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_363),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_386),
.C(n_387),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_413),
.A2(n_352),
.B(n_367),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_447),
.A2(n_435),
.B(n_316),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_373),
.B1(n_388),
.B2(n_372),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_429),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_450),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_396),
.B(n_395),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_459),
.C(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_456),
.A2(n_463),
.B1(n_469),
.B2(n_470),
.Y(n_490)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_381),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_429),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_460),
.B(n_467),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_408),
.Y(n_462)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_381),
.B1(n_377),
.B2(n_355),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_393),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_472),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_385),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_422),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_413),
.A2(n_289),
.B1(n_317),
.B2(n_303),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_422),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_471),
.A2(n_475),
.B1(n_452),
.B2(n_461),
.Y(n_505)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_473),
.B(n_474),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_375),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_398),
.B(n_350),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_402),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_482),
.B(n_494),
.C(n_500),
.Y(n_514)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_410),
.B1(n_424),
.B2(n_411),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_484),
.A2(n_488),
.B1(n_498),
.B2(n_501),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_448),
.A2(n_428),
.B1(n_412),
.B2(n_397),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_496),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_447),
.A2(n_436),
.B(n_404),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_495),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_404),
.C(n_433),
.Y(n_494)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_462),
.B(n_397),
.CI(n_288),
.CON(n_495),
.SN(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_454),
.B(n_415),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_441),
.A2(n_438),
.B1(n_472),
.B2(n_449),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_497),
.A2(n_439),
.B(n_458),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_438),
.A2(n_397),
.B1(n_426),
.B2(n_418),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_416),
.C(n_334),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_460),
.B1(n_468),
.B2(n_474),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_456),
.A2(n_417),
.B1(n_416),
.B2(n_415),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_502),
.A2(n_510),
.B1(n_296),
.B2(n_341),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_454),
.B(n_444),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_507),
.Y(n_536)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_504),
.Y(n_511)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_505),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_506),
.A2(n_457),
.B(n_453),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_298),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_298),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_508),
.B(n_509),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_298),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_465),
.A2(n_435),
.B1(n_341),
.B2(n_328),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g513 ( 
.A1(n_481),
.A2(n_461),
.B(n_467),
.Y(n_513)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_513),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_464),
.C(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_521),
.C(n_531),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_455),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_516),
.B(n_522),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_519),
.A2(n_523),
.B(n_526),
.Y(n_548)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_478),
.Y(n_520)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_482),
.C(n_494),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_466),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_504),
.B(n_445),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_524),
.B(n_512),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_496),
.B(n_445),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_525),
.B(n_541),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_435),
.B(n_370),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_527),
.A2(n_495),
.B1(n_16),
.B2(n_18),
.Y(n_556)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_528),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_476),
.A2(n_498),
.B1(n_488),
.B2(n_484),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_509),
.B(n_316),
.C(n_323),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_499),
.B(n_323),
.Y(n_532)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_532),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_477),
.B(n_319),
.Y(n_533)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_479),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_538),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_479),
.A2(n_290),
.B(n_289),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_537),
.B(n_539),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_476),
.A2(n_501),
.B1(n_493),
.B2(n_491),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_506),
.A2(n_322),
.B(n_335),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_489),
.B(n_322),
.C(n_335),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_508),
.C(n_507),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_544),
.B(n_553),
.C(n_559),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_514),
.B(n_490),
.C(n_502),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_545),
.B(n_550),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_514),
.B(n_486),
.C(n_487),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_480),
.C(n_510),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_495),
.Y(n_555)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_517),
.A2(n_15),
.B(n_18),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_558),
.B(n_533),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_521),
.B(n_18),
.C(n_540),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_532),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_539),
.Y(n_575)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_562),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_563),
.B(n_567),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_511),
.B(n_528),
.Y(n_564)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_564),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_534),
.A2(n_535),
.B1(n_526),
.B2(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_565),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_529),
.B(n_531),
.C(n_522),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_566),
.B(n_544),
.C(n_543),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_536),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_551),
.A2(n_518),
.B1(n_523),
.B2(n_538),
.Y(n_568)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_568),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_515),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_569),
.B(n_585),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_542),
.A2(n_518),
.B1(n_519),
.B2(n_511),
.Y(n_570)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_570),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_571),
.B(n_586),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_581),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_548),
.A2(n_525),
.B(n_541),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_576),
.A2(n_558),
.B(n_578),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_548),
.A2(n_536),
.B(n_555),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_578),
.A2(n_557),
.B(n_549),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_564),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_546),
.B(n_552),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_584),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_552),
.B(n_554),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_566),
.B(n_550),
.C(n_545),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_567),
.Y(n_587)
);

XNOR2x1_ASAP7_75t_L g600 ( 
.A(n_587),
.B(n_547),
.Y(n_600)
);

AOI21x1_ASAP7_75t_L g619 ( 
.A1(n_591),
.A2(n_571),
.B(n_583),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_580),
.A2(n_542),
.B(n_565),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_594),
.A2(n_601),
.B(n_606),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_572),
.A2(n_554),
.B(n_561),
.Y(n_595)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_547),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_598),
.B(n_599),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_553),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_583),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_580),
.A2(n_561),
.B(n_556),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_569),
.B(n_559),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_602),
.B(n_604),
.Y(n_608)
);

XOR2x2_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_572),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_574),
.B(n_586),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_574),
.B(n_585),
.Y(n_605)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_605),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_575),
.A2(n_584),
.B(n_577),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_614),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_589),
.A2(n_579),
.B(n_576),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_611),
.A2(n_619),
.B(n_603),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_590),
.A2(n_597),
.B1(n_568),
.B2(n_573),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_616),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_573),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_591),
.A2(n_593),
.B1(n_606),
.B2(n_577),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_593),
.A2(n_570),
.B1(n_581),
.B2(n_582),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_617),
.B(n_618),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_600),
.B(n_587),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_620),
.B(n_598),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_621),
.A2(n_612),
.B(n_595),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_609),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_592),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_624),
.B(n_628),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_594),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_625),
.B(n_627),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_601),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_617),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_610),
.B(n_596),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_629),
.B(n_596),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_630),
.B(n_609),
.C(n_613),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_635),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_623),
.Y(n_634)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_634),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_637),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_633),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_641),
.B(n_630),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_638),
.Y(n_642)
);

OAI321xp33_ASAP7_75t_L g644 ( 
.A1(n_642),
.A2(n_643),
.A3(n_640),
.B1(n_632),
.B2(n_639),
.C(n_634),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_645),
.B(n_626),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_618),
.B(n_620),
.Y(n_647)
);


endmodule