module real_aes_15653_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_0), .A2(n_99), .B1(n_517), .B2(n_1203), .C(n_1206), .Y(n_1202) );
AOI22xp33_ASAP7_75t_SL g1220 ( .A1(n_0), .A2(n_201), .B1(n_1221), .B2(n_1223), .Y(n_1220) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1), .Y(n_1655) );
OAI211xp5_ASAP7_75t_L g1689 ( .A1(n_1), .A2(n_1194), .B(n_1690), .C(n_1695), .Y(n_1689) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_2), .A2(n_82), .B1(n_1446), .B2(n_1449), .Y(n_1471) );
INVx1_ASAP7_75t_L g1263 ( .A(n_3), .Y(n_1263) );
INVx1_ASAP7_75t_L g327 ( .A(n_4), .Y(n_327) );
AND2x2_ASAP7_75t_L g436 ( .A(n_4), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g465 ( .A(n_4), .B(n_216), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_4), .B(n_337), .Y(n_502) );
INVx1_ASAP7_75t_L g1149 ( .A(n_5), .Y(n_1149) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_5), .A2(n_10), .B1(n_485), .B2(n_1169), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_6), .A2(n_231), .B1(n_887), .B2(n_890), .Y(n_886) );
OAI22xp33_ASAP7_75t_L g918 ( .A1(n_6), .A2(n_231), .B1(n_919), .B2(n_922), .Y(n_918) );
INVx1_ASAP7_75t_L g1107 ( .A(n_7), .Y(n_1107) );
INVx1_ASAP7_75t_L g1192 ( .A(n_8), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1227 ( .A1(n_8), .A2(n_86), .B1(n_1228), .B2(n_1230), .Y(n_1227) );
INVx1_ASAP7_75t_L g1730 ( .A(n_9), .Y(n_1730) );
OA222x2_ASAP7_75t_L g1739 ( .A1(n_9), .A2(n_132), .B1(n_158), .B2(n_476), .C1(n_1740), .C2(n_1742), .Y(n_1739) );
INVx1_ASAP7_75t_L g1158 ( .A(n_10), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1679 ( .A1(n_11), .A2(n_149), .B1(n_1680), .B2(n_1682), .Y(n_1679) );
INVx1_ASAP7_75t_L g1691 ( .A(n_11), .Y(n_1691) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_12), .A2(n_303), .B1(n_362), .B2(n_367), .C(n_373), .Y(n_361) );
OAI21xp33_ASAP7_75t_SL g475 ( .A1(n_12), .A2(n_476), .B(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g879 ( .A(n_13), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_14), .A2(n_85), .B1(n_517), .B2(n_1051), .C(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_SL g1226 ( .A1(n_14), .A2(n_174), .B1(n_544), .B2(n_994), .Y(n_1226) );
INVx2_ASAP7_75t_L g357 ( .A(n_15), .Y(n_357) );
INVx1_ASAP7_75t_L g1262 ( .A(n_16), .Y(n_1262) );
OAI322xp33_ASAP7_75t_L g1266 ( .A1(n_16), .A2(n_1267), .A3(n_1272), .B1(n_1273), .B2(n_1276), .C1(n_1282), .C2(n_1284), .Y(n_1266) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_17), .Y(n_807) );
INVx1_ASAP7_75t_L g836 ( .A(n_18), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1724 ( .A1(n_19), .A2(n_160), .B1(n_1721), .B2(n_1725), .Y(n_1724) );
INVxp67_ASAP7_75t_SL g1756 ( .A(n_19), .Y(n_1756) );
AOI221xp5_ASAP7_75t_L g1256 ( .A1(n_20), .A2(n_200), .B1(n_657), .B2(n_1183), .C(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1275 ( .A(n_20), .Y(n_1275) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_21), .A2(n_254), .B1(n_407), .B2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g469 ( .A(n_21), .Y(n_469) );
INVx1_ASAP7_75t_L g1347 ( .A(n_22), .Y(n_1347) );
OAI211xp5_ASAP7_75t_L g874 ( .A1(n_23), .A2(n_824), .B(n_875), .C(n_878), .Y(n_874) );
INVx1_ASAP7_75t_L g917 ( .A(n_23), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_24), .A2(n_282), .B1(n_407), .B2(n_410), .Y(n_1108) );
INVxp67_ASAP7_75t_SL g1110 ( .A(n_24), .Y(n_1110) );
INVx1_ASAP7_75t_L g742 ( .A(n_25), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_25), .A2(n_130), .B1(n_768), .B2(n_770), .C(n_771), .Y(n_767) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_26), .Y(n_322) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_26), .B(n_320), .Y(n_1440) );
INVx1_ASAP7_75t_L g846 ( .A(n_27), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_28), .A2(n_193), .B1(n_562), .B2(n_564), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_28), .A2(n_265), .B1(n_610), .B2(n_613), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_29), .A2(n_264), .B1(n_962), .B2(n_1260), .Y(n_1259) );
INVxp67_ASAP7_75t_L g1271 ( .A(n_29), .Y(n_1271) );
INVx1_ASAP7_75t_L g1022 ( .A(n_30), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_30), .A2(n_59), .B1(n_749), .B2(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1237 ( .A(n_31), .Y(n_1237) );
OAI211xp5_ASAP7_75t_SL g1343 ( .A1(n_32), .A2(n_1344), .B(n_1346), .C(n_1349), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_32), .A2(n_239), .B1(n_989), .B2(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1100 ( .A(n_33), .Y(n_1100) );
INVx1_ASAP7_75t_L g755 ( .A(n_34), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_34), .A2(n_45), .B1(n_362), .B2(n_367), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_35), .A2(n_262), .B1(n_962), .B2(n_963), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_35), .A2(n_200), .B1(n_544), .B2(n_547), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_36), .A2(n_66), .B1(n_1439), .B2(n_1456), .Y(n_1470) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_37), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_37), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g1720 ( .A1(n_38), .A2(n_236), .B1(n_1219), .B2(n_1721), .Y(n_1720) );
INVxp67_ASAP7_75t_SL g1749 ( .A(n_38), .Y(n_1749) );
INVx1_ASAP7_75t_L g1310 ( .A(n_39), .Y(n_1310) );
INVx1_ASAP7_75t_L g1671 ( .A(n_40), .Y(n_1671) );
AOI21xp33_ASAP7_75t_L g1696 ( .A1(n_40), .A2(n_655), .B(n_658), .Y(n_1696) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_41), .A2(n_386), .B1(n_794), .B2(n_797), .Y(n_793) );
INVx1_ASAP7_75t_L g814 ( .A(n_41), .Y(n_814) );
INVx1_ASAP7_75t_L g1307 ( .A(n_42), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1330 ( .A1(n_42), .A2(n_230), .B1(n_518), .B2(n_1172), .C(n_1331), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1353 ( .A1(n_43), .A2(n_109), .B1(n_1197), .B2(n_1354), .C(n_1355), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_43), .A2(n_109), .B1(n_1381), .B2(n_1383), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_44), .A2(n_167), .B1(n_455), .B2(n_612), .Y(n_660) );
INVx1_ASAP7_75t_L g707 ( .A(n_44), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g746 ( .A1(n_45), .A2(n_271), .B1(n_479), .B2(n_747), .C(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g1086 ( .A(n_46), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g1359 ( .A1(n_47), .A2(n_223), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_47), .A2(n_305), .B1(n_544), .B2(n_995), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_48), .Y(n_334) );
XNOR2xp5_ASAP7_75t_L g1714 ( .A(n_49), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1664 ( .A(n_50), .Y(n_1664) );
OAI22xp5_ASAP7_75t_L g1687 ( .A1(n_50), .A2(n_273), .B1(n_1344), .B2(n_1688), .Y(n_1687) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_51), .A2(n_293), .B1(n_1041), .B2(n_1042), .C(n_1043), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_51), .A2(n_156), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI21xp5_ASAP7_75t_L g1092 ( .A1(n_52), .A2(n_544), .B(n_1043), .Y(n_1092) );
INVxp67_ASAP7_75t_SL g1118 ( .A(n_52), .Y(n_1118) );
INVx1_ASAP7_75t_L g1147 ( .A(n_53), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_53), .A2(n_164), .B1(n_485), .B2(n_1172), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_54), .A2(n_173), .B1(n_379), .B2(n_386), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_54), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_55), .A2(n_102), .B1(n_1439), .B2(n_1456), .Y(n_1455) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_56), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_57), .A2(n_222), .B1(n_1439), .B2(n_1456), .Y(n_1476) );
INVx1_ASAP7_75t_L g801 ( .A(n_58), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_58), .A2(n_61), .B1(n_602), .B2(n_612), .Y(n_825) );
INVx1_ASAP7_75t_L g1046 ( .A(n_59), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_60), .A2(n_188), .B1(n_601), .B2(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g701 ( .A(n_60), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_61), .A2(n_297), .B1(n_563), .B2(n_788), .C(n_789), .Y(n_787) );
OAI222xp33_ASAP7_75t_L g933 ( .A1(n_62), .A2(n_77), .B1(n_934), .B2(n_938), .C1(n_945), .C2(n_953), .Y(n_933) );
INVx1_ASAP7_75t_L g981 ( .A(n_62), .Y(n_981) );
INVxp67_ASAP7_75t_SL g751 ( .A(n_63), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_63), .A2(n_386), .B1(n_773), .B2(n_775), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_64), .A2(n_219), .B1(n_362), .B2(n_367), .C(n_373), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_64), .A2(n_282), .B1(n_479), .B2(n_747), .C(n_749), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_65), .A2(n_252), .B1(n_379), .B2(n_386), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_65), .Y(n_1314) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_67), .A2(n_414), .B(n_417), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_67), .A2(n_98), .B1(n_515), .B2(n_517), .C(n_519), .Y(n_514) );
INVx1_ASAP7_75t_L g530 ( .A(n_68), .Y(n_530) );
INVx1_ASAP7_75t_L g1023 ( .A(n_69), .Y(n_1023) );
OAI21xp33_ASAP7_75t_L g1075 ( .A1(n_69), .A2(n_476), .B(n_479), .Y(n_1075) );
CKINVDCx5p33_ASAP7_75t_R g1287 ( .A(n_70), .Y(n_1287) );
INVx1_ASAP7_75t_L g1252 ( .A(n_71), .Y(n_1252) );
OAI211xp5_ASAP7_75t_L g1288 ( .A1(n_71), .A2(n_1228), .B(n_1232), .C(n_1289), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_72), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_73), .A2(n_206), .B1(n_1439), .B2(n_1456), .Y(n_1483) );
INVx1_ASAP7_75t_L g757 ( .A(n_74), .Y(n_757) );
OAI222xp33_ASAP7_75t_L g760 ( .A1(n_74), .A2(n_259), .B1(n_271), .B2(n_383), .C1(n_761), .C2(n_762), .Y(n_760) );
AOI21xp33_ASAP7_75t_L g1358 ( .A1(n_75), .A2(n_485), .B(n_1206), .Y(n_1358) );
INVx1_ASAP7_75t_L g1365 ( .A(n_75), .Y(n_1365) );
XOR2x2_ASAP7_75t_L g343 ( .A(n_76), .B(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g1464 ( .A1(n_76), .A2(n_215), .B1(n_1446), .B2(n_1449), .Y(n_1464) );
INVx1_ASAP7_75t_L g983 ( .A(n_77), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g1465 ( .A1(n_78), .A2(n_92), .B1(n_1439), .B2(n_1466), .Y(n_1465) );
AO22x1_ASAP7_75t_L g1445 ( .A1(n_79), .A2(n_224), .B1(n_1446), .B2(n_1449), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_80), .A2(n_115), .B1(n_632), .B2(n_634), .C(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g673 ( .A(n_80), .Y(n_673) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_81), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_83), .A2(n_177), .B1(n_972), .B2(n_989), .Y(n_1210) );
INVx1_ASAP7_75t_L g638 ( .A(n_84), .Y(n_638) );
OAI221xp5_ASAP7_75t_SL g684 ( .A1(n_84), .A2(n_112), .B1(n_365), .B2(n_569), .C(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_85), .A2(n_238), .B1(n_994), .B2(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1190 ( .A(n_86), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_87), .A2(n_286), .B1(n_770), .B2(n_1034), .C(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1431 ( .A(n_87), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_88), .A2(n_183), .B1(n_379), .B2(n_386), .Y(n_378) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_88), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g1727 ( .A1(n_89), .A2(n_107), .B1(n_562), .B2(n_1041), .C(n_1043), .Y(n_1727) );
AOI22xp33_ASAP7_75t_SL g1757 ( .A1(n_89), .A2(n_236), .B1(n_612), .B2(n_613), .Y(n_1757) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_90), .A2(n_136), .B1(n_294), .B2(n_388), .C1(n_419), .C2(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g522 ( .A(n_90), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_91), .Y(n_738) );
INVx1_ASAP7_75t_L g1303 ( .A(n_93), .Y(n_1303) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_93), .A2(n_172), .B1(n_1323), .B2(n_1325), .C(n_1327), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g808 ( .A1(n_94), .A2(n_133), .B1(n_362), .B2(n_367), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_94), .A2(n_257), .B1(n_747), .B2(n_749), .Y(n_826) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_95), .Y(n_946) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_95), .A2(n_247), .B1(n_544), .B2(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1678 ( .A(n_96), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1694 ( .A1(n_96), .A2(n_221), .B1(n_602), .B2(n_612), .Y(n_1694) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_97), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_98), .A2(n_192), .B1(n_391), .B2(n_394), .C(n_398), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_99), .A2(n_241), .B1(n_557), .B2(n_564), .Y(n_1224) );
INVx1_ASAP7_75t_L g320 ( .A(n_100), .Y(n_320) );
INVx1_ASAP7_75t_L g796 ( .A(n_101), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_101), .A2(n_297), .B1(n_455), .B2(n_612), .Y(n_820) );
INVx1_ASAP7_75t_L g752 ( .A(n_103), .Y(n_752) );
AO221x2_ASAP7_75t_L g1537 ( .A1(n_104), .A2(n_295), .B1(n_1446), .B2(n_1449), .C(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g360 ( .A(n_105), .Y(n_360) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_105), .A2(n_450), .B(n_459), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_106), .A2(n_138), .B1(n_653), .B2(n_657), .C(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g692 ( .A(n_106), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g1747 ( .A1(n_107), .A2(n_142), .B1(n_657), .B2(n_1693), .C(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g839 ( .A(n_108), .Y(n_839) );
INVx1_ASAP7_75t_L g1156 ( .A(n_110), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_110), .A2(n_147), .B1(n_455), .B2(n_612), .Y(n_1170) );
XOR2x2_ASAP7_75t_L g1392 ( .A(n_111), .B(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g648 ( .A(n_112), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_113), .Y(n_1144) );
INVx1_ASAP7_75t_L g970 ( .A(n_114), .Y(n_970) );
INVx1_ASAP7_75t_L g667 ( .A(n_115), .Y(n_667) );
INVx1_ASAP7_75t_L g1406 ( .A(n_116), .Y(n_1406) );
INVx1_ASAP7_75t_L g1411 ( .A(n_117), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_118), .A2(n_203), .B1(n_613), .B2(n_1174), .Y(n_1352) );
INVx1_ASAP7_75t_L g1368 ( .A(n_118), .Y(n_1368) );
OAI221xp5_ASAP7_75t_L g1137 ( .A1(n_119), .A2(n_250), .B1(n_379), .B2(n_386), .C(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1175 ( .A(n_119), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_120), .A2(n_527), .B1(n_528), .B2(n_622), .Y(n_526) );
INVx1_ASAP7_75t_L g622 ( .A(n_120), .Y(n_622) );
INVx1_ASAP7_75t_L g1410 ( .A(n_121), .Y(n_1410) );
INVx1_ASAP7_75t_L g642 ( .A(n_122), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_122), .A2(n_681), .B(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g1673 ( .A1(n_123), .A2(n_245), .B1(n_1042), .B2(n_1674), .Y(n_1673) );
AOI21xp33_ASAP7_75t_L g1692 ( .A1(n_123), .A2(n_662), .B(n_1693), .Y(n_1692) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_124), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_125), .A2(n_175), .B1(n_407), .B2(n_410), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_125), .A2(n_248), .B1(n_462), .B2(n_471), .Y(n_1420) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_126), .A2(n_281), .B1(n_894), .B2(n_895), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_126), .A2(n_281), .B1(n_902), .B2(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g1249 ( .A(n_127), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_128), .A2(n_189), .B1(n_379), .B2(n_386), .Y(n_1398) );
INVxp67_ASAP7_75t_SL g1418 ( .A(n_128), .Y(n_1418) );
AO22x1_ASAP7_75t_L g1461 ( .A1(n_129), .A2(n_298), .B1(n_1446), .B2(n_1449), .Y(n_1461) );
INVx1_ASAP7_75t_L g724 ( .A(n_130), .Y(n_724) );
INVx1_ASAP7_75t_L g942 ( .A(n_131), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_131), .A2(n_179), .B1(n_997), .B2(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1736 ( .A(n_132), .Y(n_1736) );
INVx1_ASAP7_75t_L g815 ( .A(n_133), .Y(n_815) );
AOI221xp5_ASAP7_75t_SL g652 ( .A1(n_134), .A2(n_277), .B1(n_653), .B2(n_657), .C(n_658), .Y(n_652) );
INVx1_ASAP7_75t_L g704 ( .A(n_134), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_135), .Y(n_650) );
INVx1_ASAP7_75t_L g489 ( .A(n_136), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_137), .A2(n_184), .B1(n_496), .B2(n_944), .C(n_1245), .Y(n_1244) );
INVxp67_ASAP7_75t_L g1268 ( .A(n_137), .Y(n_1268) );
INVx1_ASAP7_75t_L g708 ( .A(n_138), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_139), .A2(n_305), .B1(n_662), .B2(n_1169), .C(n_1351), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_139), .A2(n_223), .B1(n_544), .B2(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1030 ( .A(n_140), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_140), .A2(n_151), .B1(n_1054), .B2(n_1055), .Y(n_1053) );
INVx1_ASAP7_75t_L g1140 ( .A(n_141), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_141), .A2(n_289), .B1(n_462), .B2(n_471), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1722 ( .A1(n_142), .A2(n_165), .B1(n_547), .B2(n_559), .C(n_1723), .Y(n_1722) );
AOI221xp5_ASAP7_75t_L g1304 ( .A1(n_143), .A2(n_172), .B1(n_770), .B2(n_1305), .C(n_1306), .Y(n_1304) );
INVx1_ASAP7_75t_L g1335 ( .A(n_143), .Y(n_1335) );
AO22x1_ASAP7_75t_L g1438 ( .A1(n_144), .A2(n_299), .B1(n_1439), .B2(n_1443), .Y(n_1438) );
CKINVDCx16_ASAP7_75t_R g1539 ( .A(n_145), .Y(n_1539) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_146), .Y(n_536) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_146), .A2(n_373), .B1(n_379), .B2(n_566), .C(n_575), .Y(n_565) );
INVx1_ASAP7_75t_L g1151 ( .A(n_147), .Y(n_1151) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_148), .A2(n_557), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g596 ( .A(n_148), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1697 ( .A1(n_149), .A2(n_245), .B1(n_602), .B2(n_612), .Y(n_1697) );
INVx1_ASAP7_75t_L g574 ( .A(n_150), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_150), .A2(n_193), .B1(n_599), .B2(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g1039 ( .A(n_151), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_152), .A2(n_307), .B1(n_388), .B2(n_563), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1127 ( .A(n_152), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1397 ( .A1(n_153), .A2(n_248), .B1(n_362), .B2(n_367), .C(n_373), .Y(n_1397) );
INVxp67_ASAP7_75t_SL g1416 ( .A(n_153), .Y(n_1416) );
INVx1_ASAP7_75t_L g803 ( .A(n_154), .Y(n_803) );
INVx1_ASAP7_75t_L g1090 ( .A(n_155), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g1031 ( .A1(n_156), .A2(n_269), .B1(n_559), .B2(n_1032), .C(n_1034), .Y(n_1031) );
INVx1_ASAP7_75t_L g882 ( .A(n_157), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g906 ( .A1(n_157), .A2(n_854), .B(n_907), .C(n_909), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g1732 ( .A1(n_158), .A2(n_159), .B1(n_798), .B2(n_1369), .C(n_1733), .Y(n_1732) );
INVxp67_ASAP7_75t_SL g1744 ( .A(n_159), .Y(n_1744) );
INVxp33_ASAP7_75t_SL g1750 ( .A(n_160), .Y(n_1750) );
INVx2_ASAP7_75t_L g1442 ( .A(n_161), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_161), .B(n_266), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_161), .B(n_1448), .Y(n_1450) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_162), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_162), .A2(n_279), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g1340 ( .A(n_163), .B(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1155 ( .A(n_164), .Y(n_1155) );
INVx1_ASAP7_75t_L g1754 ( .A(n_165), .Y(n_1754) );
INVx1_ASAP7_75t_L g1176 ( .A(n_166), .Y(n_1176) );
INVx1_ASAP7_75t_L g691 ( .A(n_167), .Y(n_691) );
INVx1_ASAP7_75t_L g1098 ( .A(n_168), .Y(n_1098) );
OAI221xp5_ASAP7_75t_L g1312 ( .A1(n_169), .A2(n_242), .B1(n_362), .B2(n_367), .C(n_373), .Y(n_1312) );
INVx1_ASAP7_75t_L g1339 ( .A(n_169), .Y(n_1339) );
OAI21xp5_ASAP7_75t_SL g1015 ( .A1(n_170), .A2(n_1016), .B(n_1017), .Y(n_1015) );
INVx1_ASAP7_75t_L g1045 ( .A(n_170), .Y(n_1045) );
INVx1_ASAP7_75t_L g837 ( .A(n_171), .Y(n_837) );
INVx1_ASAP7_75t_L g1069 ( .A(n_173), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g1201 ( .A(n_174), .Y(n_1201) );
OAI211xp5_ASAP7_75t_L g1413 ( .A1(n_175), .A2(n_1016), .B(n_1414), .C(n_1417), .Y(n_1413) );
INVx1_ASAP7_75t_L g1735 ( .A(n_176), .Y(n_1735) );
OAI22xp5_ASAP7_75t_L g1758 ( .A1(n_176), .A2(n_202), .B1(n_462), .B2(n_471), .Y(n_1758) );
OAI211xp5_ASAP7_75t_L g1180 ( .A1(n_177), .A2(n_957), .B(n_1181), .C(n_1189), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_178), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_179), .A2(n_311), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx2_ASAP7_75t_L g359 ( .A(n_180), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_180), .B(n_357), .Y(n_382) );
INVx1_ASAP7_75t_L g424 ( .A(n_180), .Y(n_424) );
INVx1_ASAP7_75t_L g1386 ( .A(n_181), .Y(n_1386) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_182), .A2(n_373), .B(n_1020), .C(n_1021), .Y(n_1019) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_182), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_183), .Y(n_429) );
INVxp67_ASAP7_75t_L g1278 ( .A(n_184), .Y(n_1278) );
INVx1_ASAP7_75t_L g717 ( .A(n_185), .Y(n_717) );
OAI221xp5_ASAP7_75t_SL g1195 ( .A1(n_186), .A2(n_267), .B1(n_934), .B2(n_1196), .C(n_1198), .Y(n_1195) );
INVx1_ASAP7_75t_L g1214 ( .A(n_186), .Y(n_1214) );
INVx1_ASAP7_75t_L g1159 ( .A(n_187), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_187), .A2(n_284), .B1(n_636), .B2(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g705 ( .A(n_188), .Y(n_705) );
INVxp67_ASAP7_75t_SL g1415 ( .A(n_189), .Y(n_1415) );
INVx1_ASAP7_75t_L g941 ( .A(n_190), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_190), .A2(n_311), .B1(n_998), .B2(n_1000), .Y(n_999) );
BUFx3_ASAP7_75t_L g351 ( .A(n_191), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_192), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g400 ( .A(n_194), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_195), .A2(n_199), .B1(n_1446), .B2(n_1449), .Y(n_1484) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_196), .A2(n_257), .B1(n_554), .B2(n_805), .C(n_806), .Y(n_804) );
OAI211xp5_ASAP7_75t_L g811 ( .A1(n_196), .A2(n_812), .B(n_813), .C(n_816), .Y(n_811) );
OAI21xp5_ASAP7_75t_SL g971 ( .A1(n_197), .A2(n_972), .B(n_973), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_198), .Y(n_790) );
XOR2xp5_ASAP7_75t_L g1177 ( .A(n_199), .B(n_1178), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_201), .A2(n_241), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
INVx1_ASAP7_75t_L g1729 ( .A(n_202), .Y(n_1729) );
INVx1_ASAP7_75t_L g1375 ( .A(n_203), .Y(n_1375) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_204), .Y(n_1209) );
INVx1_ASAP7_75t_L g1106 ( .A(n_205), .Y(n_1106) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_207), .Y(n_535) );
INVx1_ASAP7_75t_L g1404 ( .A(n_208), .Y(n_1404) );
INVx1_ASAP7_75t_L g1661 ( .A(n_209), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_210), .Y(n_732) );
INVx1_ASAP7_75t_L g967 ( .A(n_211), .Y(n_967) );
OAI211xp5_ASAP7_75t_L g1141 ( .A1(n_212), .A2(n_348), .B(n_373), .C(n_1142), .Y(n_1141) );
INVxp33_ASAP7_75t_SL g1165 ( .A(n_212), .Y(n_1165) );
INVx1_ASAP7_75t_L g1396 ( .A(n_213), .Y(n_1396) );
INVx1_ASAP7_75t_L g1348 ( .A(n_214), .Y(n_1348) );
BUFx3_ASAP7_75t_L g337 ( .A(n_216), .Y(n_337) );
INVx1_ASAP7_75t_L g437 ( .A(n_216), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g1541 ( .A(n_217), .Y(n_1541) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_218), .A2(n_233), .B1(n_1446), .B2(n_1449), .Y(n_1475) );
INVxp67_ASAP7_75t_SL g1131 ( .A(n_219), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g956 ( .A1(n_220), .A2(n_957), .B(n_959), .C(n_965), .Y(n_956) );
INVx1_ASAP7_75t_L g987 ( .A(n_220), .Y(n_987) );
INVx1_ASAP7_75t_L g1672 ( .A(n_221), .Y(n_1672) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_225), .B(n_617), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_226), .Y(n_637) );
INVx1_ASAP7_75t_L g549 ( .A(n_227), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_228), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g1298 ( .A1(n_229), .A2(n_291), .B1(n_770), .B2(n_1299), .C(n_1300), .Y(n_1298) );
INVx1_ASAP7_75t_L g1328 ( .A(n_229), .Y(n_1328) );
INVx1_ASAP7_75t_L g1301 ( .A(n_230), .Y(n_1301) );
INVx1_ASAP7_75t_L g853 ( .A(n_232), .Y(n_853) );
XOR2xp5_ASAP7_75t_L g1293 ( .A(n_233), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g403 ( .A(n_234), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_235), .Y(n_570) );
XOR2x2_ASAP7_75t_L g930 ( .A(n_237), .B(n_931), .Y(n_930) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_238), .Y(n_1199) );
AOI211xp5_ASAP7_75t_L g1400 ( .A1(n_240), .A2(n_1041), .B(n_1401), .C(n_1403), .Y(n_1400) );
INVx1_ASAP7_75t_L g1428 ( .A(n_240), .Y(n_1428) );
INVxp67_ASAP7_75t_SL g1318 ( .A(n_242), .Y(n_1318) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_243), .A2(n_301), .B1(n_1446), .B2(n_1449), .Y(n_1454) );
AO22x1_ASAP7_75t_L g1460 ( .A1(n_244), .A2(n_251), .B1(n_1439), .B2(n_1456), .Y(n_1460) );
INVx1_ASAP7_75t_L g354 ( .A(n_246), .Y(n_354) );
INVx1_ASAP7_75t_L g372 ( .A(n_246), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_247), .A2(n_279), .B1(n_496), .B2(n_653), .C(n_662), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_249), .Y(n_728) );
INVxp67_ASAP7_75t_SL g1163 ( .A(n_250), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1650 ( .A1(n_251), .A2(n_1651), .B1(n_1652), .B2(n_1701), .Y(n_1650) );
INVxp67_ASAP7_75t_L g1701 ( .A(n_251), .Y(n_1701) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_251), .A2(n_1708), .B1(n_1713), .B2(n_1759), .Y(n_1707) );
INVx1_ASAP7_75t_L g1321 ( .A(n_252), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_253), .A2(n_285), .B1(n_407), .B2(n_410), .Y(n_1297) );
INVx1_ASAP7_75t_L g1319 ( .A(n_253), .Y(n_1319) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_254), .Y(n_443) );
INVx1_ASAP7_75t_L g844 ( .A(n_255), .Y(n_844) );
AOI21xp33_ASAP7_75t_L g1102 ( .A1(n_256), .A2(n_559), .B(n_697), .Y(n_1102) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_256), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1656 ( .A(n_258), .Y(n_1656) );
OAI221xp5_ASAP7_75t_L g1699 ( .A1(n_258), .A2(n_292), .B1(n_508), .B2(n_1197), .C(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g780 ( .A(n_259), .Y(n_780) );
INVx1_ASAP7_75t_L g1734 ( .A(n_260), .Y(n_1734) );
NOR2xp33_ASAP7_75t_L g1737 ( .A(n_260), .B(n_1016), .Y(n_1737) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_261), .Y(n_1662) );
INVxp33_ASAP7_75t_L g1274 ( .A(n_262), .Y(n_1274) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_263), .Y(n_1356) );
INVx1_ASAP7_75t_L g1280 ( .A(n_264), .Y(n_1280) );
INVx1_ASAP7_75t_L g582 ( .A(n_265), .Y(n_582) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_266), .B(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1448 ( .A(n_266), .Y(n_1448) );
INVx1_ASAP7_75t_L g1215 ( .A(n_267), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_268), .Y(n_978) );
AOI221xp5_ASAP7_75t_SL g1058 ( .A1(n_269), .A2(n_270), .B1(n_1051), .B2(n_1059), .C(n_1060), .Y(n_1058) );
INVx1_ASAP7_75t_L g1038 ( .A(n_270), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_272), .A2(n_1013), .B1(n_1014), .B2(n_1078), .Y(n_1012) );
INVx1_ASAP7_75t_L g1078 ( .A(n_272), .Y(n_1078) );
INVx1_ASAP7_75t_L g1666 ( .A(n_273), .Y(n_1666) );
INVx1_ASAP7_75t_L g841 ( .A(n_274), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g1677 ( .A(n_275), .Y(n_1677) );
XOR2x2_ASAP7_75t_L g1082 ( .A(n_276), .B(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g695 ( .A(n_277), .Y(n_695) );
INVx1_ASAP7_75t_L g1402 ( .A(n_278), .Y(n_1402) );
INVx1_ASAP7_75t_L g550 ( .A(n_280), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_280), .A2(n_476), .B1(n_604), .B2(n_614), .C(n_615), .Y(n_603) );
INVx1_ASAP7_75t_L g1255 ( .A(n_283), .Y(n_1255) );
INVx1_ASAP7_75t_L g1153 ( .A(n_284), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1337 ( .A(n_285), .Y(n_1337) );
INVx1_ASAP7_75t_L g1424 ( .A(n_286), .Y(n_1424) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
INVx1_ASAP7_75t_L g1095 ( .A(n_288), .Y(n_1095) );
INVx1_ASAP7_75t_L g1143 ( .A(n_289), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_290), .Y(n_795) );
INVx1_ASAP7_75t_L g1332 ( .A(n_291), .Y(n_1332) );
INVx1_ASAP7_75t_L g1659 ( .A(n_292), .Y(n_1659) );
INVx1_ASAP7_75t_L g1063 ( .A(n_293), .Y(n_1063) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_294), .A2(n_496), .B(n_499), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_296), .Y(n_725) );
INVx2_ASAP7_75t_L g427 ( .A(n_300), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_300), .Y(n_434) );
INVx1_ASAP7_75t_L g454 ( .A(n_300), .Y(n_454) );
XOR2x2_ASAP7_75t_L g830 ( .A(n_301), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g1308 ( .A(n_302), .Y(n_1308) );
INVx1_ASAP7_75t_L g460 ( .A(n_303), .Y(n_460) );
INVx1_ASAP7_75t_L g783 ( .A(n_304), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_306), .Y(n_552) );
INVxp67_ASAP7_75t_SL g1116 ( .A(n_307), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_308), .Y(n_1241) );
OAI21xp33_ASAP7_75t_SL g1135 ( .A1(n_309), .A2(n_1016), .B(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1139 ( .A(n_309), .Y(n_1139) );
INVx1_ASAP7_75t_L g855 ( .A(n_310), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_338), .B(n_1433), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_317), .B(n_326), .Y(n_1706) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g1712 ( .A(n_319), .B(n_322), .Y(n_1712) );
INVx1_ASAP7_75t_L g1762 ( .A(n_319), .Y(n_1762) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_322), .B(n_1762), .Y(n_1764) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g898 ( .A(n_326), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g510 ( .A(n_327), .B(n_337), .Y(n_510) );
AND2x4_ASAP7_75t_L g659 ( .A(n_327), .B(n_336), .Y(n_659) );
INVx1_ASAP7_75t_L g894 ( .A(n_328), .Y(n_894) );
AND2x4_ASAP7_75t_SL g1705 ( .A(n_328), .B(n_1706), .Y(n_1705) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_330), .B(n_335), .Y(n_329) );
BUFx4f_ASAP7_75t_L g488 ( .A(n_330), .Y(n_488) );
INVxp67_ASAP7_75t_L g741 ( .A(n_330), .Y(n_741) );
OR2x6_ASAP7_75t_L g888 ( .A(n_330), .B(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1334 ( .A(n_330), .Y(n_1334) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g521 ( .A(n_331), .Y(n_521) );
BUFx4f_ASAP7_75t_L g633 ( .A(n_331), .Y(n_633) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g439 ( .A(n_333), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g447 ( .A(n_333), .Y(n_447) );
INVx2_ASAP7_75t_L g458 ( .A(n_333), .Y(n_458) );
INVx1_ASAP7_75t_L g474 ( .A(n_333), .Y(n_474) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_333), .B(n_334), .Y(n_478) );
AND2x2_ASAP7_75t_L g498 ( .A(n_333), .B(n_334), .Y(n_498) );
INVx2_ASAP7_75t_L g440 ( .A(n_334), .Y(n_440) );
INVx1_ASAP7_75t_L g448 ( .A(n_334), .Y(n_448) );
AND2x2_ASAP7_75t_L g457 ( .A(n_334), .B(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g468 ( .A(n_334), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_334), .B(n_458), .Y(n_494) );
OR2x2_ASAP7_75t_L g595 ( .A(n_334), .B(n_447), .Y(n_595) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g877 ( .A(n_336), .Y(n_877) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g881 ( .A(n_337), .Y(n_881) );
AND2x4_ASAP7_75t_L g885 ( .A(n_337), .B(n_473), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_1008), .B2(n_1009), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_712), .B1(n_713), .B2(n_1007), .Y(n_340) );
INVx1_ASAP7_75t_L g1007 ( .A(n_341), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_524), .B1(n_710), .B2(n_711), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g710 ( .A(n_343), .Y(n_710) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_345), .B(n_441), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_389), .B(n_425), .C(n_428), .Y(n_345) );
AOI211xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_360), .B(n_361), .C(n_378), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_347), .A2(n_752), .B1(n_760), .B2(n_763), .C(n_764), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_347), .A2(n_763), .B1(n_803), .B2(n_804), .C(n_808), .Y(n_802) );
INVx2_ASAP7_75t_L g1020 ( .A(n_347), .Y(n_1020) );
AOI211xp5_ASAP7_75t_L g1085 ( .A1(n_347), .A2(n_1086), .B(n_1087), .C(n_1088), .Y(n_1085) );
AOI211xp5_ASAP7_75t_SL g1309 ( .A1(n_347), .A2(n_1310), .B(n_1311), .C(n_1312), .Y(n_1309) );
AOI211xp5_ASAP7_75t_L g1395 ( .A1(n_347), .A2(n_1396), .B(n_1397), .C(n_1398), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1731 ( .A1(n_347), .A2(n_540), .B1(n_1732), .B2(n_1736), .Y(n_1731) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g532 ( .A(n_348), .B(n_533), .Y(n_532) );
OR2x6_ASAP7_75t_L g989 ( .A(n_348), .B(n_533), .Y(n_989) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .Y(n_348) );
BUFx3_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
AND2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_409), .Y(n_408) );
INVx8_ASAP7_75t_L g545 ( .A(n_349), .Y(n_545) );
BUFx3_ASAP7_75t_L g563 ( .A(n_349), .Y(n_563) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
AND2x4_ASAP7_75t_L g384 ( .A(n_350), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_351), .Y(n_366) );
AND2x4_ASAP7_75t_L g412 ( .A(n_351), .B(n_371), .Y(n_412) );
OR2x2_ASAP7_75t_L g420 ( .A(n_351), .B(n_353), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_351), .B(n_372), .Y(n_581) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
AND2x6_ASAP7_75t_L g363 ( .A(n_355), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g368 ( .A(n_355), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
AND2x4_ASAP7_75t_L g686 ( .A(n_355), .B(n_506), .Y(n_686) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_356), .B(n_424), .Y(n_423) );
NAND3x1_ASAP7_75t_L g850 ( .A(n_356), .B(n_424), .C(n_851), .Y(n_850) );
OR2x4_ASAP7_75t_L g902 ( .A(n_356), .B(n_420), .Y(n_902) );
INVx1_ASAP7_75t_L g905 ( .A(n_356), .Y(n_905) );
AND2x4_ASAP7_75t_L g908 ( .A(n_356), .B(n_412), .Y(n_908) );
OR2x6_ASAP7_75t_L g923 ( .A(n_356), .B(n_700), .Y(n_923) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
NAND2xp33_ASAP7_75t_SL g560 ( .A(n_357), .B(n_359), .Y(n_560) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g404 ( .A(n_359), .B(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_359), .Y(n_927) );
AND3x4_ASAP7_75t_L g992 ( .A(n_359), .B(n_405), .C(n_426), .Y(n_992) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_363), .A2(n_368), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_363), .A2(n_368), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_363), .A2(n_368), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
AOI221xp5_ASAP7_75t_L g1728 ( .A1(n_363), .A2(n_368), .B1(n_766), .B2(n_1729), .C(n_1730), .Y(n_1728) );
AND2x2_ASAP7_75t_L g982 ( .A(n_364), .B(n_686), .Y(n_982) );
NAND2x1_ASAP7_75t_L g1291 ( .A(n_364), .B(n_686), .Y(n_1291) );
AND2x4_ASAP7_75t_SL g1382 ( .A(n_364), .B(n_686), .Y(n_1382) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_366), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g388 ( .A(n_366), .B(n_370), .Y(n_388) );
BUFx2_ASAP7_75t_L g913 ( .A(n_366), .Y(n_913) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g685 ( .A(n_369), .Y(n_685) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_372), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_373), .Y(n_766) );
OR2x6_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g416 ( .A(n_374), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g794 ( .A1(n_374), .A2(n_422), .B1(n_573), .B2(n_795), .C(n_796), .Y(n_794) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_375), .Y(n_397) );
BUFx3_ASAP7_75t_L g569 ( .A(n_375), .Y(n_569) );
BUFx2_ASAP7_75t_L g916 ( .A(n_376), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_379), .Y(n_1105) );
OR2x6_ASAP7_75t_SL g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g387 ( .A(n_381), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_381), .Y(n_542) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
OR2x2_ASAP7_75t_L g671 ( .A(n_382), .B(n_513), .Y(n_671) );
INVx3_ASAP7_75t_L g675 ( .A(n_383), .Y(n_675) );
BUFx2_ASAP7_75t_L g843 ( .A(n_383), .Y(n_843) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_383), .Y(n_1222) );
INVx1_ASAP7_75t_L g1270 ( .A(n_383), .Y(n_1270) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_384), .Y(n_393) );
BUFx8_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_384), .Y(n_697) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_387), .B(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g1104 ( .A1(n_387), .A2(n_1105), .B1(n_1106), .B2(n_1107), .C(n_1108), .Y(n_1104) );
INVx5_ASAP7_75t_L g399 ( .A(n_388), .Y(n_399) );
BUFx3_ASAP7_75t_L g770 ( .A(n_388), .Y(n_770) );
BUFx12f_ASAP7_75t_L g788 ( .A(n_388), .Y(n_788) );
BUFx3_ASAP7_75t_L g998 ( .A(n_388), .Y(n_998) );
BUFx2_ASAP7_75t_L g1721 ( .A(n_388), .Y(n_1721) );
NOR3xp33_ASAP7_75t_SL g389 ( .A(n_390), .B(n_406), .C(n_413), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g792 ( .A(n_393), .Y(n_792) );
INVx2_ASAP7_75t_L g840 ( .A(n_393), .Y(n_840) );
AND2x4_ASAP7_75t_L g904 ( .A(n_393), .B(n_905), .Y(n_904) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_393), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g1374 ( .A(n_393), .Y(n_1374) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g1091 ( .A(n_396), .Y(n_1091) );
INVx4_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g555 ( .A(n_397), .Y(n_555) );
OR2x2_ASAP7_75t_L g678 ( .A(n_397), .B(n_671), .Y(n_678) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_397), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_397), .A2(n_404), .B1(n_790), .B2(n_791), .C(n_792), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_401), .B2(n_403), .C(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g564 ( .A(n_399), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_400), .A2(n_520), .B1(n_522), .B2(n_523), .Y(n_519) );
INVx2_ASAP7_75t_L g1219 ( .A(n_401), .Y(n_1219) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_402), .B(n_807), .Y(n_806) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_402), .Y(n_1042) );
INVx1_ASAP7_75t_L g1681 ( .A(n_402), .Y(n_1681) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_403), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g771 ( .A1(n_404), .A2(n_569), .B1(n_703), .B2(n_732), .C(n_736), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_404), .A2(n_693), .B1(n_1147), .B2(n_1148), .C(n_1149), .Y(n_1146) );
OAI221xp5_ASAP7_75t_L g1300 ( .A1(n_404), .A2(n_569), .B1(n_1301), .B2(n_1302), .C(n_1303), .Y(n_1300) );
OAI21xp33_ASAP7_75t_L g1401 ( .A1(n_404), .A2(n_1148), .B(n_1402), .Y(n_1401) );
INVx3_ASAP7_75t_L g912 ( .A(n_405), .Y(n_912) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_408), .A2(n_411), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_408), .A2(n_411), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AND2x2_ASAP7_75t_L g411 ( .A(n_409), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g547 ( .A(n_412), .Y(n_547) );
BUFx2_ASAP7_75t_L g995 ( .A(n_412), .Y(n_995) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_412), .Y(n_1003) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_412), .Y(n_1033) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_412), .Y(n_1041) );
INVx2_ASAP7_75t_L g1378 ( .A(n_412), .Y(n_1378) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .Y(n_417) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_419), .Y(n_1028) );
INVx3_ASAP7_75t_L g1152 ( .A(n_419), .Y(n_1152) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_420), .Y(n_573) );
BUFx3_ASAP7_75t_L g761 ( .A(n_420), .Y(n_761) );
BUFx3_ASAP7_75t_L g774 ( .A(n_420), .Y(n_774) );
OR2x4_ASAP7_75t_L g921 ( .A(n_420), .B(n_905), .Y(n_921) );
INVx3_ASAP7_75t_L g558 ( .A(n_421), .Y(n_558) );
INVx2_ASAP7_75t_SL g576 ( .A(n_421), .Y(n_576) );
AND2x4_ASAP7_75t_L g974 ( .A(n_421), .B(n_670), .Y(n_974) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_421), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_421), .Y(n_1094) );
INVx3_ASAP7_75t_L g1148 ( .A(n_421), .Y(n_1148) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_422), .A2(n_567), .B1(n_570), .B2(n_571), .C(n_574), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_422), .A2(n_569), .B1(n_725), .B2(n_738), .C(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g1043 ( .A(n_422), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_422), .A2(n_774), .B1(n_1091), .B2(n_1155), .C(n_1156), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_422), .A2(n_569), .B1(n_573), .B2(n_1307), .C(n_1308), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1409 ( .A1(n_422), .A2(n_569), .B1(n_774), .B2(n_1410), .C(n_1411), .Y(n_1409) );
INVx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g709 ( .A(n_423), .B(n_501), .Y(n_709) );
O2A1O1Ixp5_ASAP7_75t_L g932 ( .A1(n_425), .A2(n_933), .B(n_956), .C(n_971), .Y(n_932) );
INVx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g585 ( .A(n_426), .Y(n_585) );
OAI31xp33_ASAP7_75t_SL g1136 ( .A1(n_426), .A2(n_1137), .A3(n_1141), .B(n_1145), .Y(n_1136) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_427), .B(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g529 ( .A1(n_430), .A2(n_444), .B1(n_530), .B2(n_531), .C1(n_535), .C2(n_536), .Y(n_529) );
NAND2xp33_ASAP7_75t_SL g779 ( .A(n_430), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g812 ( .A(n_430), .Y(n_812) );
INVx1_ASAP7_75t_L g1071 ( .A(n_430), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_430), .B(n_1106), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_430), .B(n_1163), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_430), .B(n_1418), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1745 ( .A(n_430), .Y(n_1745) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_435), .Y(n_430) );
AND2x4_ASAP7_75t_L g444 ( .A(n_431), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g533 ( .A(n_432), .Y(n_533) );
OR2x2_ASAP7_75t_L g749 ( .A(n_432), .B(n_472), .Y(n_749) );
INVx1_ASAP7_75t_L g899 ( .A(n_432), .Y(n_899) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g513 ( .A(n_433), .Y(n_513) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
AND2x2_ASAP7_75t_L g445 ( .A(n_436), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_436), .B(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g639 ( .A(n_436), .Y(n_639) );
AND2x4_ASAP7_75t_SL g937 ( .A(n_436), .B(n_497), .Y(n_937) );
AND2x4_ASAP7_75t_L g958 ( .A(n_436), .B(n_602), .Y(n_958) );
AND2x4_ASAP7_75t_L g969 ( .A(n_436), .B(n_438), .Y(n_969) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_436), .B(n_455), .Y(n_1345) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_437), .Y(n_889) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
INVx2_ASAP7_75t_L g1247 ( .A(n_438), .Y(n_1247) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g518 ( .A(n_439), .Y(n_518) );
INVx2_ASAP7_75t_L g656 ( .A(n_439), .Y(n_656) );
AND2x4_ASAP7_75t_L g896 ( .A(n_439), .B(n_889), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_482), .Y(n_441) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_449), .C(n_475), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_444), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_444), .B(n_807), .Y(n_810) );
INVx3_ASAP7_75t_L g1016 ( .A(n_444), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_444), .B(n_1337), .Y(n_1336) );
BUFx6f_ASAP7_75t_L g966 ( .A(n_445), .Y(n_966) );
INVx1_ASAP7_75t_L g1251 ( .A(n_445), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_446), .B(n_465), .Y(n_508) );
INVx3_ASAP7_75t_L g600 ( .A(n_446), .Y(n_600) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_446), .Y(n_612) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g534 ( .A(n_451), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g750 ( .A1(n_451), .A2(n_504), .B1(n_751), .B2(n_752), .C1(n_753), .C2(n_755), .Y(n_750) );
AOI211xp5_ASAP7_75t_L g1073 ( .A1(n_451), .A2(n_1074), .B(n_1075), .C(n_1076), .Y(n_1073) );
AOI222xp33_ASAP7_75t_L g1130 ( .A1(n_451), .A2(n_504), .B1(n_753), .B2(n_1086), .C1(n_1107), .C2(n_1131), .Y(n_1130) );
AOI21xp33_ASAP7_75t_L g1164 ( .A1(n_451), .A2(n_1165), .B(n_1166), .Y(n_1164) );
AOI222xp33_ASAP7_75t_L g1317 ( .A1(n_451), .A2(n_461), .B1(n_470), .B2(n_1310), .C1(n_1318), .C2(n_1319), .Y(n_1317) );
AOI222xp33_ASAP7_75t_L g1414 ( .A1(n_451), .A2(n_504), .B1(n_753), .B2(n_1396), .C1(n_1415), .C2(n_1416), .Y(n_1414) );
INVxp67_ASAP7_75t_L g1742 ( .A(n_451), .Y(n_1742) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
AOI332xp33_ASAP7_75t_L g813 ( .A1(n_452), .A2(n_455), .A3(n_505), .B1(n_507), .B2(n_753), .B3(n_803), .C1(n_814), .C2(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g476 ( .A(n_453), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g754 ( .A(n_453), .B(n_477), .Y(n_754) );
INVx1_ASAP7_75t_L g506 ( .A(n_454), .Y(n_506) );
INVx1_ASAP7_75t_L g851 ( .A(n_454), .Y(n_851) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g1361 ( .A(n_456), .Y(n_1361) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_457), .Y(n_602) );
BUFx3_ASAP7_75t_L g613 ( .A(n_457), .Y(n_613) );
BUFx3_ASAP7_75t_L g636 ( .A(n_457), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_469), .B2(n_470), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_461), .A2(n_470), .B1(n_546), .B2(n_549), .Y(n_615) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g748 ( .A(n_462), .Y(n_748) );
HB1xp67_ASAP7_75t_L g1077 ( .A(n_462), .Y(n_1077) );
NAND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g481 ( .A(n_463), .Y(n_481) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_465), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g644 ( .A(n_465), .Y(n_644) );
AND2x2_ASAP7_75t_L g646 ( .A(n_465), .B(n_647), .Y(n_646) );
AND2x6_ASAP7_75t_L g964 ( .A(n_465), .B(n_497), .Y(n_964) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g647 ( .A(n_468), .Y(n_647) );
AND2x4_ASAP7_75t_L g880 ( .A(n_468), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g955 ( .A(n_468), .Y(n_955) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g972 ( .A(n_471), .B(n_678), .Y(n_972) );
AND2x4_ASAP7_75t_L g1388 ( .A(n_471), .B(n_678), .Y(n_1388) );
INVx1_ASAP7_75t_L g649 ( .A(n_472), .Y(n_649) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g737 ( .A(n_477), .Y(n_737) );
INVx2_ASAP7_75t_SL g940 ( .A(n_477), .Y(n_940) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_478), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_479), .A2(n_588), .B(n_592), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_479), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g1752 ( .A1(n_479), .A2(n_1066), .B(n_1753), .Y(n_1752) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_480), .Y(n_597) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_480), .Y(n_608) );
INVx4_ASAP7_75t_L g730 ( .A(n_480), .Y(n_730) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_480), .Y(n_824) );
BUFx4f_ASAP7_75t_L g1357 ( .A(n_480), .Y(n_1357) );
BUFx4f_ASAP7_75t_L g1423 ( .A(n_480), .Y(n_1423) );
AOI322xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .A3(n_495), .B1(n_503), .B2(n_504), .C1(n_509), .C2(n_514), .Y(n_482) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_488), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
INVx5_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx6_ASAP7_75t_L g1751 ( .A(n_491), .Y(n_1751) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g523 ( .A(n_492), .Y(n_523) );
INVx2_ASAP7_75t_SL g726 ( .A(n_492), .Y(n_726) );
INVx4_ASAP7_75t_L g862 ( .A(n_492), .Y(n_862) );
INVx2_ASAP7_75t_L g951 ( .A(n_492), .Y(n_951) );
INVx1_ASAP7_75t_L g1200 ( .A(n_492), .Y(n_1200) );
INVx8_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g892 ( .A(n_493), .B(n_881), .Y(n_892) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_493), .Y(n_1119) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_496), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_496), .A2(n_610), .B(n_642), .C(n_643), .Y(n_641) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_497), .Y(n_516) );
BUFx3_ASAP7_75t_L g657 ( .A(n_497), .Y(n_657) );
AND2x2_ASAP7_75t_L g876 ( .A(n_497), .B(n_877), .Y(n_876) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_497), .Y(n_1169) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_497), .Y(n_1172) );
INVx1_ASAP7_75t_L g1324 ( .A(n_497), .Y(n_1324) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g1205 ( .A(n_498), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_499), .A2(n_857), .A3(n_863), .B1(n_865), .B2(n_868), .B3(n_870), .Y(n_856) );
OAI33xp33_ASAP7_75t_L g1421 ( .A1(n_499), .A2(n_744), .A3(n_1422), .B1(n_1425), .B2(n_1427), .B3(n_1430), .Y(n_1421) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
INVx2_ASAP7_75t_L g722 ( .A(n_500), .Y(n_722) );
INVx2_ASAP7_75t_L g1067 ( .A(n_500), .Y(n_1067) );
AOI222xp33_ASAP7_75t_L g1320 ( .A1(n_500), .A2(n_504), .B1(n_509), .B2(n_1321), .C1(n_1322), .C2(n_1330), .Y(n_1320) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g621 ( .A(n_501), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g1048 ( .A1(n_504), .A2(n_509), .A3(n_1049), .B1(n_1053), .B2(n_1057), .C1(n_1058), .C2(n_1065), .Y(n_1048) );
AOI332xp33_ASAP7_75t_L g1167 ( .A1(n_504), .A2(n_509), .A3(n_590), .B1(n_1168), .B2(n_1170), .B3(n_1171), .C1(n_1173), .C2(n_1175), .Y(n_1167) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g619 ( .A(n_506), .B(n_508), .Y(n_619) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_509), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g1746 ( .A1(n_509), .A2(n_1747), .B(n_1752), .C(n_1758), .Y(n_1746) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx4_ASAP7_75t_L g662 ( .A(n_510), .Y(n_662) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_510), .B(n_513), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_510), .B(n_511), .Y(n_821) );
INVx4_ASAP7_75t_L g1184 ( .A(n_510), .Y(n_1184) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g689 ( .A(n_513), .B(n_560), .Y(n_689) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_513), .Y(n_929) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g1052 ( .A(n_516), .Y(n_1052) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g1326 ( .A(n_518), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_520), .A2(n_726), .B1(n_1406), .B2(n_1431), .Y(n_1430) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g860 ( .A(n_521), .Y(n_860) );
INVx2_ASAP7_75t_SL g948 ( .A(n_521), .Y(n_948) );
BUFx6f_ASAP7_75t_L g1117 ( .A(n_521), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_523), .A2(n_1404), .B1(n_1411), .B2(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g711 ( .A(n_524), .Y(n_711) );
XOR2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_623), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .C(n_586), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_535), .A2(n_544), .B1(n_546), .B2(n_547), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_565), .B(n_583), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B(n_548), .C(n_551), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g763 ( .A(n_542), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_544), .A2(n_637), .B(n_684), .C(n_686), .Y(n_683) );
INVx8_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g669 ( .A(n_545), .Y(n_669) );
INVx3_ASAP7_75t_L g1002 ( .A(n_545), .Y(n_1002) );
INVx2_ASAP7_75t_L g1299 ( .A(n_545), .Y(n_1299) );
OAI211xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_556), .C(n_561), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_552), .A2(n_570), .B1(n_605), .B2(n_608), .C(n_609), .Y(n_604) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g762 ( .A(n_555), .Y(n_762) );
INVx3_ASAP7_75t_L g1101 ( .A(n_555), .Y(n_1101) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_558), .A2(n_728), .B1(n_743), .B2(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g769 ( .A(n_563), .Y(n_769) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_569), .A2(n_573), .B1(n_707), .B2(n_708), .Y(n_706) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_569), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_571), .A2(n_693), .B1(n_836), .B2(n_837), .Y(n_835) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_571), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_571), .A2(n_762), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_573), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_578), .B2(n_582), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_577), .A2(n_593), .B1(n_596), .B2(n_597), .C(n_598), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g1372 ( .A1(n_578), .A2(n_1356), .B1(n_1373), .B2(n_1375), .C(n_1376), .Y(n_1372) );
OAI221xp5_ASAP7_75t_L g1669 ( .A1(n_578), .A2(n_1670), .B1(n_1671), .B2(n_1672), .C(n_1673), .Y(n_1669) );
CKINVDCx8_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g776 ( .A(n_579), .Y(n_776) );
INVx3_ASAP7_75t_L g800 ( .A(n_579), .Y(n_800) );
INVx1_ASAP7_75t_L g1405 ( .A(n_579), .Y(n_1405) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g682 ( .A(n_580), .Y(n_682) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx2_ASAP7_75t_L g700 ( .A(n_581), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g1685 ( .A1(n_583), .A2(n_1686), .B(n_1698), .Y(n_1685) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_SL g1084 ( .A1(n_584), .A2(n_1085), .B(n_1104), .C(n_1109), .Y(n_1084) );
INVx1_ASAP7_75t_L g1265 ( .A(n_584), .Y(n_1265) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_585), .Y(n_809) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_585), .Y(n_1207) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_603), .C(n_616), .Y(n_586) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_593), .A2(n_839), .B1(n_844), .B2(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g735 ( .A(n_594), .Y(n_735) );
INVx2_ASAP7_75t_L g823 ( .A(n_594), .Y(n_823) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g607 ( .A(n_595), .Y(n_607) );
BUFx3_ASAP7_75t_L g819 ( .A(n_595), .Y(n_819) );
INVx1_ASAP7_75t_L g1123 ( .A(n_595), .Y(n_1123) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_595), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_597), .A2(n_791), .B1(n_799), .B2(n_819), .C(n_820), .Y(n_818) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g962 ( .A(n_600), .Y(n_962) );
INVx1_ASAP7_75t_L g1054 ( .A(n_600), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1174 ( .A(n_600), .Y(n_1174) );
INVx1_ASAP7_75t_L g1360 ( .A(n_600), .Y(n_1360) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g1188 ( .A(n_602), .Y(n_1188) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g634 ( .A(n_606), .Y(n_634) );
INVx4_ASAP7_75t_L g731 ( .A(n_606), .Y(n_731) );
INVx4_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_608), .A2(n_837), .B1(n_855), .B2(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_612), .Y(n_664) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x4_ASAP7_75t_L g977 ( .A(n_619), .B(n_681), .Y(n_977) );
INVx1_ASAP7_75t_L g1741 ( .A(n_619), .Y(n_1741) );
AOI21xp5_ASAP7_75t_SL g629 ( .A1(n_621), .A2(n_630), .B(n_651), .Y(n_629) );
BUFx2_ASAP7_75t_L g778 ( .A(n_621), .Y(n_778) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_665), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_639), .B(n_640), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g1748 ( .A1(n_632), .A2(n_1749), .B1(n_1750), .B2(n_1751), .Y(n_1748) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_633), .Y(n_1062) );
INVx4_ASAP7_75t_L g1329 ( .A(n_633), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_634), .A2(n_1402), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_636), .Y(n_963) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_636), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_636), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2x1_ASAP7_75t_L g954 ( .A(n_644), .B(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g1243 ( .A1(n_646), .A2(n_1244), .B1(n_1248), .B2(n_1249), .C1(n_1250), .C2(n_1252), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_649), .B(n_1662), .Y(n_1700) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_650), .A2(n_673), .B1(n_674), .B2(n_677), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_660), .B1(n_661), .B2(n_663), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g1050 ( .A(n_654), .Y(n_1050) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_655), .Y(n_1059) );
INVx1_ASAP7_75t_L g1258 ( .A(n_655), .Y(n_1258) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g1693 ( .A(n_656), .Y(n_1693) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g944 ( .A(n_659), .Y(n_944) );
INVx2_ASAP7_75t_L g1206 ( .A(n_659), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_664), .Y(n_1186) );
NAND3xp33_ASAP7_75t_SL g665 ( .A(n_666), .B(n_672), .C(n_679), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_668), .A2(n_967), .B1(n_970), .B2(n_974), .Y(n_973) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AND2x4_ASAP7_75t_L g1390 ( .A(n_669), .B(n_670), .Y(n_1390) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g676 ( .A(n_671), .Y(n_676) );
OR2x2_ASAP7_75t_L g681 ( .A(n_671), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx2_ASAP7_75t_L g703 ( .A(n_675), .Y(n_703) );
INVx2_ASAP7_75t_L g805 ( .A(n_675), .Y(n_805) );
INVxp67_ASAP7_75t_L g1229 ( .A(n_676), .Y(n_1229) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_687), .Y(n_679) );
BUFx3_ASAP7_75t_L g845 ( .A(n_682), .Y(n_845) );
INVx1_ASAP7_75t_L g1097 ( .A(n_682), .Y(n_1097) );
INVx2_ASAP7_75t_L g985 ( .A(n_685), .Y(n_985) );
AND2x4_ASAP7_75t_L g984 ( .A(n_686), .B(n_985), .Y(n_984) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_686), .B(n_995), .Y(n_1005) );
AND2x4_ASAP7_75t_SL g1384 ( .A(n_686), .B(n_985), .Y(n_1384) );
OAI33xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .A3(n_694), .B1(n_702), .B2(n_706), .B3(n_709), .Y(n_687) );
BUFx3_ASAP7_75t_L g1675 ( .A(n_688), .Y(n_1675) );
BUFx4f_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g834 ( .A(n_689), .Y(n_834) );
BUFx8_ASAP7_75t_L g1272 ( .A(n_689), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_701), .Y(n_694) );
INVx8_ASAP7_75t_L g997 ( .A(n_696), .Y(n_997) );
INVx5_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g798 ( .A(n_697), .Y(n_798) );
INVx2_ASAP7_75t_SL g1302 ( .A(n_697), .Y(n_1302) );
INVx2_ASAP7_75t_SL g1726 ( .A(n_697), .Y(n_1726) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_698), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g1370 ( .A(n_699), .Y(n_1370) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_700), .Y(n_1279) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_828), .B1(n_829), .B2(n_1006), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1006 ( .A(n_715), .Y(n_1006) );
XNOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_781), .Y(n_715) );
XNOR2x1_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_758), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_750), .C(n_756), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_746), .Y(n_720) );
OAI33xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .A3(n_727), .B1(n_733), .B2(n_739), .B3(n_744), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_722), .A2(n_818), .B1(n_821), .B2(n_822), .Y(n_817) );
OAI33xp33_ASAP7_75t_L g1114 ( .A1(n_722), .A2(n_1115), .A3(n_1120), .B1(n_1124), .B2(n_1126), .B3(n_1128), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_726), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_739) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_726), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_726), .A2(n_1332), .B1(n_1333), .B2(n_1335), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_727) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_729), .Y(n_864) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g1429 ( .A(n_730), .Y(n_1429) );
INVx2_ASAP7_75t_L g1755 ( .A(n_730), .Y(n_1755) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_734), .A2(n_1410), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
INVx4_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_737), .A2(n_1095), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
OAI211xp5_ASAP7_75t_L g1690 ( .A1(n_737), .A2(n_1691), .B(n_1692), .C(n_1694), .Y(n_1690) );
OAI211xp5_ASAP7_75t_SL g1695 ( .A1(n_737), .A2(n_1677), .B(n_1696), .C(n_1697), .Y(n_1695) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g1128 ( .A(n_745), .Y(n_1128) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g1161 ( .A1(n_753), .A2(n_827), .B(n_1144), .Y(n_1161) );
AOI21xp5_ASAP7_75t_L g1338 ( .A1(n_753), .A2(n_827), .B(n_1339), .Y(n_1338) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_765), .B(n_777), .C(n_779), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g1403 ( .A1(n_761), .A2(n_1404), .B1(n_1405), .B2(n_1406), .Y(n_1403) );
NOR3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .C(n_772), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_766), .B(n_787), .C(n_793), .Y(n_786) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_776), .A2(n_1151), .B1(n_1152), .B2(n_1153), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1676 ( .A1(n_776), .A2(n_843), .B1(n_1677), .B2(n_1678), .C(n_1679), .Y(n_1676) );
A2O1A1Ixp33_ASAP7_75t_L g1295 ( .A1(n_777), .A2(n_1296), .B(n_1309), .C(n_1313), .Y(n_1295) );
INVx1_ASAP7_75t_L g1412 ( .A(n_777), .Y(n_1412) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI31xp33_ASAP7_75t_SL g1017 ( .A1(n_778), .A2(n_1018), .A3(n_1019), .B(n_1024), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1717 ( .A1(n_778), .A2(n_1718), .B(n_1737), .Y(n_1717) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
XNOR2x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
OR2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_811), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_802), .B(n_809), .C(n_810), .Y(n_785) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_788), .Y(n_1223) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_790), .A2(n_795), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_800), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_838) );
OAI21xp33_ASAP7_75t_L g1342 ( .A1(n_809), .A2(n_1343), .B(n_1353), .Y(n_1342) );
INVx1_ASAP7_75t_L g1315 ( .A(n_812), .Y(n_1315) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_826), .C(n_827), .Y(n_816) );
INVx2_ASAP7_75t_L g867 ( .A(n_819), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_821), .Y(n_869) );
OAI221xp5_ASAP7_75t_L g938 ( .A1(n_823), .A2(n_939), .B1(n_941), .B2(n_942), .C(n_943), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_824), .A2(n_1090), .B1(n_1100), .B2(n_1125), .Y(n_1124) );
OR3x1_ASAP7_75t_L g1419 ( .A(n_827), .B(n_1420), .C(n_1421), .Y(n_1419) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_930), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_873), .C(n_900), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_856), .Y(n_832) );
OAI33xp33_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .A3(n_838), .B1(n_842), .B2(n_847), .B3(n_852), .Y(n_833) );
OAI22xp5_ASAP7_75t_SL g857 ( .A1(n_836), .A2(n_853), .B1(n_858), .B2(n_861), .Y(n_857) );
INVx1_ASAP7_75t_L g1034 ( .A(n_840), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_841), .A2(n_846), .B1(n_858), .B2(n_871), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_845), .A2(n_1026), .B1(n_1029), .B2(n_1030), .C(n_1031), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_845), .A2(n_1036), .B1(n_1038), .B2(n_1039), .C(n_1040), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_845), .A2(n_1268), .B1(n_1269), .B2(n_1271), .Y(n_1267) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AOI33xp33_ASAP7_75t_L g990 ( .A1(n_848), .A2(n_991), .A3(n_993), .B1(n_996), .B2(n_999), .B3(n_1001), .Y(n_990) );
BUFx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_849), .Y(n_1283) );
INVx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx3_ASAP7_75t_L g1225 ( .A(n_850), .Y(n_1225) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g872 ( .A(n_862), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g1327 ( .A1(n_862), .A2(n_1308), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
OAI221xp5_ASAP7_75t_L g1753 ( .A1(n_866), .A2(n_1754), .B1(n_1755), .B2(n_1756), .C(n_1757), .Y(n_1753) );
INVx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI31xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_886), .A3(n_893), .B(n_897), .Y(n_873) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_880), .B1(n_882), .B2(n_883), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_879), .A2(n_910), .B1(n_914), .B2(n_917), .Y(n_909) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx3_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
BUFx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
OAI31xp33_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_906), .A3(n_918), .B(n_924), .Y(n_900) );
INVx2_ASAP7_75t_SL g1665 ( .A(n_902), .Y(n_1665) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1654 ( .A1(n_904), .A2(n_1655), .B1(n_1656), .B2(n_1657), .Y(n_1654) );
NAND4xp25_ASAP7_75t_L g1653 ( .A(n_907), .B(n_1654), .C(n_1658), .D(n_1663), .Y(n_1653) );
CKINVDCx8_ASAP7_75t_R g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
BUFx3_ASAP7_75t_L g1660 ( .A(n_911), .Y(n_1660) );
AND2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
AND2x4_ASAP7_75t_L g915 ( .A(n_912), .B(n_916), .Y(n_915) );
AOI222xp33_ASAP7_75t_L g1658 ( .A1(n_914), .A2(n_1003), .B1(n_1659), .B2(n_1660), .C1(n_1661), .C2(n_1662), .Y(n_1658) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1663 ( .A1(n_920), .A2(n_1664), .B1(n_1665), .B2(n_1666), .Y(n_1663) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
BUFx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g1657 ( .A(n_923), .Y(n_1657) );
BUFx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AND2x2_ASAP7_75t_SL g925 ( .A(n_926), .B(n_928), .Y(n_925) );
AND2x4_ASAP7_75t_L g1667 ( .A(n_926), .B(n_928), .Y(n_1667) );
INVx1_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NAND3x1_ASAP7_75t_L g931 ( .A(n_932), .B(n_975), .C(n_979), .Y(n_931) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g1354 ( .A(n_935), .Y(n_1354) );
INVx4_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
BUFx3_ASAP7_75t_L g1254 ( .A(n_937), .Y(n_1254) );
INVx5_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_949), .B2(n_952), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_947), .A2(n_1098), .B1(n_1119), .B2(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
BUFx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx2_ASAP7_75t_L g1197 ( .A(n_954), .Y(n_1197) );
INVx3_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g1261 ( .A1(n_958), .A2(n_968), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B(n_964), .Y(n_959) );
AOI21xp5_ASAP7_75t_L g1181 ( .A1(n_964), .A2(n_1182), .B(n_1185), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_964), .A2(n_1254), .B1(n_1255), .B2(n_1256), .C(n_1259), .Y(n_1253) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_964), .A2(n_1350), .B(n_1352), .Y(n_1349) );
AOI211xp5_ASAP7_75t_SL g1698 ( .A1(n_964), .A2(n_1254), .B(n_1661), .C(n_1699), .Y(n_1698) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_970), .Y(n_965) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_966), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_966), .A2(n_969), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
INVx1_ASAP7_75t_L g1688 ( .A(n_966), .Y(n_1688) );
BUFx6f_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g1194 ( .A(n_969), .Y(n_1194) );
INVx2_ASAP7_75t_L g1240 ( .A(n_972), .Y(n_1240) );
INVx2_ASAP7_75t_L g1230 ( .A(n_974), .Y(n_1230) );
INVx2_ASAP7_75t_L g1284 ( .A(n_974), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_974), .A2(n_1347), .B1(n_1348), .B2(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g1208 ( .A1(n_976), .A2(n_1209), .B(n_1210), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g1285 ( .A1(n_976), .A2(n_1263), .B1(n_1286), .B2(n_1287), .C(n_1288), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g1385 ( .A1(n_976), .A2(n_1386), .B(n_1387), .Y(n_1385) );
INVx8_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
AND4x1_ASAP7_75t_SL g979 ( .A(n_980), .B(n_986), .C(n_990), .D(n_1004), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_982), .A2(n_984), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_984), .A2(n_1249), .B1(n_1255), .B2(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
INVx5_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx3_ASAP7_75t_L g1286 ( .A(n_989), .Y(n_1286) );
AOI33xp33_ASAP7_75t_L g1216 ( .A1(n_991), .A2(n_1217), .A3(n_1220), .B1(n_1224), .B2(n_1225), .B3(n_1226), .Y(n_1216) );
BUFx3_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
BUFx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1003), .Y(n_1683) );
INVx3_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx3_ASAP7_75t_L g1232 ( .A(n_1005), .Y(n_1232) );
NOR3xp33_ASAP7_75t_L g1362 ( .A(n_1005), .B(n_1363), .C(n_1380), .Y(n_1362) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
XNOR2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1234), .Y(n_1009) );
OA22x2_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1079), .B1(n_1080), .B2(n_1233), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1012), .Y(n_1233) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NOR2x1_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1047), .Y(n_1014) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1016), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1035), .C(n_1044), .Y(n_1024) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
OR2x6_ASAP7_75t_L g1228 ( .A(n_1028), .B(n_1229), .Y(n_1228) );
OAI22xp5_ASAP7_75t_SL g1060 ( .A1(n_1029), .A2(n_1061), .B1(n_1063), .B2(n_1064), .Y(n_1060) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_1033), .A2(n_1299), .B1(n_1734), .B2(n_1735), .Y(n_1733) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1037), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1068), .Y(n_1047) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1055 ( .A(n_1056), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1198 ( .A1(n_1061), .A2(n_1199), .B1(n_1200), .B2(n_1201), .C(n_1202), .Y(n_1198) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx3_ASAP7_75t_L g1426 ( .A(n_1062), .Y(n_1426) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
BUFx6f_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
AOI21xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B(n_1072), .Y(n_1068) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
XNOR2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1177), .Y(n_1080) );
XNOR2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1133), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1112), .Y(n_1083) );
OAI21xp33_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1093), .B(n_1099), .Y(n_1088) );
OAI21xp33_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B(n_1092), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1096), .B2(n_1098), .Y(n_1093) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1094), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1096), .A2(n_1148), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1101), .B(n_1102), .C(n_1103), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
NAND3xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1130), .C(n_1132), .Y(n_1112) );
NOR2xp33_ASAP7_75t_SL g1113 ( .A(n_1114), .B(n_1129), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1117), .B1(n_1118), .B2(n_1119), .Y(n_1115) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
XOR2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1176), .Y(n_1133) );
NOR2xp33_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1160), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1150), .B1(n_1154), .B2(n_1157), .Y(n_1145) );
OAI21xp5_ASAP7_75t_L g1364 ( .A1(n_1148), .A2(n_1365), .B(n_1366), .Y(n_1364) );
NAND4xp25_ASAP7_75t_SL g1160 ( .A(n_1161), .B(n_1162), .C(n_1164), .D(n_1167), .Y(n_1160) );
NAND3xp33_ASAP7_75t_SL g1178 ( .A(n_1179), .B(n_1208), .C(n_1211), .Y(n_1178) );
OAI21xp33_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1195), .B(n_1207), .Y(n_1179) );
HB1xp67_ASAP7_75t_SL g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B1(n_1192), .B2(n_1193), .Y(n_1189) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NOR3xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1227), .C(n_1231), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1216), .Y(n_1212) );
BUFx2_ASAP7_75t_SL g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g1379 ( .A(n_1225), .Y(n_1379) );
INVx2_ASAP7_75t_L g1684 ( .A(n_1225), .Y(n_1684) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_1232), .Y(n_1231) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_1235), .A2(n_1391), .B1(n_1392), .B2(n_1432), .Y(n_1234) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1235), .Y(n_1432) );
XOR2xp5_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1292), .Y(n_1235) );
XNOR2x1_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1238), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1285), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1241), .B1(n_1242), .B2(n_1264), .C(n_1266), .Y(n_1239) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1253), .C(n_1261), .Y(n_1242) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1247), .Y(n_1351) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1270), .Y(n_1670) );
CKINVDCx20_ASAP7_75t_R g1366 ( .A(n_1272), .Y(n_1366) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1278), .B1(n_1279), .B2(n_1280), .C(n_1281), .Y(n_1276) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
XNOR2xp5_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1340), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1316), .Y(n_1294) );
NOR3xp33_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .C(n_1304), .Y(n_1296) );
INVx2_ASAP7_75t_L g1723 ( .A(n_1302), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
NAND4xp25_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .C(n_1336), .D(n_1338), .Y(n_1316) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AND4x1_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1362), .C(n_1385), .D(n_1389), .Y(n_1341) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B(n_1358), .C(n_1359), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1367), .B1(n_1372), .B2(n_1379), .Y(n_1363) );
OAI21xp33_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1369), .B(n_1371), .Y(n_1367) );
INVx3_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1378), .Y(n_1674) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
AOI211x1_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1412), .B(n_1413), .C(n_1419), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1399), .Y(n_1394) );
NOR3xp33_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1407), .C(n_1408), .Y(n_1399) );
OAI221xp5_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1644), .B1(n_1648), .B2(n_1702), .C(n_1707), .Y(n_1433) );
AOI21xp5_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1557), .B(n_1601), .Y(n_1434) );
OAI211xp5_ASAP7_75t_L g1435 ( .A1(n_1436), .A2(n_1451), .B(n_1497), .C(n_1543), .Y(n_1435) );
AOI22xp5_ASAP7_75t_L g1626 ( .A1(n_1436), .A2(n_1549), .B1(n_1627), .B2(n_1633), .Y(n_1626) );
CKINVDCx5p33_ASAP7_75t_R g1436 ( .A(n_1437), .Y(n_1436) );
CKINVDCx6p67_ASAP7_75t_R g1509 ( .A(n_1437), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1437), .B(n_1469), .Y(n_1610) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1437), .B(n_1469), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1437), .B(n_1533), .Y(n_1643) );
OR2x6_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1445), .Y(n_1437) );
OR2x2_ASAP7_75t_L g1530 ( .A(n_1438), .B(n_1445), .Y(n_1530) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1439), .Y(n_1540) );
AND2x6_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1440), .B(n_1444), .Y(n_1443) );
AND2x4_ASAP7_75t_L g1446 ( .A(n_1440), .B(n_1447), .Y(n_1446) );
AND2x6_ASAP7_75t_L g1449 ( .A(n_1440), .B(n_1450), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1440), .B(n_1444), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1440), .B(n_1444), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1442), .B(n_1448), .Y(n_1447) );
OAI21xp5_ASAP7_75t_L g1761 ( .A1(n_1444), .A2(n_1762), .B(n_1763), .Y(n_1761) );
O2A1O1Ixp33_ASAP7_75t_L g1451 ( .A1(n_1452), .A2(n_1467), .B(n_1472), .C(n_1486), .Y(n_1451) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1457), .Y(n_1452) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1453), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1453), .B(n_1488), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1453), .B(n_1462), .Y(n_1494) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1453), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1453), .B(n_1525), .Y(n_1524) );
OR2x2_ASAP7_75t_L g1567 ( .A(n_1453), .B(n_1529), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1453), .B(n_1482), .Y(n_1599) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1453), .B(n_1482), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1455), .Y(n_1453) );
INVxp67_ASAP7_75t_L g1542 ( .A(n_1456), .Y(n_1542) );
HB1xp67_ASAP7_75t_L g1647 ( .A(n_1456), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1462), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1458), .B(n_1491), .Y(n_1496) );
AND3x1_ASAP7_75t_L g1513 ( .A(n_1458), .B(n_1474), .C(n_1479), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1458), .B(n_1474), .Y(n_1520) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1458), .B(n_1462), .Y(n_1632) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1459), .B(n_1474), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1459), .B(n_1491), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1459), .B(n_1462), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1461), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1462), .B(n_1491), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_1462), .B(n_1474), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1462), .B(n_1520), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1462), .B(n_1474), .Y(n_1597) );
BUFx2_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx2_ASAP7_75t_L g1479 ( .A(n_1463), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1463), .B(n_1473), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1463), .B(n_1496), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1463), .B(n_1504), .Y(n_1564) );
OR2x2_ASAP7_75t_L g1585 ( .A(n_1463), .B(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
O2A1O1Ixp33_ASAP7_75t_L g1472 ( .A1(n_1467), .A2(n_1473), .B(n_1477), .C(n_1481), .Y(n_1472) );
CKINVDCx14_ASAP7_75t_R g1467 ( .A(n_1468), .Y(n_1467) );
OAI22xp5_ASAP7_75t_L g1550 ( .A1(n_1468), .A2(n_1548), .B1(n_1551), .B2(n_1554), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1468), .B(n_1536), .Y(n_1568) );
AOI211xp5_ASAP7_75t_L g1592 ( .A1(n_1468), .A2(n_1593), .B(n_1594), .C(n_1595), .Y(n_1592) );
AOI221xp5_ASAP7_75t_L g1602 ( .A1(n_1468), .A2(n_1513), .B1(n_1603), .B2(n_1605), .C(n_1606), .Y(n_1602) );
INVx3_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1469), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1469), .B(n_1482), .Y(n_1499) );
AOI22xp5_ASAP7_75t_L g1523 ( .A1(n_1469), .A2(n_1524), .B1(n_1527), .B2(n_1528), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1469), .B(n_1482), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1469), .B(n_1488), .Y(n_1534) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1469), .B(n_1509), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1469), .B(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1469), .B(n_1509), .Y(n_1625) );
AND2x4_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1471), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_1473), .B(n_1480), .Y(n_1547) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1473), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1473), .B(n_1494), .Y(n_1630) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1474), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1526 ( .A(n_1474), .B(n_1479), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1476), .Y(n_1474) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1478), .B(n_1496), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1480), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1479), .B(n_1504), .Y(n_1503) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1479), .B(n_1547), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1479), .B(n_1496), .Y(n_1589) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1479), .B(n_1556), .Y(n_1638) );
NAND2xp5_ASAP7_75t_SL g1640 ( .A(n_1479), .B(n_1641), .Y(n_1640) );
NOR2xp33_ASAP7_75t_L g1518 ( .A(n_1480), .B(n_1519), .Y(n_1518) );
NOR2xp33_ASAP7_75t_L g1553 ( .A(n_1480), .B(n_1515), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1480), .B(n_1508), .Y(n_1563) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1480), .Y(n_1591) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1480), .B(n_1597), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1481), .B(n_1509), .Y(n_1516) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1481), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1485), .Y(n_1481) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1482), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1484), .Y(n_1482) );
OAI21xp33_ASAP7_75t_L g1486 ( .A1(n_1487), .A2(n_1489), .B(n_1492), .Y(n_1486) );
INVx2_ASAP7_75t_L g1508 ( .A(n_1488), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1488), .B(n_1509), .Y(n_1521) );
OAI211xp5_ASAP7_75t_SL g1559 ( .A1(n_1489), .A2(n_1560), .B(n_1561), .C(n_1565), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1489), .B(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
A2O1A1Ixp33_ASAP7_75t_L g1517 ( .A1(n_1490), .A2(n_1502), .B(n_1518), .C(n_1521), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_1490), .A2(n_1544), .B1(n_1545), .B2(n_1548), .C(n_1550), .Y(n_1543) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1492), .Y(n_1593) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1492), .B(n_1508), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1495), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1496), .B(n_1502), .Y(n_1556) );
AOI211xp5_ASAP7_75t_L g1497 ( .A1(n_1498), .A2(n_1500), .B(n_1505), .C(n_1522), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1498), .B(n_1502), .Y(n_1544) );
OAI322xp33_ASAP7_75t_L g1571 ( .A1(n_1498), .A2(n_1515), .A3(n_1530), .B1(n_1547), .B2(n_1572), .C1(n_1575), .C2(n_1577), .Y(n_1571) );
AND2x2_ASAP7_75t_SL g1594 ( .A(n_1498), .B(n_1513), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1498), .B(n_1501), .Y(n_1604) );
INVx2_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1503), .Y(n_1500) );
NOR2xp33_ASAP7_75t_L g1514 ( .A(n_1501), .B(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1501), .Y(n_1576) );
AOI31xp33_ASAP7_75t_L g1583 ( .A1(n_1501), .A2(n_1579), .A3(n_1584), .B(n_1587), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1501), .B(n_1513), .Y(n_1624) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
NAND2xp5_ASAP7_75t_SL g1560 ( .A(n_1502), .B(n_1527), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1502), .B(n_1582), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1503), .B(n_1576), .Y(n_1575) );
OR2x2_ASAP7_75t_L g1641 ( .A(n_1504), .B(n_1520), .Y(n_1641) );
OAI211xp5_ASAP7_75t_L g1505 ( .A1(n_1506), .A2(n_1510), .B(n_1512), .C(n_1517), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1509), .Y(n_1507) );
INVx2_ASAP7_75t_L g1549 ( .A(n_1508), .Y(n_1549) );
A2O1A1Ixp33_ASAP7_75t_L g1621 ( .A1(n_1508), .A2(n_1622), .B(n_1624), .C(n_1625), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1509), .B(n_1570), .Y(n_1569) );
NOR2xp33_ASAP7_75t_SL g1573 ( .A(n_1509), .B(n_1574), .Y(n_1573) );
NOR2xp33_ASAP7_75t_L g1615 ( .A(n_1509), .B(n_1616), .Y(n_1615) );
O2A1O1Ixp33_ASAP7_75t_L g1606 ( .A1(n_1510), .A2(n_1607), .B(n_1608), .C(n_1609), .Y(n_1606) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
OAI21xp33_ASAP7_75t_L g1512 ( .A1(n_1513), .A2(n_1514), .B(n_1516), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1516), .B(n_1532), .Y(n_1600) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1521), .Y(n_1577) );
OAI221xp5_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1530), .B1(n_1531), .B2(n_1533), .C(n_1535), .Y(n_1522) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_1530), .A2(n_1612), .B1(n_1617), .B2(n_1619), .Y(n_1611) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
CKINVDCx6p67_ASAP7_75t_R g1533 ( .A(n_1534), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1534), .B(n_1591), .Y(n_1590) );
INVx3_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVx2_ASAP7_75t_SL g1536 ( .A(n_1537), .Y(n_1536) );
OAI21xp33_ASAP7_75t_L g1565 ( .A1(n_1537), .A2(n_1566), .B(n_1568), .Y(n_1565) );
INVx2_ASAP7_75t_SL g1570 ( .A(n_1537), .Y(n_1570) );
OAI22xp5_ASAP7_75t_SL g1538 ( .A1(n_1539), .A2(n_1540), .B1(n_1541), .B2(n_1542), .Y(n_1538) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1544), .Y(n_1613) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1548), .B(n_1553), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1548), .B(n_1593), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1548), .B(n_1635), .Y(n_1634) );
INVx2_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
NAND5xp2_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1578), .C(n_1583), .D(n_1592), .E(n_1600), .Y(n_1557) );
AOI21xp5_ASAP7_75t_L g1558 ( .A1(n_1559), .A2(n_1569), .B(n_1571), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1564), .Y(n_1561) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
NAND3xp33_ASAP7_75t_L g1622 ( .A(n_1567), .B(n_1588), .C(n_1623), .Y(n_1622) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1581), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
OAI22xp5_ASAP7_75t_L g1627 ( .A1(n_1580), .A2(n_1628), .B1(n_1629), .B2(n_1631), .Y(n_1627) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1582), .Y(n_1618) );
AOI21xp33_ASAP7_75t_L g1587 ( .A1(n_1586), .A2(n_1588), .B(n_1590), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1588), .B(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
INVxp67_ASAP7_75t_SL g1595 ( .A(n_1596), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1598), .Y(n_1596) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1597), .Y(n_1607) );
CKINVDCx14_ASAP7_75t_R g1608 ( .A(n_1599), .Y(n_1608) );
NAND5xp2_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1611), .C(n_1621), .D(n_1626), .E(n_1636), .Y(n_1601) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_SL g1612 ( .A(n_1613), .B(n_1614), .Y(n_1612) );
INVxp67_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
CKINVDCx14_ASAP7_75t_R g1631 ( .A(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
OAI21xp5_ASAP7_75t_L g1636 ( .A1(n_1637), .A2(n_1639), .B(n_1642), .Y(n_1636) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVxp67_ASAP7_75t_SL g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
CKINVDCx20_ASAP7_75t_R g1644 ( .A(n_1645), .Y(n_1644) );
CKINVDCx20_ASAP7_75t_R g1645 ( .A(n_1646), .Y(n_1645) );
INVx4_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
HB1xp67_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
AOI211xp5_ASAP7_75t_L g1652 ( .A1(n_1653), .A2(n_1667), .B(n_1668), .C(n_1685), .Y(n_1652) );
OAI22xp5_ASAP7_75t_L g1668 ( .A1(n_1669), .A2(n_1675), .B1(n_1676), .B2(n_1684), .Y(n_1668) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
NOR2xp33_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1689), .Y(n_1686) );
CKINVDCx20_ASAP7_75t_R g1702 ( .A(n_1703), .Y(n_1702) );
CKINVDCx20_ASAP7_75t_R g1703 ( .A(n_1704), .Y(n_1703) );
INVx3_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
HB1xp67_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
BUFx3_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVxp33_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
HB1xp67_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
AND3x1_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1738), .C(n_1746), .Y(n_1716) );
NAND3xp33_ASAP7_75t_SL g1718 ( .A(n_1719), .B(n_1728), .C(n_1731), .Y(n_1718) );
AOI22xp5_ASAP7_75t_L g1719 ( .A1(n_1720), .A2(n_1722), .B1(n_1724), .B2(n_1727), .Y(n_1719) );
INVx2_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1739), .B(n_1743), .Y(n_1738) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
endmodule