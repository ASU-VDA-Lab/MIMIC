module fake_netlist_5_1346_n_67 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_67);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_67;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_28;
wire n_46;
wire n_24;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_38;
wire n_61;
wire n_35;
wire n_41;
wire n_32;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_20;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_49;
wire n_52;
wire n_60;
wire n_39;

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_5),
.B(n_13),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_6),
.B(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_19),
.B(n_21),
.C(n_31),
.Y(n_44)
);

OR2x6_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_51),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_50),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_47),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_45),
.C(n_44),
.Y(n_59)
);

OAI31xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_34),
.A3(n_48),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_45),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_57),
.Y(n_62)
);

AOI221xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.C(n_27),
.Y(n_63)
);

NAND4xp25_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_60),
.C(n_25),
.D(n_22),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_62),
.B(n_22),
.Y(n_65)
);

AOI222xp33_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.C1(n_23),
.C2(n_32),
.Y(n_66)
);

OR2x6_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_29),
.Y(n_67)
);


endmodule