module real_aes_6242_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_0), .A2(n_222), .B(n_226), .C(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_1), .A2(n_217), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g520 ( .A(n_1), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_2), .B(n_240), .Y(n_293) );
INVx1_ASAP7_75t_L g200 ( .A(n_3), .Y(n_200) );
AND2x6_ASAP7_75t_L g222 ( .A(n_3), .B(n_198), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_3), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g250 ( .A(n_4), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_5), .B(n_231), .Y(n_267) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_6), .A2(n_25), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g215 ( .A(n_7), .Y(n_215) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_8), .A2(n_72), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_8), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_9), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_10), .A2(n_251), .B(n_276), .C(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_11), .B(n_240), .Y(n_279) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_12), .A2(n_28), .B1(n_89), .B2(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_13), .B(n_336), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_14), .A2(n_230), .B(n_232), .C(n_236), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_15), .B(n_231), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_16), .A2(n_80), .B1(n_177), .B2(n_178), .Y(n_79) );
INVx1_ASAP7_75t_L g177 ( .A(n_16), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_16), .B(n_231), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_17), .Y(n_296) );
INVx1_ASAP7_75t_L g310 ( .A(n_18), .Y(n_310) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_19), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_20), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_21), .A2(n_80), .B1(n_178), .B2(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_21), .Y(n_522) );
INVx1_ASAP7_75t_L g333 ( .A(n_22), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_23), .A2(n_180), .B1(n_186), .B2(n_187), .Y(n_179) );
INVx1_ASAP7_75t_L g186 ( .A(n_23), .Y(n_186) );
INVx2_ASAP7_75t_L g220 ( .A(n_24), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_26), .A2(n_44), .B1(n_170), .B2(n_174), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_27), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g191 ( .A1(n_28), .A2(n_41), .B1(n_52), .B2(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_28), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_29), .A2(n_230), .B(n_289), .C(n_291), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_30), .Y(n_150) );
INVxp67_ASAP7_75t_L g334 ( .A(n_31), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g287 ( .A(n_32), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_33), .A2(n_226), .B(n_309), .C(n_315), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_34), .A2(n_49), .B1(n_152), .B2(n_157), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_35), .Y(n_83) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_36), .A2(n_248), .B(n_249), .C(n_252), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_37), .A2(n_181), .B1(n_182), .B2(n_185), .Y(n_180) );
INVx1_ASAP7_75t_L g185 ( .A(n_37), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_38), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_39), .Y(n_330) );
INVx1_ASAP7_75t_L g224 ( .A(n_40), .Y(n_224) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_41), .A2(n_63), .B1(n_89), .B2(n_93), .Y(n_98) );
INVxp67_ASAP7_75t_L g195 ( .A(n_41), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g246 ( .A(n_42), .Y(n_246) );
INVx1_ASAP7_75t_L g198 ( .A(n_43), .Y(n_198) );
INVx1_ASAP7_75t_L g214 ( .A(n_45), .Y(n_214) );
INVx1_ASAP7_75t_SL g290 ( .A(n_46), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_46), .A2(n_80), .B1(n_178), .B2(n_290), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_47), .A2(n_67), .B1(n_163), .B2(n_167), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_48), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_50), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g299 ( .A(n_51), .Y(n_299) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_52), .A2(n_71), .B1(n_89), .B2(n_90), .Y(n_96) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_53), .A2(n_217), .B(n_245), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_54), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_55), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_56), .A2(n_217), .B(n_273), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_57), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_58), .A2(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g274 ( .A(n_59), .Y(n_274) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_60), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_61), .A2(n_217), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g277 ( .A(n_62), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_64), .Y(n_125) );
INVx2_ASAP7_75t_L g212 ( .A(n_65), .Y(n_212) );
INVx1_ASAP7_75t_L g264 ( .A(n_66), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_68), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_69), .A2(n_226), .B(n_298), .C(n_301), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_70), .Y(n_113) );
INVx1_ASAP7_75t_L g184 ( .A(n_72), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_73), .B(n_210), .Y(n_254) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx2_ASAP7_75t_L g233 ( .A(n_75), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_76), .Y(n_127) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_188), .B1(n_201), .B2(n_507), .C(n_510), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_179), .Y(n_78) );
INVx1_ASAP7_75t_L g178 ( .A(n_80), .Y(n_178) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_140), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_105), .C(n_126), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_99), .B2(n_100), .Y(n_82) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
INVx2_ASAP7_75t_L g166 ( .A(n_86), .Y(n_166) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g104 ( .A(n_87), .B(n_92), .Y(n_104) );
AND2x2_ASAP7_75t_L g145 ( .A(n_87), .B(n_111), .Y(n_145) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_98), .Y(n_112) );
AND2x2_ASAP7_75t_L g117 ( .A(n_88), .B(n_92), .Y(n_117) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
INVx1_ASAP7_75t_L g159 ( .A(n_92), .Y(n_159) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2x1p5_ASAP7_75t_L g103 ( .A(n_95), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g149 ( .A(n_95), .B(n_145), .Y(n_149) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g110 ( .A(n_96), .Y(n_110) );
INVx1_ASAP7_75t_L g119 ( .A(n_96), .Y(n_119) );
INVx1_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_96), .B(n_98), .Y(n_160) );
AND2x2_ASAP7_75t_L g118 ( .A(n_97), .B(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g156 ( .A(n_98), .B(n_139), .Y(n_156) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g155 ( .A(n_104), .B(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g168 ( .A(n_104), .B(n_118), .Y(n_168) );
OAI222xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_113), .B1(n_114), .B2(n_120), .C1(n_121), .C2(n_125), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
INVx1_ASAP7_75t_L g131 ( .A(n_111), .Y(n_131) );
AND2x4_ASAP7_75t_L g123 ( .A(n_112), .B(n_124), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g130 ( .A(n_112), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g136 ( .A(n_117), .Y(n_136) );
AND2x2_ASAP7_75t_L g144 ( .A(n_118), .B(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g165 ( .A(n_118), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_132), .B2(n_133), .Y(n_126) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_135), .Y(n_134) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_161), .Y(n_140) );
OAI221xp5_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_146), .B1(n_147), .B2(n_150), .C(n_151), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g173 ( .A(n_145), .B(n_156), .Y(n_173) );
AND2x4_ASAP7_75t_L g175 ( .A(n_145), .B(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_162), .B(n_169), .Y(n_161) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx11_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_180), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
AND3x1_ASAP7_75t_SL g190 ( .A(n_191), .B(n_196), .C(n_199), .Y(n_190) );
INVxp67_ASAP7_75t_L g515 ( .A(n_191), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_SL g517 ( .A(n_196), .Y(n_517) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_196), .A2(n_218), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g526 ( .A(n_196), .Y(n_526) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_197), .B(n_200), .Y(n_519) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_199), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_433), .Y(n_203) );
NOR4xp25_ASAP7_75t_L g204 ( .A(n_205), .B(n_375), .C(n_405), .D(n_415), .Y(n_204) );
OAI211xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_280), .B(n_338), .C(n_365), .Y(n_205) );
OAI222xp33_ASAP7_75t_L g460 ( .A1(n_206), .A2(n_380), .B1(n_461), .B2(n_462), .C1(n_463), .C2(n_464), .Y(n_460) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_255), .Y(n_206) );
AOI33xp33_ASAP7_75t_L g386 ( .A1(n_207), .A2(n_373), .A3(n_374), .B1(n_387), .B2(n_392), .B3(n_394), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g443 ( .A1(n_207), .A2(n_444), .B(n_446), .C(n_448), .Y(n_443) );
OR2x2_ASAP7_75t_L g459 ( .A(n_207), .B(n_445), .Y(n_459) );
INVx1_ASAP7_75t_L g492 ( .A(n_207), .Y(n_492) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_242), .Y(n_207) );
INVx2_ASAP7_75t_L g369 ( .A(n_208), .Y(n_369) );
AND2x2_ASAP7_75t_L g385 ( .A(n_208), .B(n_271), .Y(n_385) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_208), .Y(n_420) );
AND2x2_ASAP7_75t_L g449 ( .A(n_208), .B(n_242), .Y(n_449) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_216), .B(n_239), .Y(n_208) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_209), .A2(n_272), .B(n_279), .Y(n_271) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_209), .A2(n_285), .B(n_293), .Y(n_284) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx4_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g326 ( .A(n_211), .Y(n_326) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_212), .B(n_213), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx2_ASAP7_75t_L g328 ( .A(n_217), .Y(n_328) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_222), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_218), .B(n_222), .Y(n_261) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g314 ( .A(n_219), .Y(n_314) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
INVx1_ASAP7_75t_L g237 ( .A(n_220), .Y(n_237) );
INVx1_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_221), .Y(n_235) );
INVx3_ASAP7_75t_L g251 ( .A(n_221), .Y(n_251) );
INVx4_ASAP7_75t_SL g238 ( .A(n_222), .Y(n_238) );
BUFx3_ASAP7_75t_L g315 ( .A(n_222), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_225), .B(n_229), .C(n_238), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g245 ( .A1(n_225), .A2(n_238), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_225), .A2(n_238), .B(n_274), .C(n_275), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_225), .A2(n_238), .B(n_287), .C(n_288), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_225), .A2(n_238), .B(n_330), .C(n_331), .Y(n_329) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
BUFx3_ASAP7_75t_L g253 ( .A(n_227), .Y(n_253) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_230), .B(n_290), .Y(n_289) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g248 ( .A(n_231), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_234), .B(n_277), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_234), .A2(n_311), .B1(n_333), .B2(n_334), .Y(n_332) );
INVx4_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_241), .B(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_241), .A2(n_295), .B(n_302), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_241), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g349 ( .A(n_242), .Y(n_349) );
BUFx3_ASAP7_75t_L g357 ( .A(n_242), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_242), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g368 ( .A(n_242), .B(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_242), .B(n_256), .Y(n_397) );
AND2x2_ASAP7_75t_L g466 ( .A(n_242), .B(n_400), .Y(n_466) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_254), .Y(n_242) );
INVx1_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
INVx2_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_243), .A2(n_261), .B(n_307), .C(n_308), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx5_ASAP7_75t_L g311 ( .A(n_251), .Y(n_311) );
INVx2_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
INVx2_ASAP7_75t_SL g360 ( .A(n_255), .Y(n_360) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_271), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_256), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g402 ( .A(n_256), .Y(n_402) );
AND2x2_ASAP7_75t_L g413 ( .A(n_256), .B(n_369), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_256), .B(n_398), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_256), .B(n_400), .Y(n_445) );
AND2x2_ASAP7_75t_L g504 ( .A(n_256), .B(n_449), .Y(n_504) );
INVx4_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g374 ( .A(n_257), .B(n_271), .Y(n_374) );
AND2x2_ASAP7_75t_L g384 ( .A(n_257), .B(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g406 ( .A(n_257), .Y(n_406) );
AND3x2_ASAP7_75t_L g465 ( .A(n_257), .B(n_466), .C(n_467), .Y(n_465) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_269), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_262), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_261), .A2(n_296), .B(n_297), .Y(n_295) );
O2A1O1Ixp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_267), .C(n_268), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_265), .A2(n_268), .B(n_299), .C(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
INVx1_ASAP7_75t_SL g400 ( .A(n_271), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_271), .B(n_349), .C(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_318), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_281), .A2(n_384), .B(n_436), .C(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_305), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_283), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g452 ( .A(n_283), .Y(n_452) );
AND2x2_ASAP7_75t_L g473 ( .A(n_283), .B(n_320), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_283), .B(n_382), .Y(n_501) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_294), .Y(n_283) );
AND2x2_ASAP7_75t_L g346 ( .A(n_284), .B(n_337), .Y(n_346) );
INVx2_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_320), .Y(n_373) );
AND2x2_ASAP7_75t_L g423 ( .A(n_284), .B(n_305), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_284), .Y(n_427) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_SL g337 ( .A(n_294), .Y(n_337) );
BUFx2_ASAP7_75t_L g363 ( .A(n_294), .Y(n_363) );
AND2x2_ASAP7_75t_L g490 ( .A(n_294), .B(n_305), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
INVx3_ASAP7_75t_SL g320 ( .A(n_305), .Y(n_320) );
AND2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g352 ( .A(n_305), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g382 ( .A(n_305), .B(n_342), .Y(n_382) );
OR2x2_ASAP7_75t_L g391 ( .A(n_305), .B(n_337), .Y(n_391) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_305), .Y(n_409) );
AND2x2_ASAP7_75t_L g414 ( .A(n_305), .B(n_367), .Y(n_414) );
AND2x2_ASAP7_75t_L g442 ( .A(n_305), .B(n_322), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_305), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g480 ( .A(n_305), .B(n_321), .Y(n_480) );
OR2x6_ASAP7_75t_L g305 ( .A(n_306), .B(n_316), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_312), .C(n_313), .Y(n_309) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_314), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g404 ( .A(n_320), .B(n_353), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_320), .B(n_346), .Y(n_432) );
AND2x2_ASAP7_75t_L g450 ( .A(n_320), .B(n_367), .Y(n_450) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_337), .Y(n_321) );
AND2x2_ASAP7_75t_L g351 ( .A(n_322), .B(n_337), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_322), .B(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
OR2x2_ASAP7_75t_L g437 ( .A(n_322), .B(n_357), .Y(n_437) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_327), .B(n_335), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_328), .Y(n_509) );
INVx1_ASAP7_75t_L g344 ( .A(n_335), .Y(n_344) );
AND2x2_ASAP7_75t_L g372 ( .A(n_337), .B(n_342), .Y(n_372) );
INVx1_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
AND2x2_ASAP7_75t_L g475 ( .A(n_337), .B(n_353), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_347), .B1(n_350), .B2(n_354), .C1(n_358), .C2(n_361), .Y(n_338) );
INVx1_ASAP7_75t_L g470 ( .A(n_339), .Y(n_470) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_345), .Y(n_339) );
AND2x2_ASAP7_75t_L g366 ( .A(n_340), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g377 ( .A(n_340), .B(n_346), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_340), .B(n_368), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_340), .A2(n_416), .B1(n_421), .B2(n_422), .C1(n_430), .C2(n_432), .Y(n_415) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g403 ( .A(n_342), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_342), .B(n_423), .Y(n_463) );
AND2x2_ASAP7_75t_L g474 ( .A(n_342), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_345), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_347), .B(n_398), .Y(n_461) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_349), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g419 ( .A(n_349), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx3_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_352), .A2(n_455), .B(n_458), .C(n_460), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_352), .B(n_389), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_352), .B(n_372), .Y(n_494) );
AND2x2_ASAP7_75t_L g367 ( .A(n_353), .B(n_363), .Y(n_367) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_357), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g446 ( .A(n_357), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g485 ( .A(n_357), .B(n_385), .Y(n_485) );
INVx1_ASAP7_75t_L g497 ( .A(n_357), .Y(n_497) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_360), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g478 ( .A(n_363), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_368), .B(n_370), .C(n_374), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_366), .A2(n_396), .B1(n_411), .B2(n_414), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_367), .B(n_381), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_367), .B(n_389), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_368), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g431 ( .A(n_368), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_368), .B(n_418), .Y(n_438) );
INVx2_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NOR4xp25_ASAP7_75t_L g376 ( .A(n_373), .B(n_377), .C(n_378), .D(n_381), .Y(n_376) );
INVx1_ASAP7_75t_SL g447 ( .A(n_374), .Y(n_447) );
AND2x2_ASAP7_75t_L g491 ( .A(n_374), .B(n_492), .Y(n_491) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_383), .B(n_386), .C(n_395), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_382), .B(n_452), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_384), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
INVx1_ASAP7_75t_SL g457 ( .A(n_385), .Y(n_457) );
AND2x2_ASAP7_75t_L g496 ( .A(n_385), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_389), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_393), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_394), .B(n_419), .Y(n_479) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_401), .B(n_403), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g499 ( .A(n_399), .Y(n_499) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_400), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_410), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_406), .Y(n_418) );
OR2x2_ASAP7_75t_L g456 ( .A(n_406), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI21xp33_ASAP7_75t_SL g451 ( .A1(n_409), .A2(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_413), .A2(n_440), .B1(n_443), .B2(n_450), .C(n_451), .Y(n_439) );
INVx1_ASAP7_75t_SL g483 ( .A(n_414), .Y(n_483) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OR2x2_ASAP7_75t_L g430 ( .A(n_418), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_427), .B2(n_428), .Y(n_422) );
INVx1_ASAP7_75t_L g462 ( .A(n_423), .Y(n_462) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_426), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NOR4xp25_ASAP7_75t_L g433 ( .A(n_434), .B(n_468), .C(n_481), .D(n_493), .Y(n_433) );
NAND3xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_439), .C(n_454), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_437), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_444), .B(n_449), .Y(n_453) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI221xp5_ASAP7_75t_SL g481 ( .A1(n_456), .A2(n_482), .B1(n_483), .B2(n_484), .C(n_486), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_458), .A2(n_473), .B(n_474), .C(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_459), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_476) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_471), .C(n_472), .Y(n_468) );
INVx1_ASAP7_75t_L g487 ( .A(n_480), .Y(n_487) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_488), .B(n_491), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI221xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_495), .B1(n_498), .B2(n_500), .C(n_502), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
OAI322xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .A3(n_516), .B1(n_518), .B2(n_520), .C1(n_521), .C2(n_523), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
endmodule