module fake_jpeg_28443_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_40),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_28),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_64),
.B1(n_68),
.B2(n_22),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_35),
.B(n_33),
.C(n_25),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_36),
.B1(n_44),
.B2(n_20),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_41),
.B1(n_24),
.B2(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_72),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_17),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_94),
.B1(n_70),
.B2(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_35),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_92),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_97),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_33),
.B(n_24),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_24),
.B(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_36),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_48),
.A2(n_23),
.B1(n_44),
.B2(n_32),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_36),
.Y(n_100)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_20),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_63),
.B1(n_57),
.B2(n_51),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_115),
.B1(n_84),
.B2(n_102),
.Y(n_137)
);

CKINVDCx10_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_99),
.B1(n_78),
.B2(n_92),
.C(n_13),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_44),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_80),
.C(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_84),
.B1(n_90),
.B2(n_76),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_5),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_114),
.CON(n_135),
.SN(n_135)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_153),
.B(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_119),
.B1(n_118),
.B2(n_120),
.Y(n_167)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_107),
.B(n_75),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_82),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_159),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_107),
.B(n_83),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_127),
.B1(n_119),
.B2(n_123),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_179),
.B1(n_159),
.B2(n_138),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_169),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_108),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_177),
.C(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_175),
.B1(n_176),
.B2(n_136),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_129),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_122),
.B1(n_112),
.B2(n_101),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_101),
.B1(n_102),
.B2(n_124),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_125),
.C(n_113),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_130),
.B1(n_6),
.B2(n_8),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_168),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_156),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_194),
.C(n_161),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_160),
.B(n_146),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_198),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_173),
.B1(n_163),
.B2(n_130),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_157),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_181),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_147),
.C(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_143),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_142),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_200),
.B1(n_179),
.B2(n_176),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_91),
.CI(n_155),
.CON(n_200),
.SN(n_200)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_200),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_172),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_187),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_167),
.B1(n_175),
.B2(n_170),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_194),
.B1(n_193),
.B2(n_198),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_171),
.B(n_164),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_189),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_214),
.B(n_195),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_223),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_219),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_184),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_208),
.C(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_206),
.C(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_230),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_209),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_236),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_211),
.B1(n_216),
.B2(n_217),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_237),
.B(n_232),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_228),
.B(n_231),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_233),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.A3(n_225),
.B1(n_173),
.B2(n_163),
.C1(n_14),
.C2(n_15),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_16),
.A3(n_82),
.B1(n_9),
.B2(n_5),
.C1(n_6),
.C2(n_20),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_242),
.C(n_16),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_6),
.B1(n_9),
.B2(n_20),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_9),
.Y(n_250)
);


endmodule