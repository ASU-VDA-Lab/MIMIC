module fake_jpeg_22872_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_10),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_35),
.B1(n_34),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_61),
.B1(n_31),
.B2(n_20),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_35),
.B1(n_36),
.B2(n_19),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_21),
.B1(n_26),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_74),
.B1(n_82),
.B2(n_83),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_69),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_33),
.B1(n_21),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_33),
.B1(n_26),
.B2(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_32),
.B1(n_18),
.B2(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_23),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_23),
.B1(n_36),
.B2(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_18),
.B1(n_37),
.B2(n_27),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_98),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_13),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_90),
.A2(n_120),
.B(n_6),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_64),
.B1(n_62),
.B2(n_56),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_29),
.C(n_24),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_53),
.Y(n_148)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_106),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_0),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_0),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_109),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_2),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_115),
.B1(n_103),
.B2(n_104),
.Y(n_135)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_6),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_75),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_125),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_132),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_112),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_105),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

AO21x2_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_68),
.B(n_65),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_135),
.B1(n_142),
.B2(n_154),
.Y(n_164)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_131),
.Y(n_169)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_85),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_77),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_69),
.B1(n_79),
.B2(n_58),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_86),
.B1(n_96),
.B2(n_9),
.Y(n_189)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_75),
.A3(n_60),
.B1(n_53),
.B2(n_9),
.Y(n_144)
);

XOR2x2_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_120),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_118),
.B(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_179),
.B(n_184),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_119),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_102),
.C(n_116),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_143),
.C(n_137),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_102),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_166),
.A2(n_178),
.B(n_96),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_120),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_170),
.B1(n_146),
.B2(n_126),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_121),
.B1(n_114),
.B2(n_101),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_99),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_102),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_180),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_109),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_100),
.B(n_95),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_116),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_127),
.A2(n_88),
.B(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_88),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_106),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_127),
.B1(n_135),
.B2(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_195),
.B1(n_203),
.B2(n_208),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_193),
.B(n_199),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_168),
.B1(n_167),
.B2(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_201),
.C(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_144),
.B1(n_123),
.B2(n_124),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_202),
.B(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_133),
.C(n_155),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_123),
.B(n_145),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_154),
.B1(n_130),
.B2(n_86),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_173),
.C(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_130),
.B1(n_86),
.B2(n_147),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_139),
.C(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_146),
.CI(n_126),
.CON(n_215),
.SN(n_215)
);

NOR4xp25_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_178),
.C(n_165),
.D(n_158),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_179),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_122),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_177),
.B(n_166),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_222),
.B(n_229),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_225),
.B(n_218),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_204),
.B1(n_200),
.B2(n_198),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_198),
.B1(n_204),
.B2(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_183),
.B1(n_160),
.B2(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_190),
.B1(n_200),
.B2(n_216),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_235),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_202),
.B(n_178),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_219),
.B(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_201),
.C(n_211),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_251),
.C(n_220),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_224),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_196),
.C(n_194),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_192),
.B1(n_215),
.B2(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_215),
.B1(n_172),
.B2(n_159),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_261),
.B1(n_234),
.B2(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_237),
.B(n_231),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_194),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_222),
.A2(n_172),
.B1(n_159),
.B2(n_163),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_255),
.B(n_253),
.C(n_261),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_266),
.B(n_276),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_226),
.B1(n_237),
.B2(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_259),
.B1(n_250),
.B2(n_246),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_220),
.C(n_241),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_228),
.C(n_219),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_238),
.C(n_242),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_274),
.C(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_225),
.C(n_227),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_243),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_244),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_259),
.B1(n_246),
.B2(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_264),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_282),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_252),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_270),
.C(n_268),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_290),
.Y(n_299)
);

AOI31xp33_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_262),
.A3(n_254),
.B(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_258),
.B(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_284),
.C(n_285),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_289),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_249),
.B(n_267),
.C(n_258),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_256),
.B1(n_249),
.B2(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_274),
.C(n_272),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_279),
.C(n_291),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.Y(n_311)
);

NOR2x1_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_295),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_287),
.B1(n_290),
.B2(n_269),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_247),
.B(n_260),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_297),
.A3(n_299),
.B1(n_294),
.B2(n_288),
.C1(n_296),
.C2(n_129),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_297),
.B(n_131),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_315),
.A3(n_140),
.B1(n_138),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_308),
.A3(n_312),
.B1(n_131),
.B2(n_129),
.C1(n_140),
.C2(n_138),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_7),
.C(n_8),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_15),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_11),
.Y(n_320)
);


endmodule