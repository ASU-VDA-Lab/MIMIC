module fake_ariane_1518_n_2756 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2756);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2756;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_762;
wire n_1468;
wire n_1661;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_2640;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_727;
wire n_699;
wire n_590;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1524;
wire n_1476;
wire n_2016;
wire n_1856;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_2676;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2372;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2105;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_272),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_52),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_186),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_478),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_582),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_566),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_94),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_470),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_304),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_130),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_296),
.Y(n_595)
);

BUFx2_ASAP7_75t_SL g596 ( 
.A(n_565),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_522),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_573),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_409),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_49),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_291),
.Y(n_601)
);

BUFx2_ASAP7_75t_SL g602 ( 
.A(n_285),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_374),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_257),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_295),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_451),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_407),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_266),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_580),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_251),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_577),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_395),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_429),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_295),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_175),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_13),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_237),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_282),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_263),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_116),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_327),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g623 ( 
.A(n_557),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_578),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_90),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_270),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_232),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_506),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_233),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_123),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_413),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_339),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_178),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_270),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_344),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_132),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_315),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_33),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_92),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_446),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_335),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_432),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_73),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_77),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_347),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_382),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_156),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_19),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_481),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_179),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_439),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_203),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_430),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_456),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_118),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_567),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_377),
.Y(n_660)
);

CKINVDCx16_ASAP7_75t_R g661 ( 
.A(n_570),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_571),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_426),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_371),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_430),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_575),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_561),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_81),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_296),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_8),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_345),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_289),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_356),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_347),
.Y(n_674)
);

INVx4_ASAP7_75t_R g675 ( 
.A(n_435),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_388),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_181),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_230),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_191),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_491),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_198),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_367),
.Y(n_682)
);

BUFx5_ASAP7_75t_L g683 ( 
.A(n_545),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_281),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_124),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_310),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_548),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_474),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_131),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_248),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_253),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_367),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_568),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_302),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_251),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_560),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_248),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_250),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_42),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_135),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_226),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_354),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_576),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_385),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_419),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_443),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_225),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_3),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_237),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_249),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_177),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_453),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_127),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_479),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_477),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_355),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_202),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_227),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_343),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_246),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_551),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_54),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_157),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_473),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_480),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_432),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_304),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_422),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_427),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_342),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_581),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_463),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_523),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_329),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_366),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_423),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_381),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_541),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_100),
.Y(n_740)
);

CKINVDCx6p67_ASAP7_75t_R g741 ( 
.A(n_443),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_466),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_95),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_7),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_56),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_253),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_455),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_118),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_153),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_59),
.Y(n_750)
);

CKINVDCx14_ASAP7_75t_R g751 ( 
.A(n_379),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_143),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_399),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_98),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_516),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_317),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_572),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_510),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_317),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_56),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_472),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_529),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_157),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_205),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_39),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_483),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_245),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_380),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_471),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_96),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_115),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_405),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_420),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_579),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_473),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_518),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_52),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_319),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_527),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_309),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_290),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_227),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_434),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_264),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_390),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_459),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_264),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_521),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_481),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_346),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_67),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_403),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_520),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_88),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_174),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_278),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_569),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_404),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_134),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_225),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_482),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_396),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_425),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_467),
.Y(n_804)
);

BUFx8_ASAP7_75t_SL g805 ( 
.A(n_204),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_482),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_380),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_390),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_147),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_475),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_397),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_379),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_204),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_421),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_438),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_110),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_195),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_414),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_267),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_286),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_423),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_94),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_348),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_574),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_505),
.Y(n_825)
);

CKINVDCx14_ASAP7_75t_R g826 ( 
.A(n_245),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_117),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_29),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_544),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_593),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_751),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_593),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_652),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_826),
.Y(n_834)
);

CKINVDCx14_ASAP7_75t_R g835 ( 
.A(n_637),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_652),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

CKINVDCx14_ASAP7_75t_R g838 ( 
.A(n_637),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_715),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_591),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_805),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_711),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_715),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_711),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_715),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_664),
.Y(n_846)
);

INVxp67_ASAP7_75t_SL g847 ( 
.A(n_711),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_715),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_805),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_715),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_715),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_711),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_712),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_712),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_623),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_755),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_712),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_587),
.Y(n_858)
);

INVxp33_ASAP7_75t_SL g859 ( 
.A(n_651),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_661),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_741),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_712),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_599),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_603),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_607),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_741),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_616),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_744),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_617),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_829),
.Y(n_870)
);

INVxp33_ASAP7_75t_SL g871 ( 
.A(n_654),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_619),
.Y(n_872)
);

CKINVDCx14_ASAP7_75t_R g873 ( 
.A(n_637),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_620),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_687),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_625),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_631),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_633),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_768),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_634),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_591),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_744),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_635),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_687),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_639),
.Y(n_885)
);

CKINVDCx16_ASAP7_75t_R g886 ( 
.A(n_787),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_643),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_656),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_744),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_632),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_657),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_722),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_669),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_722),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_674),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_676),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_678),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_681),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_682),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_686),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_697),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_698),
.Y(n_902)
);

INVxp33_ASAP7_75t_L g903 ( 
.A(n_668),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_702),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_722),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_704),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_709),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_744),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_773),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_773),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_710),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_824),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_773),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_727),
.Y(n_914)
);

BUFx5_ASAP7_75t_L g915 ( 
.A(n_644),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_776),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_728),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_730),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_666),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_738),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_760),
.Y(n_921)
);

INVxp33_ASAP7_75t_SL g922 ( 
.A(n_585),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_740),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_632),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_773),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_803),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_803),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_803),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_803),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_743),
.Y(n_930)
);

BUFx8_ASAP7_75t_SL g931 ( 
.A(n_840),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_916),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_916),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_842),
.B(n_667),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_919),
.B(n_673),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_837),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_919),
.B(n_930),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_839),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_916),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_916),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_841),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_916),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_843),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_845),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_882),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_841),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_848),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_850),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_851),
.A2(n_696),
.B(n_680),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_856),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_836),
.B(n_673),
.Y(n_951)
);

BUFx8_ASAP7_75t_L g952 ( 
.A(n_856),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_830),
.B(n_691),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_882),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_889),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_844),
.B(n_691),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_889),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_908),
.Y(n_958)
);

OA21x2_ASAP7_75t_L g959 ( 
.A1(n_852),
.A2(n_757),
.B(n_705),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_908),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_909),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_720),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_909),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_846),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_910),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_840),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_849),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_929),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_910),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_913),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_857),
.B(n_720),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_915),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_862),
.B(n_771),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_915),
.Y(n_975)
);

CKINVDCx6p67_ASAP7_75t_R g976 ( 
.A(n_831),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_915),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_879),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_852),
.A2(n_788),
.B(n_774),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_833),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_913),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_859),
.A2(n_685),
.B1(n_706),
.B2(n_655),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_834),
.B(n_797),
.Y(n_983)
);

BUFx8_ASAP7_75t_SL g984 ( 
.A(n_881),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_849),
.Y(n_985)
);

OAI22x1_ASAP7_75t_SL g986 ( 
.A1(n_881),
.A2(n_685),
.B1(n_706),
.B2(n_655),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_925),
.A2(n_662),
.B(n_793),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_925),
.Y(n_989)
);

OAI22x1_ASAP7_75t_SL g990 ( 
.A1(n_890),
.A2(n_767),
.B1(n_786),
.B2(n_723),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_928),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_928),
.A2(n_662),
.B(n_771),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_929),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_853),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_853),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_927),
.B(n_776),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_944),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_977),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_948),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_964),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_946),
.B(n_838),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_931),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_970),
.B(n_892),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_937),
.B(n_873),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_937),
.B(n_935),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_944),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_938),
.B(n_752),
.C(n_749),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_948),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_948),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_946),
.B(n_855),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_938),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_944),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_943),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_944),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_944),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_984),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_943),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_964),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_944),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_936),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_944),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_977),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_936),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_947),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_937),
.B(n_776),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_992),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_947),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_946),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_967),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_935),
.B(n_903),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_992),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_992),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_967),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_978),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_949),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_951),
.B(n_858),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_967),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_985),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_947),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_966),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_949),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_935),
.B(n_863),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_949),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_985),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_947),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_947),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_976),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_949),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_947),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_949),
.B(n_776),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_951),
.B(n_864),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_955),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_985),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_994),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_994),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_976),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_983),
.B(n_894),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_973),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_994),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_988),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_954),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_954),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_954),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_951),
.B(n_894),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_963),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_987),
.A2(n_868),
.B(n_854),
.Y(n_1068)
);

NAND2xp33_ASAP7_75t_L g1069 ( 
.A(n_973),
.B(n_855),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_955),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_988),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_963),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_965),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_970),
.B(n_834),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_987),
.A2(n_926),
.B(n_854),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_988),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_965),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_988),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_955),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_976),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_941),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_971),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_956),
.B(n_905),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_971),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_991),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_941),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_998),
.B(n_973),
.Y(n_1087)
);

INVxp33_ASAP7_75t_L g1088 ( 
.A(n_1031),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1012),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_999),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_999),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_998),
.B(n_975),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1041),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1012),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1014),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1066),
.A2(n_982),
.B1(n_870),
.B2(n_884),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1003),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1001),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1014),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1009),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1009),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1000),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1018),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_998),
.B(n_975),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1010),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1003),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1010),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1059),
.B(n_905),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1003),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1002),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_1021),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1018),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_1000),
.B(n_978),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1005),
.B(n_922),
.Y(n_1114)
);

AND2x6_ASAP7_75t_L g1115 ( 
.A(n_1036),
.B(n_1042),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_998),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1067),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1063),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1019),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1083),
.B(n_922),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_997),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1021),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1067),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1023),
.B(n_975),
.Y(n_1124)
);

CKINVDCx11_ASAP7_75t_R g1125 ( 
.A(n_1048),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1026),
.Y(n_1126)
);

CKINVDCx6p67_ASAP7_75t_R g1127 ( 
.A(n_1058),
.Y(n_1127)
);

XNOR2x2_ASAP7_75t_R g1128 ( 
.A(n_1011),
.B(n_982),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1063),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1072),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1023),
.B(n_1060),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1064),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1021),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1017),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1021),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_1031),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1072),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1073),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1006),
.B(n_912),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1037),
.A2(n_871),
.B1(n_859),
.B2(n_726),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1060),
.A2(n_737),
.B1(n_783),
.B2(n_871),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1064),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1080),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1019),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1073),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1065),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1035),
.B(n_886),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1077),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1077),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1082),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1006),
.B(n_912),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1037),
.B(n_860),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1074),
.B(n_870),
.C(n_860),
.Y(n_1153)
);

OAI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1081),
.A2(n_884),
.B1(n_875),
.B2(n_726),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1065),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1057),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1057),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1023),
.B(n_977),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1061),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1029),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1023),
.B(n_977),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_SL g1162 ( 
.A(n_1086),
.B(n_763),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1082),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1061),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1084),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1062),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1037),
.B(n_956),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1084),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1085),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1056),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1037),
.B(n_956),
.Y(n_1171)
);

AO22x2_ASAP7_75t_L g1172 ( 
.A1(n_1036),
.A2(n_990),
.B1(n_986),
.B2(n_602),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1004),
.B(n_952),
.Y(n_1173)
);

INVx8_ASAP7_75t_L g1174 ( 
.A(n_1071),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1056),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1030),
.Y(n_1176)
);

INVxp33_ASAP7_75t_L g1177 ( 
.A(n_1043),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1024),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1053),
.B(n_956),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_987),
.B(n_934),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1024),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_SL g1183 ( 
.A(n_1076),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1013),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1043),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1053),
.B(n_1060),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1025),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1078),
.Y(n_1188)
);

INVxp33_ASAP7_75t_L g1189 ( 
.A(n_1008),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1013),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1025),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1026),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1025),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1069),
.B(n_952),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_997),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1025),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1034),
.B(n_875),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_997),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1008),
.A2(n_723),
.B1(n_745),
.B2(n_733),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1028),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1015),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1038),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1028),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1028),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_997),
.B(n_1007),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1015),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1028),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1040),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1040),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1039),
.B(n_866),
.C(n_861),
.Y(n_1210)
);

XNOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1045),
.B(n_890),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1026),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1040),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1027),
.A2(n_934),
.B(n_959),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1040),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1050),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1026),
.B(n_956),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1016),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1055),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_997),
.B(n_915),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1050),
.Y(n_1221)
);

NAND2x1_ASAP7_75t_L g1222 ( 
.A(n_1026),
.B(n_996),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1044),
.A2(n_745),
.B1(n_763),
.B2(n_733),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_997),
.B(n_915),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1026),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1144),
.B(n_924),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1118),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1114),
.B(n_924),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1186),
.B(n_1044),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1089),
.B(n_1049),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1114),
.B(n_952),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1110),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1110),
.B(n_1134),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1113),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1120),
.A2(n_1050),
.B(n_1016),
.C(n_1046),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1136),
.B(n_952),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1109),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1118),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1099),
.Y(n_1240)
);

AND2x2_ASAP7_75t_SL g1241 ( 
.A(n_1223),
.B(n_986),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1136),
.B(n_952),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1102),
.B(n_950),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1109),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1109),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1113),
.B(n_921),
.Y(n_1247)
);

AO221x1_ASAP7_75t_L g1248 ( 
.A1(n_1154),
.A2(n_742),
.B1(n_950),
.B2(n_990),
.C(n_764),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_L g1249 ( 
.A(n_1116),
.B(n_1007),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1112),
.B(n_1049),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1117),
.B(n_1050),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1123),
.B(n_1020),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1130),
.B(n_1020),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1108),
.B(n_861),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1120),
.B(n_950),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_L g1256 ( 
.A(n_1134),
.B(n_866),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1137),
.Y(n_1257)
);

AND2x6_ASAP7_75t_L g1258 ( 
.A(n_1194),
.B(n_1027),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1113),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1119),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1179),
.B(n_950),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1138),
.Y(n_1262)
);

BUFx5_ASAP7_75t_L g1263 ( 
.A(n_1115),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1160),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_L g1265 ( 
.A(n_1116),
.B(n_1007),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1116),
.B(n_1007),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1088),
.B(n_767),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1171),
.B(n_962),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1171),
.B(n_962),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1145),
.Y(n_1270)
);

BUFx5_ASAP7_75t_L g1271 ( 
.A(n_1115),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1129),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1132),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1167),
.B(n_962),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1148),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1132),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1149),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1150),
.Y(n_1278)
);

NOR3xp33_ASAP7_75t_L g1279 ( 
.A(n_1153),
.B(n_1141),
.C(n_1139),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1088),
.B(n_1177),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1093),
.B(n_962),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1177),
.B(n_786),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1168),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1142),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1151),
.B(n_798),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1109),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1140),
.B(n_974),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1146),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1169),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1146),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1155),
.Y(n_1292)
);

OAI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1140),
.A2(n_648),
.B1(n_688),
.B2(n_615),
.C(n_601),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1116),
.B(n_1007),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1197),
.B(n_798),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1180),
.B(n_1022),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1155),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_L g1298 ( 
.A(n_1152),
.B(n_769),
.C(n_766),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1147),
.B(n_980),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1170),
.B(n_1047),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1182),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1170),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1225),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1173),
.B(n_1007),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1173),
.B(n_1054),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1175),
.B(n_1051),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1174),
.B(n_980),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1185),
.B(n_972),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1189),
.B(n_1054),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1189),
.B(n_1054),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1194),
.B(n_1160),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1174),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1219),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1156),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1156),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1157),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_SL g1317 ( 
.A(n_1166),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1157),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1175),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1178),
.B(n_972),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1096),
.B(n_800),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1219),
.B(n_800),
.Y(n_1322)
);

INVxp33_ASAP7_75t_L g1323 ( 
.A(n_1211),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1115),
.A2(n_1026),
.B1(n_972),
.B2(n_974),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1121),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1159),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1115),
.B(n_1022),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1159),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1178),
.B(n_972),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1164),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1174),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1164),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1090),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1115),
.A2(n_972),
.B1(n_974),
.B2(n_737),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1202),
.B(n_1054),
.Y(n_1335)
);

NOR3xp33_ASAP7_75t_L g1336 ( 
.A(n_1162),
.B(n_815),
.C(n_796),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1122),
.B(n_974),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1090),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1143),
.B(n_1054),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1133),
.B(n_980),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1143),
.B(n_1054),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1091),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1091),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1100),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_SL g1345 ( 
.A(n_1126),
.B(n_824),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1100),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1133),
.B(n_953),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1097),
.B(n_953),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1188),
.B(n_1070),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_SL g1350 ( 
.A(n_1166),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1225),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1097),
.B(n_953),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1106),
.B(n_1046),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1101),
.Y(n_1354)
);

NOR3xp33_ASAP7_75t_L g1355 ( 
.A(n_1162),
.B(n_816),
.C(n_770),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1106),
.B(n_1047),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1111),
.B(n_1051),
.Y(n_1357)
);

INVxp33_ASAP7_75t_SL g1358 ( 
.A(n_1098),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1111),
.B(n_1052),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1101),
.B(n_1052),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1176),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1105),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1105),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1107),
.B(n_1052),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1176),
.B(n_1183),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1107),
.B(n_915),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1191),
.B(n_915),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1135),
.B(n_1126),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1191),
.B(n_915),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1204),
.B(n_1032),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1204),
.B(n_1032),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1121),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1187),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1209),
.B(n_1033),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1209),
.B(n_1033),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1210),
.B(n_1223),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1184),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1192),
.B(n_865),
.Y(n_1378)
);

BUFx5_ASAP7_75t_L g1379 ( 
.A(n_1135),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1192),
.B(n_867),
.Y(n_1380)
);

INVxp33_ASAP7_75t_L g1381 ( 
.A(n_1125),
.Y(n_1381)
);

NAND2xp33_ASAP7_75t_L g1382 ( 
.A(n_1121),
.B(n_1070),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1193),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1127),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1215),
.B(n_1070),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1215),
.B(n_1070),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1221),
.B(n_1070),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1199),
.B(n_585),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1225),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1098),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1217),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1221),
.B(n_1070),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1196),
.B(n_604),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1200),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1203),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1207),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1208),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1184),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1213),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1212),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1125),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1212),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1121),
.B(n_1079),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1190),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1216),
.B(n_605),
.C(n_604),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1212),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1195),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_L g1408 ( 
.A(n_1195),
.B(n_1079),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1195),
.B(n_1079),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1190),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1201),
.B(n_1079),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1201),
.Y(n_1412)
);

NAND2xp33_ASAP7_75t_L g1413 ( 
.A(n_1195),
.B(n_1079),
.Y(n_1413)
);

BUFx5_ASAP7_75t_L g1414 ( 
.A(n_1198),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1172),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_SL g1416 ( 
.A(n_1128),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1206),
.B(n_1079),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1206),
.B(n_1068),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1198),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1212),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1218),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1218),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1181),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1198),
.B(n_605),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1241),
.A2(n_1172),
.B1(n_606),
.B2(n_595),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1231),
.B(n_1198),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1227),
.Y(n_1427)
);

OAI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1228),
.A2(n_612),
.B1(n_828),
.B2(n_610),
.C(n_608),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1240),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1245),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1257),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1307),
.B(n_1172),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1307),
.B(n_1205),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1321),
.B(n_1205),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1238),
.A2(n_1131),
.B1(n_1092),
.B2(n_1104),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1232),
.Y(n_1436)
);

AO22x2_ASAP7_75t_L g1437 ( 
.A1(n_1415),
.A2(n_777),
.B1(n_784),
.B2(n_782),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1239),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1307),
.B(n_869),
.Y(n_1439)
);

AO22x2_ASAP7_75t_L g1440 ( 
.A1(n_1288),
.A2(n_789),
.B1(n_801),
.B2(n_790),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1262),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1327),
.A2(n_1131),
.B(n_1158),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1270),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1255),
.B(n_1181),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1275),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1247),
.B(n_595),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1260),
.B(n_1087),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1277),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1272),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1295),
.A2(n_1092),
.B1(n_1104),
.B2(n_1087),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1278),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1226),
.B(n_1286),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1273),
.Y(n_1453)
);

AO22x2_ASAP7_75t_L g1454 ( 
.A1(n_1423),
.A2(n_818),
.B1(n_827),
.B2(n_823),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1284),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1234),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1290),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1355),
.A2(n_759),
.B1(n_874),
.B2(n_872),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_SL g1459 ( 
.A(n_1264),
.B(n_824),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1293),
.A2(n_1388),
.B1(n_1322),
.B2(n_1254),
.C(n_1376),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1301),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1276),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1282),
.A2(n_612),
.B1(n_828),
.B2(n_610),
.C(n_608),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1302),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1280),
.B(n_876),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1319),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1259),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1336),
.A2(n_878),
.B1(n_880),
.B2(n_877),
.Y(n_1468)
);

AO22x2_ASAP7_75t_L g1469 ( 
.A1(n_1261),
.A2(n_885),
.B1(n_887),
.B2(n_883),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1313),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1299),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1279),
.A2(n_893),
.B1(n_895),
.B2(n_891),
.C(n_888),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1243),
.A2(n_897),
.B1(n_898),
.B2(n_896),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1238),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1384),
.B(n_1222),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1283),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1283),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1317),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1312),
.B(n_899),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1281),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1328),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1330),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1331),
.B(n_1224),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1342),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1298),
.A2(n_901),
.B1(n_902),
.B2(n_900),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1233),
.B(n_1311),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1389),
.B(n_1220),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1285),
.Y(n_1488)
);

AND2x6_ASAP7_75t_SL g1489 ( 
.A(n_1365),
.B(n_904),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1267),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1361),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1317),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1343),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1344),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1358),
.B(n_1220),
.Y(n_1495)
);

AO22x2_ASAP7_75t_L g1496 ( 
.A1(n_1236),
.A2(n_907),
.B1(n_911),
.B2(n_906),
.Y(n_1496)
);

AO22x2_ASAP7_75t_L g1497 ( 
.A1(n_1242),
.A2(n_917),
.B1(n_918),
.B2(n_914),
.Y(n_1497)
);

AND2x6_ASAP7_75t_L g1498 ( 
.A(n_1389),
.B(n_991),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1373),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_L g1500 ( 
.A(n_1379),
.B(n_1124),
.Y(n_1500)
);

AND2x6_ASAP7_75t_L g1501 ( 
.A(n_1303),
.B(n_920),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1383),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1268),
.B(n_923),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1394),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1396),
.Y(n_1505)
);

OAI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1256),
.A2(n_592),
.B1(n_594),
.B2(n_588),
.C(n_586),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1269),
.B(n_600),
.Y(n_1507)
);

NAND2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1303),
.B(n_1351),
.Y(n_1508)
);

AO22x2_ASAP7_75t_L g1509 ( 
.A1(n_1248),
.A2(n_596),
.B1(n_1224),
.B2(n_675),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1289),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1391),
.B(n_1274),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1334),
.A2(n_613),
.B1(n_622),
.B2(n_618),
.C(n_614),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1291),
.Y(n_1514)
);

AO22x2_ASAP7_75t_L g1515 ( 
.A1(n_1377),
.A2(n_1124),
.B1(n_606),
.B2(n_595),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1399),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1292),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1390),
.A2(n_627),
.B1(n_629),
.B2(n_626),
.C(n_621),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1347),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1395),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1252),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1381),
.B(n_636),
.C(n_630),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1297),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1351),
.B(n_1401),
.Y(n_1524)
);

AO22x2_ASAP7_75t_L g1525 ( 
.A1(n_1398),
.A2(n_606),
.B1(n_958),
.B2(n_957),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1252),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1237),
.B(n_945),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1378),
.B(n_1158),
.Y(n_1528)
);

AO22x2_ASAP7_75t_L g1529 ( 
.A1(n_1404),
.A2(n_958),
.B1(n_961),
.B2(n_957),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_L g1530 ( 
.A(n_1237),
.B(n_945),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1416),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1314),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1308),
.B(n_638),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1253),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1378),
.B(n_640),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1380),
.B(n_641),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1253),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1315),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1296),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1393),
.A2(n_642),
.B1(n_649),
.B2(n_647),
.C(n_646),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1350),
.Y(n_1541)
);

AO22x2_ASAP7_75t_L g1542 ( 
.A1(n_1410),
.A2(n_958),
.B1(n_961),
.B2(n_957),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1380),
.B(n_1161),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1296),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1237),
.B(n_945),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1350),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1316),
.Y(n_1547)
);

AND2x6_ASAP7_75t_L g1548 ( 
.A(n_1324),
.B(n_945),
.Y(n_1548)
);

OAI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1405),
.A2(n_645),
.B1(n_660),
.B2(n_658),
.C(n_653),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1416),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1318),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1258),
.A2(n_1345),
.B1(n_1323),
.B2(n_1424),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1320),
.B(n_650),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1326),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1246),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1332),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1333),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1338),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_L g1559 ( 
.A(n_1339),
.B(n_1214),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1246),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1346),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1354),
.Y(n_1562)
);

BUFx8_ASAP7_75t_L g1563 ( 
.A(n_1246),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1412),
.A2(n_969),
.B1(n_981),
.B2(n_961),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1362),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1363),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1340),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1329),
.B(n_663),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1348),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1287),
.B(n_1161),
.Y(n_1570)
);

AO22x2_ASAP7_75t_L g1571 ( 
.A1(n_1421),
.A2(n_981),
.B1(n_993),
.B2(n_969),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_SL g1572 ( 
.A(n_1287),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1352),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1249),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1229),
.B(n_665),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1341),
.B(n_969),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1422),
.Y(n_1577)
);

AO22x2_ASAP7_75t_L g1578 ( 
.A1(n_1304),
.A2(n_1305),
.B1(n_1310),
.B2(n_1309),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1345),
.A2(n_677),
.B1(n_679),
.B2(n_672),
.C(n_671),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1251),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1349),
.B(n_1287),
.Y(n_1581)
);

AO22x2_ASAP7_75t_L g1582 ( 
.A1(n_1229),
.A2(n_993),
.B1(n_981),
.B2(n_927),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1335),
.Y(n_1583)
);

AO22x2_ASAP7_75t_L g1584 ( 
.A1(n_1230),
.A2(n_1250),
.B1(n_1418),
.B2(n_1306),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1230),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1250),
.Y(n_1586)
);

AO22x2_ASAP7_75t_L g1587 ( 
.A1(n_1418),
.A2(n_993),
.B1(n_926),
.B2(n_1068),
.Y(n_1587)
);

OR2x6_ASAP7_75t_SL g1588 ( 
.A(n_1337),
.B(n_670),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1300),
.Y(n_1589)
);

AO22x2_ASAP7_75t_L g1590 ( 
.A1(n_1306),
.A2(n_1068),
.B1(n_2),
.B2(n_0),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1258),
.B(n_684),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1370),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1370),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1235),
.A2(n_689),
.B1(n_694),
.B2(n_692),
.C(n_690),
.Y(n_1594)
);

AO22x2_ASAP7_75t_L g1595 ( 
.A1(n_1360),
.A2(n_1068),
.B1(n_2),
.B2(n_0),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1407),
.B(n_695),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1371),
.A2(n_700),
.B1(n_701),
.B2(n_699),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1411),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1265),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1411),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1374),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1375),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1407),
.B(n_707),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1375),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1419),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1258),
.B(n_708),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1258),
.B(n_713),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1367),
.A2(n_716),
.B(n_714),
.Y(n_1608)
);

AO22x2_ASAP7_75t_L g1609 ( 
.A1(n_1360),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_1609)
);

AO22x1_ASAP7_75t_L g1610 ( 
.A1(n_1244),
.A2(n_718),
.B1(n_719),
.B2(n_717),
.Y(n_1610)
);

NOR2xp67_ASAP7_75t_L g1611 ( 
.A(n_1400),
.B(n_609),
.Y(n_1611)
);

OAI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1367),
.A2(n_729),
.B1(n_731),
.B2(n_725),
.C(n_724),
.Y(n_1612)
);

AO22x2_ASAP7_75t_L g1613 ( 
.A1(n_1364),
.A2(n_1417),
.B1(n_1357),
.B2(n_1359),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1417),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1366),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1369),
.A2(n_746),
.B1(n_747),
.B2(n_736),
.C(n_735),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1364),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1385),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1419),
.B(n_721),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1385),
.A2(n_806),
.B(n_814),
.C(n_785),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1414),
.B(n_1325),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1325),
.B(n_955),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1386),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1325),
.B(n_955),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1386),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1528),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1460),
.B(n_1372),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1452),
.A2(n_1271),
.B1(n_1263),
.B2(n_1368),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1490),
.B(n_1372),
.Y(n_1629)
);

AOI21xp33_ASAP7_75t_L g1630 ( 
.A1(n_1434),
.A2(n_1369),
.B(n_1356),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1574),
.A2(n_1408),
.B(n_1382),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_SL g1632 ( 
.A(n_1531),
.B(n_1263),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1524),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1528),
.Y(n_1634)
);

AND2x6_ASAP7_75t_L g1635 ( 
.A(n_1543),
.B(n_1372),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1428),
.A2(n_1413),
.B(n_1387),
.C(n_1392),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1599),
.A2(n_1392),
.B(n_1387),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1426),
.A2(n_1409),
.B(n_1403),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1552),
.B(n_1379),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1474),
.A2(n_1353),
.B1(n_1294),
.B2(n_1266),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1480),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1500),
.A2(n_1271),
.B(n_1263),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1442),
.A2(n_1271),
.B(n_1263),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1476),
.A2(n_1406),
.B(n_1420),
.C(n_1402),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1585),
.A2(n_1271),
.B(n_1263),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1586),
.A2(n_1271),
.B(n_1414),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1477),
.B(n_1414),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1435),
.A2(n_1075),
.B(n_750),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1444),
.A2(n_1414),
.B(n_1379),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1584),
.A2(n_1414),
.B(n_1379),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1582),
.A2(n_1075),
.B(n_940),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1446),
.B(n_748),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1471),
.B(n_753),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1465),
.B(n_754),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1459),
.B(n_1379),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1433),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1439),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1511),
.B(n_756),
.Y(n_1658)
);

O2A1O1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1463),
.A2(n_940),
.B(n_933),
.C(n_765),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1575),
.A2(n_1075),
.B(n_772),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1470),
.B(n_1075),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1495),
.B(n_761),
.Y(n_1662)
);

AO21x1_ASAP7_75t_L g1663 ( 
.A1(n_1591),
.A2(n_1607),
.B(n_1606),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1584),
.A2(n_1593),
.B(n_1592),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_SL g1665 ( 
.A(n_1436),
.B(n_775),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1563),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1543),
.B(n_609),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1555),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1501),
.A2(n_778),
.B1(n_781),
.B2(n_780),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1567),
.B(n_791),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1450),
.A2(n_794),
.B(n_792),
.Y(n_1671)
);

INVx5_ASAP7_75t_L g1672 ( 
.A(n_1498),
.Y(n_1672)
);

AO21x1_ASAP7_75t_L g1673 ( 
.A1(n_1521),
.A2(n_940),
.B(n_933),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1519),
.B(n_1569),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1508),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1540),
.A2(n_933),
.B(n_799),
.C(n_802),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1573),
.B(n_1526),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1534),
.B(n_795),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1478),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1601),
.A2(n_1604),
.B(n_1602),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1550),
.B(n_804),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1537),
.B(n_807),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1588),
.B(n_808),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1456),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1539),
.B(n_809),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1467),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1580),
.A2(n_979),
.B(n_959),
.Y(n_1687)
);

AOI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1582),
.A2(n_979),
.B(n_960),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1544),
.A2(n_825),
.B(n_611),
.Y(n_1689)
);

AOI22x1_ASAP7_75t_L g1690 ( 
.A1(n_1609),
.A2(n_810),
.B1(n_812),
.B2(n_811),
.Y(n_1690)
);

BUFx4f_ASAP7_75t_L g1691 ( 
.A(n_1501),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1440),
.B(n_813),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1440),
.B(n_817),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1520),
.B(n_819),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1615),
.A2(n_590),
.B(n_589),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1622),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1559),
.A2(n_598),
.B(n_597),
.Y(n_1697)
);

AOI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1587),
.A2(n_960),
.B(n_955),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1621),
.A2(n_628),
.B(n_624),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1579),
.B(n_821),
.C(n_820),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1458),
.B(n_822),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1427),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1429),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1430),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1622),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1518),
.B(n_659),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1572),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1625),
.A2(n_703),
.B(n_693),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1512),
.A2(n_995),
.B(n_732),
.C(n_739),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1613),
.A2(n_758),
.B(n_734),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1613),
.A2(n_779),
.B(n_762),
.Y(n_1711)
);

AOI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1587),
.A2(n_1578),
.B(n_1469),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1608),
.A2(n_995),
.B(n_960),
.C(n_968),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1431),
.B(n_1441),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1458),
.B(n_5),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1501),
.A2(n_996),
.B1(n_995),
.B2(n_683),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1491),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1618),
.A2(n_995),
.B(n_942),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1623),
.A2(n_995),
.B(n_942),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1438),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1589),
.A2(n_995),
.B(n_942),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1447),
.A2(n_942),
.B(n_932),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1596),
.A2(n_996),
.B(n_939),
.Y(n_1723)
);

AOI22x1_ASAP7_75t_L g1724 ( 
.A1(n_1609),
.A2(n_960),
.B1(n_968),
.B2(n_955),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1570),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1443),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1445),
.B(n_960),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1448),
.B(n_960),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1612),
.B(n_968),
.C(n_960),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1451),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1598),
.A2(n_942),
.B(n_932),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1489),
.B(n_6),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1475),
.B(n_968),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1455),
.B(n_1457),
.Y(n_1735)
);

AO21x1_ASAP7_75t_L g1736 ( 
.A1(n_1487),
.A2(n_683),
.B(n_968),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1461),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1483),
.B(n_968),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1479),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1600),
.A2(n_942),
.B(n_932),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1614),
.A2(n_1486),
.B(n_1594),
.Y(n_1741)
);

AND2x6_ASAP7_75t_L g1742 ( 
.A(n_1464),
.B(n_942),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1503),
.B(n_6),
.Y(n_1743)
);

INVxp33_ASAP7_75t_SL g1744 ( 
.A(n_1546),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1475),
.B(n_932),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1578),
.A2(n_932),
.B(n_939),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1473),
.B(n_7),
.Y(n_1747)
);

BUFx8_ASAP7_75t_L g1748 ( 
.A(n_1603),
.Y(n_1748)
);

NOR2x1_ASAP7_75t_L g1749 ( 
.A(n_1522),
.B(n_932),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1616),
.A2(n_989),
.B(n_932),
.C(n_939),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1483),
.B(n_683),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1499),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1620),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1469),
.B(n_9),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1624),
.A2(n_939),
.B(n_989),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1502),
.B(n_10),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1504),
.B(n_11),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1624),
.A2(n_939),
.B(n_989),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1581),
.A2(n_939),
.B(n_989),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1505),
.B(n_12),
.Y(n_1760)
);

OAI321xp33_ASAP7_75t_L g1761 ( 
.A1(n_1425),
.A2(n_1506),
.A3(n_1549),
.B1(n_1432),
.B2(n_1472),
.C(n_1597),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1513),
.B(n_12),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1516),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_L g1764 ( 
.A(n_1610),
.B(n_13),
.C(n_14),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1581),
.A2(n_939),
.B(n_989),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_R g1766 ( 
.A(n_1492),
.B(n_485),
.Y(n_1766)
);

BUFx4f_ASAP7_75t_L g1767 ( 
.A(n_1498),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1507),
.B(n_14),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1498),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1553),
.B(n_15),
.Y(n_1770)
);

INVx11_ASAP7_75t_L g1771 ( 
.A(n_1548),
.Y(n_1771)
);

CKINVDCx6p67_ASAP7_75t_R g1772 ( 
.A(n_1432),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1449),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1468),
.B(n_1485),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1568),
.B(n_15),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1453),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1466),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1533),
.B(n_16),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1619),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1590),
.A2(n_989),
.B(n_488),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1590),
.A2(n_989),
.B(n_489),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1611),
.B(n_683),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1605),
.A2(n_490),
.B(n_486),
.Y(n_1783)
);

OAI321xp33_ASAP7_75t_L g1784 ( 
.A1(n_1583),
.A2(n_683),
.A3(n_19),
.B1(n_21),
.B2(n_17),
.C(n_18),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1576),
.A2(n_493),
.B(n_492),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1576),
.A2(n_495),
.B(n_494),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1595),
.A2(n_497),
.B(n_496),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1560),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1595),
.A2(n_499),
.B(n_498),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1548),
.A2(n_996),
.B(n_20),
.Y(n_1790)
);

AO32x1_ASAP7_75t_L g1791 ( 
.A1(n_1481),
.A2(n_22),
.A3(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1468),
.B(n_22),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1529),
.A2(n_501),
.B(n_500),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1541),
.B(n_23),
.C(n_24),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1462),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1529),
.A2(n_503),
.B(n_502),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1527),
.A2(n_996),
.B(n_24),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1482),
.B(n_25),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1530),
.A2(n_996),
.B(n_25),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1545),
.A2(n_996),
.B(n_26),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1485),
.B(n_26),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1542),
.A2(n_507),
.B(n_504),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1542),
.A2(n_509),
.B(n_508),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1454),
.B(n_1437),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1454),
.B(n_27),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1484),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1493),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1807)
);

AOI22x1_ASAP7_75t_L g1808 ( 
.A1(n_1617),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1437),
.B(n_1494),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1515),
.B(n_30),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1515),
.B(n_31),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1547),
.B(n_32),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1714),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1674),
.B(n_1551),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1677),
.B(n_1554),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1702),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1641),
.B(n_1556),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1672),
.B(n_1557),
.Y(n_1818)
);

NOR3xp33_ASAP7_75t_SL g1819 ( 
.A(n_1794),
.B(n_1617),
.C(n_1561),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1662),
.A2(n_1768),
.B(n_1671),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1735),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1733),
.B(n_1558),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1809),
.B(n_1562),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1764),
.A2(n_1566),
.B(n_1577),
.C(n_1565),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1631),
.A2(n_1571),
.B(n_1564),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1696),
.B(n_1705),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1744),
.B(n_32),
.Y(n_1827)
);

BUFx12f_ASAP7_75t_L g1828 ( 
.A(n_1666),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1761),
.A2(n_1510),
.B(n_1514),
.C(n_1488),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1703),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1648),
.A2(n_1571),
.B(n_1564),
.Y(n_1831)
);

A2O1A1Ixp33_ASAP7_75t_SL g1832 ( 
.A1(n_1665),
.A2(n_1517),
.B(n_1532),
.C(n_1523),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1715),
.B(n_1496),
.Y(n_1833)
);

AO22x1_ASAP7_75t_L g1834 ( 
.A1(n_1732),
.A2(n_1509),
.B1(n_1538),
.B2(n_1496),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1720),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1637),
.A2(n_1497),
.B(n_1525),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1672),
.B(n_1497),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1676),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1810),
.A2(n_37),
.B(n_34),
.C(n_36),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1629),
.B(n_36),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1773),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1776),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1739),
.B(n_37),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1811),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_R g1845 ( 
.A(n_1707),
.B(n_511),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1686),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1795),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1804),
.B(n_38),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1704),
.Y(n_1849)
);

OAI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1790),
.A2(n_42),
.B(n_41),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1706),
.A2(n_996),
.B(n_40),
.Y(n_1851)
);

AND2x6_ASAP7_75t_L g1852 ( 
.A(n_1769),
.B(n_683),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1707),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1778),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1726),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1657),
.B(n_43),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1788),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1801),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.C(n_47),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1642),
.A2(n_45),
.B(n_46),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1684),
.B(n_47),
.Y(n_1860)
);

OA22x2_ASAP7_75t_L g1861 ( 
.A1(n_1774),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1730),
.Y(n_1862)
);

INVx5_ASAP7_75t_L g1863 ( 
.A(n_1672),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1737),
.B(n_48),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1696),
.B(n_50),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1767),
.B(n_51),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1649),
.A2(n_51),
.B(n_53),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1679),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1633),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1752),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1652),
.B(n_53),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1748),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1767),
.B(n_54),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1763),
.B(n_55),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1805),
.A2(n_996),
.B1(n_58),
.B2(n_55),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1680),
.B(n_57),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1729),
.A2(n_57),
.B(n_58),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1650),
.A2(n_59),
.B(n_60),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1627),
.B(n_60),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1664),
.A2(n_61),
.B(n_62),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1770),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1683),
.B(n_1748),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1775),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1883)
);

NOR3xp33_ASAP7_75t_L g1884 ( 
.A(n_1784),
.B(n_64),
.C(n_65),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1633),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1633),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1792),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1709),
.A2(n_69),
.B(n_66),
.C(n_68),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1743),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1771),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1696),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1777),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1643),
.A2(n_72),
.B(n_73),
.Y(n_1893)
);

AO21x1_ASAP7_75t_L g1894 ( 
.A1(n_1787),
.A2(n_74),
.B(n_75),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1640),
.A2(n_74),
.B(n_75),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_R g1896 ( 
.A(n_1691),
.B(n_583),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1806),
.B(n_76),
.Y(n_1897)
);

A2O1A1Ixp33_ASAP7_75t_L g1898 ( 
.A1(n_1659),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1806),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_SL g1900 ( 
.A1(n_1808),
.A2(n_78),
.B(n_79),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1705),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1754),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1902)
);

NAND2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1691),
.B(n_512),
.Y(n_1903)
);

A2O1A1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1753),
.A2(n_83),
.B(n_80),
.C(n_82),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1762),
.B(n_82),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1725),
.B(n_83),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1690),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1626),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1741),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1705),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1812),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1756),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1727),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1807),
.B(n_87),
.C(n_88),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1757),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1717),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1760),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1646),
.A2(n_87),
.B(n_89),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_L g1919 ( 
.A(n_1779),
.B(n_89),
.C(n_90),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1728),
.Y(n_1920)
);

INVxp67_ASAP7_75t_SL g1921 ( 
.A(n_1647),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1681),
.B(n_91),
.Y(n_1922)
);

A2O1A1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1710),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1923)
);

BUFx8_ASAP7_75t_L g1924 ( 
.A(n_1701),
.Y(n_1924)
);

INVxp33_ASAP7_75t_SL g1925 ( 
.A(n_1669),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1635),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1653),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1769),
.B(n_93),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1675),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1675),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1645),
.A2(n_95),
.B(n_96),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1747),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1932)
);

A2O1A1Ixp33_ASAP7_75t_SL g1933 ( 
.A1(n_1798),
.A2(n_100),
.B(n_97),
.C(n_99),
.Y(n_1933)
);

INVx5_ASAP7_75t_L g1934 ( 
.A(n_1635),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1658),
.B(n_101),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1626),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1654),
.A2(n_101),
.B(n_102),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1789),
.A2(n_1781),
.B(n_1780),
.C(n_1678),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1634),
.B(n_102),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1700),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1940)
);

O2A1O1Ixp5_ASAP7_75t_L g1941 ( 
.A1(n_1711),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1750),
.A2(n_106),
.B(n_107),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1636),
.A2(n_106),
.B(n_107),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1682),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1634),
.Y(n_1945)
);

NAND2x1p5_ASAP7_75t_L g1946 ( 
.A(n_1668),
.B(n_513),
.Y(n_1946)
);

A2O1A1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1689),
.A2(n_111),
.B(n_108),
.C(n_109),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1685),
.B(n_1656),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1670),
.B(n_111),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1656),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1712),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1656),
.B(n_112),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1692),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1713),
.A2(n_116),
.B(n_117),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1693),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1694),
.B(n_119),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1738),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1628),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1661),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1630),
.A2(n_122),
.B(n_123),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_L g1961 ( 
.A(n_1742),
.B(n_124),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1772),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1667),
.B(n_125),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1663),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1638),
.A2(n_125),
.B(n_126),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1639),
.B(n_126),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1660),
.A2(n_127),
.B(n_128),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1766),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1668),
.Y(n_1969)
);

OR2x6_ASAP7_75t_L g1970 ( 
.A(n_1793),
.B(n_514),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1635),
.Y(n_1971)
);

O2A1O1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1655),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1632),
.B(n_129),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1635),
.B(n_131),
.Y(n_1974)
);

OAI22x1_ASAP7_75t_L g1975 ( 
.A1(n_1724),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_1975)
);

NOR3xp33_ASAP7_75t_L g1976 ( 
.A(n_1749),
.B(n_136),
.C(n_137),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1698),
.A2(n_517),
.B(n_515),
.Y(n_1977)
);

AO22x1_ASAP7_75t_L g1978 ( 
.A1(n_1742),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1734),
.Y(n_1979)
);

BUFx8_ASAP7_75t_L g1980 ( 
.A(n_1742),
.Y(n_1980)
);

AND2x2_ASAP7_75t_SL g1981 ( 
.A(n_1734),
.B(n_138),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1977),
.A2(n_1651),
.B(n_1796),
.Y(n_1982)
);

BUFx12f_ASAP7_75t_L g1983 ( 
.A(n_1968),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1961),
.A2(n_1820),
.B(n_1938),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1891),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_R g1986 ( 
.A(n_1845),
.B(n_1697),
.Y(n_1986)
);

OAI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1825),
.A2(n_1878),
.B(n_1836),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1831),
.A2(n_1803),
.B(n_1802),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1820),
.A2(n_1723),
.B(n_1719),
.Y(n_1989)
);

AO21x2_ASAP7_75t_L g1990 ( 
.A1(n_1964),
.A2(n_1673),
.B(n_1736),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1863),
.B(n_1745),
.Y(n_1991)
);

A2O1A1Ixp33_ASAP7_75t_L g1992 ( 
.A1(n_1949),
.A2(n_1783),
.B(n_1786),
.C(n_1785),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1819),
.B(n_1751),
.C(n_1708),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1868),
.Y(n_1994)
);

CKINVDCx11_ASAP7_75t_R g1995 ( 
.A(n_1828),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1942),
.A2(n_1688),
.B(n_1746),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1925),
.A2(n_1742),
.B1(n_1782),
.B2(n_1716),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1830),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1849),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1922),
.A2(n_1695),
.B(n_1799),
.C(n_1797),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1892),
.Y(n_2001)
);

INVx5_ASAP7_75t_L g2002 ( 
.A(n_1863),
.Y(n_2002)
);

OR2x6_ASAP7_75t_L g2003 ( 
.A(n_1903),
.B(n_1644),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1863),
.B(n_1759),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1970),
.A2(n_1718),
.B(n_1791),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1855),
.Y(n_2006)
);

O2A1O1Ixp5_ASAP7_75t_L g2007 ( 
.A1(n_1943),
.A2(n_1800),
.B(n_1722),
.C(n_1699),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_L g2008 ( 
.A1(n_1893),
.A2(n_1867),
.B(n_1931),
.Y(n_2008)
);

AOI221x1_ASAP7_75t_L g2009 ( 
.A1(n_1880),
.A2(n_1740),
.B1(n_1731),
.B2(n_1721),
.C(n_1687),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1846),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1816),
.Y(n_2011)
);

NOR2x1_ASAP7_75t_SL g2012 ( 
.A(n_1934),
.B(n_1791),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1835),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1970),
.A2(n_1758),
.B(n_1755),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1895),
.A2(n_1765),
.B(n_139),
.Y(n_2015)
);

AOI221x1_ASAP7_75t_L g2016 ( 
.A1(n_1880),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1970),
.A2(n_140),
.B(n_141),
.Y(n_2017)
);

AND3x4_ASAP7_75t_L g2018 ( 
.A(n_1916),
.B(n_1884),
.C(n_1929),
.Y(n_2018)
);

BUFx12f_ASAP7_75t_L g2019 ( 
.A(n_1872),
.Y(n_2019)
);

AO21x2_ASAP7_75t_L g2020 ( 
.A1(n_1837),
.A2(n_524),
.B(n_519),
.Y(n_2020)
);

OAI22x1_ASAP7_75t_L g2021 ( 
.A1(n_1833),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_2021)
);

AO31x2_ASAP7_75t_L g2022 ( 
.A1(n_1951),
.A2(n_526),
.A3(n_528),
.B(n_525),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1953),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1954),
.A2(n_146),
.B(n_147),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1953),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1932),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_2026)
);

OAI22x1_ASAP7_75t_L g2027 ( 
.A1(n_1813),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1821),
.B(n_152),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1862),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1870),
.Y(n_2030)
);

BUFx12f_ASAP7_75t_L g2031 ( 
.A(n_1924),
.Y(n_2031)
);

AND2x6_ASAP7_75t_L g2032 ( 
.A(n_1971),
.B(n_530),
.Y(n_2032)
);

AO22x2_ASAP7_75t_L g2033 ( 
.A1(n_1823),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1850),
.A2(n_154),
.B(n_155),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1934),
.B(n_531),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_SL g2036 ( 
.A(n_1962),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1877),
.A2(n_158),
.B(n_159),
.Y(n_2037)
);

OAI22x1_ASAP7_75t_L g2038 ( 
.A1(n_1912),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_2038)
);

CKINVDCx11_ASAP7_75t_R g2039 ( 
.A(n_1857),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1857),
.B(n_160),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_SL g2041 ( 
.A1(n_1909),
.A2(n_161),
.B(n_162),
.Y(n_2041)
);

OAI21x1_ASAP7_75t_L g2042 ( 
.A1(n_1918),
.A2(n_533),
.B(n_532),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1850),
.A2(n_1967),
.B(n_1919),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_1839),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1981),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1817),
.B(n_165),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1899),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1840),
.B(n_1979),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1921),
.A2(n_166),
.B(n_167),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_SL g2050 ( 
.A1(n_1904),
.A2(n_166),
.B(n_167),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1975),
.A2(n_168),
.B(n_169),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1841),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1978),
.A2(n_168),
.B(n_169),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1859),
.A2(n_535),
.B(n_534),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1851),
.A2(n_170),
.B(n_171),
.Y(n_2055)
);

INVx5_ASAP7_75t_L g2056 ( 
.A(n_1852),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_1826),
.B(n_536),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1919),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1876),
.A2(n_1973),
.B(n_1965),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1842),
.Y(n_2060)
);

AOI221x1_ASAP7_75t_L g2061 ( 
.A1(n_1914),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.C(n_175),
.Y(n_2061)
);

AOI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1834),
.A2(n_173),
.B(n_176),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1847),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1915),
.B(n_176),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1917),
.B(n_177),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1888),
.A2(n_178),
.B(n_179),
.Y(n_2066)
);

AOI21xp33_ASAP7_75t_L g2067 ( 
.A1(n_1832),
.A2(n_180),
.B(n_181),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1818),
.A2(n_180),
.B(n_182),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1913),
.A2(n_538),
.B(n_537),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1894),
.A2(n_182),
.B(n_183),
.Y(n_2070)
);

A2O1A1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_1963),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1814),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1815),
.B(n_184),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1920),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1848),
.B(n_185),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1979),
.B(n_187),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_1980),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1891),
.Y(n_2078)
);

OAI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1941),
.A2(n_540),
.B(n_539),
.Y(n_2079)
);

AOI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_1844),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2080)
);

INVx1_ASAP7_75t_SL g2081 ( 
.A(n_1869),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1959),
.A2(n_188),
.B(n_189),
.Y(n_2082)
);

CKINVDCx6p67_ASAP7_75t_R g2083 ( 
.A(n_1885),
.Y(n_2083)
);

BUFx4_ASAP7_75t_SL g2084 ( 
.A(n_1905),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1937),
.A2(n_1879),
.B1(n_1838),
.B2(n_1875),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_1960),
.A2(n_190),
.B(n_191),
.Y(n_2086)
);

OAI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1898),
.A2(n_192),
.B(n_193),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1923),
.A2(n_192),
.B(n_193),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1871),
.B(n_194),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1926),
.B(n_542),
.Y(n_2090)
);

NOR4xp25_ASAP7_75t_L g2091 ( 
.A(n_1887),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_1824),
.A2(n_546),
.B(n_543),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1911),
.Y(n_2093)
);

O2A1O1Ixp5_ASAP7_75t_SL g2094 ( 
.A1(n_1928),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2094)
);

AOI21x1_ASAP7_75t_L g2095 ( 
.A1(n_1897),
.A2(n_197),
.B(n_199),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1958),
.A2(n_199),
.B(n_200),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1875),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2097)
);

AO21x1_ASAP7_75t_L g2098 ( 
.A1(n_1902),
.A2(n_201),
.B(n_203),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_1988),
.A2(n_1900),
.B(n_1936),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_2056),
.B(n_1908),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2056),
.B(n_1908),
.Y(n_2101)
);

OA21x2_ASAP7_75t_L g2102 ( 
.A1(n_1984),
.A2(n_1945),
.B(n_1974),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2011),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1998),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_L g2105 ( 
.A1(n_1982),
.A2(n_1957),
.B(n_1966),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2045),
.A2(n_1861),
.B1(n_1858),
.B2(n_1907),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2018),
.A2(n_2000),
.B1(n_2085),
.B2(n_2071),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_2010),
.Y(n_2108)
);

O2A1O1Ixp33_ASAP7_75t_L g2109 ( 
.A1(n_2023),
.A2(n_1933),
.B(n_1890),
.C(n_1881),
.Y(n_2109)
);

OAI21x1_ASAP7_75t_L g2110 ( 
.A1(n_1987),
.A2(n_1946),
.B(n_1972),
.Y(n_2110)
);

OAI21x1_ASAP7_75t_L g2111 ( 
.A1(n_1996),
.A2(n_1874),
.B(n_1864),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1999),
.B(n_1822),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2093),
.B(n_1927),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2006),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_L g2115 ( 
.A1(n_2014),
.A2(n_1829),
.B(n_1940),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2013),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1994),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1995),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1992),
.A2(n_1976),
.B(n_1947),
.Y(n_2119)
);

BUFx12f_ASAP7_75t_L g2120 ( 
.A(n_2031),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_1985),
.Y(n_2121)
);

OA21x2_ASAP7_75t_L g2122 ( 
.A1(n_2005),
.A2(n_1906),
.B(n_1952),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_2039),
.B(n_1969),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_2008),
.A2(n_1930),
.B(n_1955),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_1989),
.A2(n_1873),
.B(n_1866),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2029),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2043),
.A2(n_1980),
.B(n_1889),
.Y(n_2127)
);

AO21x2_ASAP7_75t_L g2128 ( 
.A1(n_2034),
.A2(n_1948),
.B(n_1843),
.Y(n_2128)
);

BUFx2_ASAP7_75t_L g2129 ( 
.A(n_2077),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_2009),
.A2(n_2092),
.B(n_2079),
.Y(n_2130)
);

OA21x2_ASAP7_75t_L g2131 ( 
.A1(n_2009),
.A2(n_1939),
.B(n_1901),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2030),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2047),
.Y(n_2133)
);

INVx3_ASAP7_75t_SL g2134 ( 
.A(n_2083),
.Y(n_2134)
);

AO21x2_ASAP7_75t_L g2135 ( 
.A1(n_1990),
.A2(n_1950),
.B(n_1883),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2004),
.A2(n_1854),
.B(n_1944),
.Y(n_2136)
);

BUFx8_ASAP7_75t_SL g2137 ( 
.A(n_2019),
.Y(n_2137)
);

CKINVDCx11_ASAP7_75t_R g2138 ( 
.A(n_1983),
.Y(n_2138)
);

OA21x2_ASAP7_75t_L g2139 ( 
.A1(n_2016),
.A2(n_1865),
.B(n_1856),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2084),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2033),
.A2(n_1924),
.B1(n_1935),
.B2(n_1956),
.Y(n_2141)
);

AO21x1_ASAP7_75t_L g2142 ( 
.A1(n_2025),
.A2(n_1860),
.B(n_1827),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_SL g2143 ( 
.A1(n_2012),
.A2(n_1853),
.B(n_1896),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2001),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2062),
.A2(n_1865),
.B(n_1882),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_2036),
.Y(n_2146)
);

AOI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2091),
.A2(n_1886),
.B1(n_1891),
.B2(n_1910),
.C(n_207),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_L g2148 ( 
.A1(n_2059),
.A2(n_1852),
.B(n_1910),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2072),
.B(n_1910),
.Y(n_2149)
);

OAI21x1_ASAP7_75t_L g2150 ( 
.A1(n_2017),
.A2(n_1852),
.B(n_549),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_1991),
.A2(n_1852),
.B(n_550),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_2016),
.A2(n_205),
.B(n_206),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_2048),
.Y(n_2153)
);

OAI21x1_ASAP7_75t_L g2154 ( 
.A1(n_2069),
.A2(n_552),
.B(n_547),
.Y(n_2154)
);

OAI21x1_ASAP7_75t_SL g2155 ( 
.A1(n_2098),
.A2(n_2087),
.B(n_2095),
.Y(n_2155)
);

OA21x2_ASAP7_75t_L g2156 ( 
.A1(n_2070),
.A2(n_206),
.B(n_207),
.Y(n_2156)
);

BUFx12f_ASAP7_75t_L g2157 ( 
.A(n_2075),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2056),
.B(n_208),
.Y(n_2158)
);

OAI21x1_ASAP7_75t_L g2159 ( 
.A1(n_2054),
.A2(n_554),
.B(n_553),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_L g2160 ( 
.A1(n_2042),
.A2(n_556),
.B(n_555),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2074),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2052),
.Y(n_2162)
);

CKINVDCx11_ASAP7_75t_R g2163 ( 
.A(n_2081),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2060),
.Y(n_2164)
);

NAND2x1p5_ASAP7_75t_L g2165 ( 
.A(n_2002),
.B(n_558),
.Y(n_2165)
);

NOR2xp67_ASAP7_75t_SL g2166 ( 
.A(n_2002),
.B(n_208),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2063),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2028),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2073),
.B(n_209),
.Y(n_2169)
);

OAI21x1_ASAP7_75t_L g2170 ( 
.A1(n_2007),
.A2(n_562),
.B(n_559),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_2015),
.A2(n_564),
.B(n_563),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2133),
.Y(n_2172)
);

NAND2x1p5_ASAP7_75t_L g2173 ( 
.A(n_2148),
.B(n_2002),
.Y(n_2173)
);

INVx4_ASAP7_75t_SL g2174 ( 
.A(n_2158),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_2108),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2104),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_2122),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2103),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2158),
.Y(n_2179)
);

BUFx2_ASAP7_75t_R g2180 ( 
.A(n_2137),
.Y(n_2180)
);

BUFx5_ASAP7_75t_L g2181 ( 
.A(n_2100),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2153),
.B(n_2100),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2107),
.A2(n_2033),
.B1(n_2055),
.B2(n_2066),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2142),
.A2(n_2097),
.B1(n_2058),
.B2(n_2044),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2103),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2114),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_2158),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2130),
.A2(n_2051),
.B(n_2053),
.Y(n_2188)
);

BUFx2_ASAP7_75t_R g2189 ( 
.A(n_2137),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2126),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_2163),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_2106),
.A2(n_1993),
.B1(n_2086),
.B2(n_2080),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2168),
.B(n_2046),
.Y(n_2193)
);

INVx2_ASAP7_75t_SL g2194 ( 
.A(n_2117),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_2102),
.Y(n_2195)
);

OAI21xp33_ASAP7_75t_L g2196 ( 
.A1(n_2119),
.A2(n_2050),
.B(n_2041),
.Y(n_2196)
);

AO21x2_ASAP7_75t_L g2197 ( 
.A1(n_2155),
.A2(n_2049),
.B(n_2037),
.Y(n_2197)
);

CKINVDCx11_ASAP7_75t_R g2198 ( 
.A(n_2120),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2117),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2141),
.A2(n_2026),
.B1(n_2003),
.B2(n_1997),
.Y(n_2200)
);

INVx5_ASAP7_75t_L g2201 ( 
.A(n_2120),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_2122),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2102),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_2102),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2132),
.B(n_2089),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2162),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2141),
.A2(n_2003),
.B1(n_2096),
.B2(n_2088),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_2148),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2122),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2164),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2116),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2167),
.Y(n_2212)
);

INVx5_ASAP7_75t_L g2213 ( 
.A(n_2100),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2116),
.Y(n_2214)
);

AOI21x1_ASAP7_75t_L g2215 ( 
.A1(n_2127),
.A2(n_2021),
.B(n_2038),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2196),
.A2(n_2128),
.B1(n_2156),
.B2(n_2139),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2195),
.Y(n_2217)
);

AOI21xp33_ASAP7_75t_L g2218 ( 
.A1(n_2197),
.A2(n_2183),
.B(n_2192),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2182),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2172),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2176),
.Y(n_2221)
);

OAI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2184),
.A2(n_2152),
.B(n_2125),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2182),
.B(n_2129),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_2198),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2186),
.Y(n_2225)
);

OAI22xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2202),
.A2(n_2113),
.B1(n_2112),
.B2(n_2118),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2195),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2190),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2195),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_SL g2230 ( 
.A(n_2180),
.B(n_2118),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2206),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2198),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2197),
.A2(n_2128),
.B1(n_2156),
.B2(n_2139),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2210),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2200),
.A2(n_2147),
.B1(n_2139),
.B2(n_2027),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2197),
.A2(n_2156),
.B1(n_2145),
.B2(n_2135),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2191),
.A2(n_2140),
.B1(n_2134),
.B2(n_2146),
.Y(n_2237)
);

AOI22xp33_ASAP7_75t_L g2238 ( 
.A1(n_2207),
.A2(n_2145),
.B1(n_2135),
.B2(n_2157),
.Y(n_2238)
);

OAI21xp33_ASAP7_75t_L g2239 ( 
.A1(n_2177),
.A2(n_2169),
.B(n_2109),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2203),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_2224),
.B(n_2174),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2220),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_2219),
.B(n_2174),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_2224),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2220),
.Y(n_2245)
);

OR2x6_ASAP7_75t_L g2246 ( 
.A(n_2224),
.B(n_2237),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2221),
.Y(n_2247)
);

NAND2xp33_ASAP7_75t_R g2248 ( 
.A(n_2232),
.B(n_2146),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_R g2249 ( 
.A(n_2230),
.B(n_2138),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_R g2250 ( 
.A(n_2223),
.B(n_2138),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_R g2251 ( 
.A(n_2223),
.B(n_2201),
.Y(n_2251)
);

INVx4_ASAP7_75t_SL g2252 ( 
.A(n_2246),
.Y(n_2252)
);

INVx4_ASAP7_75t_L g2253 ( 
.A(n_2246),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2244),
.B(n_2239),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2241),
.B(n_2219),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2243),
.B(n_2175),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2242),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2243),
.B(n_2175),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2249),
.Y(n_2259)
);

OR2x6_ASAP7_75t_SL g2260 ( 
.A(n_2252),
.B(n_2189),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2257),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2253),
.B(n_2255),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2254),
.B(n_2245),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2256),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2254),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2256),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2252),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2253),
.B(n_2239),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2252),
.B(n_2247),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2265),
.B(n_2261),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_2260),
.B(n_2259),
.Y(n_2271)
);

NAND3xp33_ASAP7_75t_L g2272 ( 
.A(n_2268),
.B(n_2267),
.C(n_2218),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2262),
.B(n_2253),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2263),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2264),
.B(n_2258),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2267),
.B(n_2222),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2266),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2263),
.B(n_2250),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2269),
.B(n_2221),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2269),
.B(n_2251),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2265),
.B(n_2225),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2281),
.Y(n_2282)
);

AND2x4_ASAP7_75t_SL g2283 ( 
.A(n_2273),
.B(n_2123),
.Y(n_2283)
);

INVx1_ASAP7_75t_SL g2284 ( 
.A(n_2271),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2280),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2274),
.B(n_2225),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_2276),
.B(n_2277),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2275),
.B(n_2134),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2270),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2270),
.B(n_2228),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2285),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2290),
.Y(n_2292)
);

NAND3xp33_ASAP7_75t_L g2293 ( 
.A(n_2289),
.B(n_2272),
.C(n_2278),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2282),
.B(n_2279),
.Y(n_2294)
);

CKINVDCx16_ASAP7_75t_R g2295 ( 
.A(n_2291),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2292),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2294),
.B(n_2284),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2293),
.B(n_2284),
.Y(n_2298)
);

OAI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2295),
.A2(n_2287),
.B1(n_2288),
.B2(n_2283),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2298),
.B(n_2286),
.Y(n_2300)
);

XOR2x2_ASAP7_75t_L g2301 ( 
.A(n_2298),
.B(n_2237),
.Y(n_2301)
);

OAI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2297),
.A2(n_2286),
.B(n_2279),
.Y(n_2302)
);

O2A1O1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2296),
.A2(n_2040),
.B(n_2065),
.C(n_2064),
.Y(n_2303)
);

AOI21xp33_ASAP7_75t_L g2304 ( 
.A1(n_2298),
.A2(n_1986),
.B(n_2236),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2301),
.Y(n_2305)
);

AOI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2300),
.A2(n_2235),
.B1(n_2248),
.B2(n_2157),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2302),
.B(n_2205),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2303),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_R g2309 ( 
.A(n_2299),
.B(n_2201),
.Y(n_2309)
);

OAI21xp33_ASAP7_75t_SL g2310 ( 
.A1(n_2304),
.A2(n_2235),
.B(n_2194),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2300),
.B(n_2228),
.Y(n_2311)
);

AOI21xp33_ASAP7_75t_SL g2312 ( 
.A1(n_2299),
.A2(n_2123),
.B(n_209),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2300),
.B(n_2205),
.Y(n_2313)
);

OAI322xp33_ASAP7_75t_SL g2314 ( 
.A1(n_2300),
.A2(n_2193),
.A3(n_2234),
.B1(n_2231),
.B2(n_2229),
.C1(n_2217),
.C2(n_2227),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2313),
.Y(n_2315)
);

INVxp67_ASAP7_75t_SL g2316 ( 
.A(n_2305),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2311),
.Y(n_2317)
);

AOI322xp5_ASAP7_75t_L g2318 ( 
.A1(n_2310),
.A2(n_2216),
.A3(n_2233),
.B1(n_2238),
.B2(n_2202),
.C1(n_2209),
.C2(n_2204),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2312),
.B(n_2201),
.Y(n_2319)
);

AOI322xp5_ASAP7_75t_L g2320 ( 
.A1(n_2308),
.A2(n_2203),
.A3(n_2204),
.B1(n_2201),
.B2(n_2229),
.C1(n_2217),
.C2(n_2227),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2307),
.Y(n_2321)
);

OAI221xp5_ASAP7_75t_SL g2322 ( 
.A1(n_2306),
.A2(n_2082),
.B1(n_2201),
.B2(n_2024),
.C(n_2217),
.Y(n_2322)
);

OAI22xp33_ASAP7_75t_SL g2323 ( 
.A1(n_2314),
.A2(n_2215),
.B1(n_2229),
.B2(n_2227),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2309),
.A2(n_2061),
.B(n_2226),
.Y(n_2324)
);

NOR2x1_ASAP7_75t_L g2325 ( 
.A(n_2305),
.B(n_2240),
.Y(n_2325)
);

OAI221xp5_ASAP7_75t_L g2326 ( 
.A1(n_2306),
.A2(n_2215),
.B1(n_2240),
.B2(n_2166),
.C(n_2068),
.Y(n_2326)
);

NOR2x1_ASAP7_75t_L g2327 ( 
.A(n_2305),
.B(n_2240),
.Y(n_2327)
);

NAND3xp33_ASAP7_75t_L g2328 ( 
.A(n_2316),
.B(n_2067),
.C(n_2163),
.Y(n_2328)
);

NOR3xp33_ASAP7_75t_SL g2329 ( 
.A(n_2315),
.B(n_210),
.C(n_211),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2319),
.B(n_2199),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2325),
.A2(n_2194),
.B1(n_2204),
.B2(n_2203),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2317),
.Y(n_2332)
);

AOI221xp5_ASAP7_75t_L g2333 ( 
.A1(n_2323),
.A2(n_2231),
.B1(n_2234),
.B2(n_2212),
.C(n_2076),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2327),
.A2(n_2170),
.B(n_2188),
.Y(n_2334)
);

NOR3xp33_ASAP7_75t_L g2335 ( 
.A(n_2321),
.B(n_2322),
.C(n_2326),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2324),
.Y(n_2336)
);

NOR3xp33_ASAP7_75t_L g2337 ( 
.A(n_2318),
.B(n_2035),
.C(n_2159),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2320),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2316),
.A2(n_2170),
.B(n_2188),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_SL g2340 ( 
.A(n_2317),
.B(n_2165),
.C(n_2094),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2316),
.B(n_210),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2316),
.B(n_211),
.Y(n_2342)
);

HB1xp67_ASAP7_75t_L g2343 ( 
.A(n_2332),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2341),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2330),
.B(n_2182),
.Y(n_2345)
);

XOR2x2_ASAP7_75t_L g2346 ( 
.A(n_2342),
.B(n_2165),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2338),
.B(n_2035),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_SL g2348 ( 
.A1(n_2336),
.A2(n_2090),
.B(n_212),
.Y(n_2348)
);

O2A1O1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2335),
.A2(n_2143),
.B(n_214),
.C(n_212),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2328),
.A2(n_213),
.B(n_214),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2340),
.A2(n_213),
.B(n_215),
.Y(n_2351)
);

NAND4xp25_ASAP7_75t_L g2352 ( 
.A(n_2333),
.B(n_2090),
.C(n_217),
.D(n_215),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2331),
.Y(n_2353)
);

AOI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2337),
.A2(n_2334),
.B1(n_2329),
.B2(n_2339),
.C(n_2208),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2338),
.A2(n_2187),
.B1(n_2179),
.B2(n_2208),
.Y(n_2355)
);

AOI322xp5_ASAP7_75t_L g2356 ( 
.A1(n_2336),
.A2(n_2057),
.A3(n_2187),
.B1(n_2179),
.B2(n_2208),
.C1(n_2101),
.C2(n_2213),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2343),
.A2(n_216),
.B(n_217),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2349),
.A2(n_2111),
.B(n_2171),
.Y(n_2358)
);

AOI322xp5_ASAP7_75t_L g2359 ( 
.A1(n_2344),
.A2(n_2347),
.A3(n_2353),
.B1(n_2354),
.B2(n_2345),
.C1(n_2350),
.C2(n_2348),
.Y(n_2359)
);

NAND4xp25_ASAP7_75t_SL g2360 ( 
.A(n_2351),
.B(n_219),
.C(n_216),
.D(n_218),
.Y(n_2360)
);

AOI221xp5_ASAP7_75t_L g2361 ( 
.A1(n_2355),
.A2(n_2057),
.B1(n_2208),
.B2(n_220),
.C(n_218),
.Y(n_2361)
);

AOI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2352),
.A2(n_2032),
.B1(n_2136),
.B2(n_2111),
.Y(n_2362)
);

AOI221xp5_ASAP7_75t_L g2363 ( 
.A1(n_2346),
.A2(n_2208),
.B1(n_221),
.B2(n_219),
.C(n_220),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2356),
.A2(n_221),
.B(n_222),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2343),
.B(n_222),
.Y(n_2365)
);

OAI211xp5_ASAP7_75t_L g2366 ( 
.A1(n_2343),
.A2(n_226),
.B(n_223),
.C(n_224),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2343),
.B(n_2179),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2343),
.B(n_2174),
.Y(n_2368)
);

NOR3xp33_ASAP7_75t_L g2369 ( 
.A(n_2343),
.B(n_2160),
.C(n_2159),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2343),
.B(n_223),
.Y(n_2370)
);

OAI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2343),
.A2(n_2187),
.B1(n_2179),
.B2(n_2131),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_2343),
.B(n_2160),
.C(n_2154),
.Y(n_2372)
);

NOR2xp67_ASAP7_75t_L g2373 ( 
.A(n_2343),
.B(n_224),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2343),
.A2(n_2171),
.B(n_2136),
.Y(n_2374)
);

AOI221x1_ASAP7_75t_L g2375 ( 
.A1(n_2350),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2343),
.Y(n_2376)
);

A2O1A1Ixp33_ASAP7_75t_L g2377 ( 
.A1(n_2351),
.A2(n_2110),
.B(n_2154),
.C(n_2124),
.Y(n_2377)
);

NOR4xp25_ASAP7_75t_L g2378 ( 
.A(n_2344),
.B(n_231),
.C(n_228),
.D(n_229),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2373),
.Y(n_2379)
);

OAI211xp5_ASAP7_75t_SL g2380 ( 
.A1(n_2376),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2380)
);

NAND4xp25_ASAP7_75t_L g2381 ( 
.A(n_2359),
.B(n_2375),
.C(n_2370),
.D(n_2363),
.Y(n_2381)
);

NOR3xp33_ASAP7_75t_L g2382 ( 
.A(n_2365),
.B(n_234),
.C(n_235),
.Y(n_2382)
);

OAI211xp5_ASAP7_75t_L g2383 ( 
.A1(n_2366),
.A2(n_238),
.B(n_235),
.C(n_236),
.Y(n_2383)
);

NOR4xp25_ASAP7_75t_L g2384 ( 
.A(n_2360),
.B(n_239),
.C(n_236),
.D(n_238),
.Y(n_2384)
);

OAI21xp33_ASAP7_75t_L g2385 ( 
.A1(n_2368),
.A2(n_2187),
.B(n_2179),
.Y(n_2385)
);

NAND4xp25_ASAP7_75t_SL g2386 ( 
.A(n_2361),
.B(n_241),
.C(n_239),
.D(n_240),
.Y(n_2386)
);

OAI221xp5_ASAP7_75t_L g2387 ( 
.A1(n_2367),
.A2(n_2378),
.B1(n_2357),
.B2(n_2364),
.C(n_2362),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2358),
.Y(n_2388)
);

AOI322xp5_ASAP7_75t_L g2389 ( 
.A1(n_2377),
.A2(n_2187),
.A3(n_2101),
.B1(n_2213),
.B2(n_2144),
.C1(n_2078),
.C2(n_2022),
.Y(n_2389)
);

OAI211xp5_ASAP7_75t_SL g2390 ( 
.A1(n_2374),
.A2(n_2371),
.B(n_2369),
.C(n_2372),
.Y(n_2390)
);

AOI21xp33_ASAP7_75t_L g2391 ( 
.A1(n_2376),
.A2(n_240),
.B(n_241),
.Y(n_2391)
);

XNOR2xp5_ASAP7_75t_L g2392 ( 
.A(n_2373),
.B(n_242),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2373),
.A2(n_2032),
.B1(n_2020),
.B2(n_2131),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2373),
.Y(n_2394)
);

O2A1O1Ixp5_ASAP7_75t_SL g2395 ( 
.A1(n_2376),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_2395)
);

AOI222xp33_ASAP7_75t_L g2396 ( 
.A1(n_2376),
.A2(n_2032),
.B1(n_2174),
.B2(n_2115),
.C1(n_2150),
.C2(n_2110),
.Y(n_2396)
);

NOR3xp33_ASAP7_75t_L g2397 ( 
.A(n_2376),
.B(n_243),
.C(n_244),
.Y(n_2397)
);

OAI211xp5_ASAP7_75t_L g2398 ( 
.A1(n_2376),
.A2(n_249),
.B(n_246),
.C(n_247),
.Y(n_2398)
);

AOI211xp5_ASAP7_75t_L g2399 ( 
.A1(n_2376),
.A2(n_252),
.B(n_247),
.C(n_250),
.Y(n_2399)
);

O2A1O1Ixp33_ASAP7_75t_L g2400 ( 
.A1(n_2376),
.A2(n_255),
.B(n_252),
.C(n_254),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2376),
.B(n_254),
.Y(n_2401)
);

AOI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2376),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_2402)
);

INVx2_ASAP7_75t_SL g2403 ( 
.A(n_2368),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2378),
.B(n_256),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_R g2405 ( 
.A(n_2376),
.B(n_258),
.Y(n_2405)
);

NAND3xp33_ASAP7_75t_L g2406 ( 
.A(n_2373),
.B(n_259),
.C(n_260),
.Y(n_2406)
);

AOI322xp5_ASAP7_75t_L g2407 ( 
.A1(n_2376),
.A2(n_2101),
.A3(n_2213),
.B1(n_2022),
.B2(n_2161),
.C1(n_2121),
.C2(n_2178),
.Y(n_2407)
);

A2O1A1Ixp33_ASAP7_75t_L g2408 ( 
.A1(n_2376),
.A2(n_2124),
.B(n_2130),
.C(n_261),
.Y(n_2408)
);

AOI211xp5_ASAP7_75t_L g2409 ( 
.A1(n_2376),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_2409)
);

AOI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2376),
.A2(n_265),
.B1(n_262),
.B2(n_263),
.C(n_266),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2376),
.A2(n_262),
.B(n_265),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2373),
.A2(n_2032),
.B1(n_2131),
.B2(n_1985),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2376),
.B(n_267),
.Y(n_2413)
);

AOI221xp5_ASAP7_75t_L g2414 ( 
.A1(n_2376),
.A2(n_271),
.B1(n_268),
.B2(n_269),
.C(n_272),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2373),
.A2(n_1985),
.B1(n_2161),
.B2(n_2178),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2401),
.B(n_268),
.C(n_269),
.Y(n_2416)
);

NAND4xp75_ASAP7_75t_L g2417 ( 
.A(n_2404),
.B(n_274),
.C(n_271),
.D(n_273),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_SL g2418 ( 
.A(n_2405),
.B(n_2173),
.C(n_273),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2392),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2413),
.Y(n_2420)
);

NAND4xp75_ASAP7_75t_L g2421 ( 
.A(n_2403),
.B(n_276),
.C(n_274),
.D(n_275),
.Y(n_2421)
);

OAI222xp33_ASAP7_75t_L g2422 ( 
.A1(n_2387),
.A2(n_2173),
.B1(n_2213),
.B2(n_2121),
.C1(n_2149),
.C2(n_279),
.Y(n_2422)
);

NOR3xp33_ASAP7_75t_L g2423 ( 
.A(n_2379),
.B(n_275),
.C(n_276),
.Y(n_2423)
);

OAI21xp33_ASAP7_75t_L g2424 ( 
.A1(n_2381),
.A2(n_2151),
.B(n_2173),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2394),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2400),
.A2(n_2411),
.B(n_2398),
.Y(n_2426)
);

NOR3xp33_ASAP7_75t_L g2427 ( 
.A(n_2406),
.B(n_277),
.C(n_278),
.Y(n_2427)
);

NOR2x1_ASAP7_75t_L g2428 ( 
.A(n_2380),
.B(n_277),
.Y(n_2428)
);

INVx2_ASAP7_75t_SL g2429 ( 
.A(n_2388),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2386),
.B(n_279),
.Y(n_2430)
);

AOI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2390),
.A2(n_2382),
.B1(n_2383),
.B2(n_2397),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2399),
.Y(n_2432)
);

NAND3xp33_ASAP7_75t_L g2433 ( 
.A(n_2409),
.B(n_280),
.C(n_281),
.Y(n_2433)
);

NOR2x1_ASAP7_75t_L g2434 ( 
.A(n_2391),
.B(n_280),
.Y(n_2434)
);

NAND4xp75_ASAP7_75t_L g2435 ( 
.A(n_2402),
.B(n_284),
.C(n_282),
.D(n_283),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2384),
.B(n_283),
.Y(n_2436)
);

NOR3xp33_ASAP7_75t_L g2437 ( 
.A(n_2410),
.B(n_284),
.C(n_285),
.Y(n_2437)
);

NAND3xp33_ASAP7_75t_L g2438 ( 
.A(n_2395),
.B(n_286),
.C(n_287),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2414),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2408),
.Y(n_2440)
);

NOR3x1_ASAP7_75t_L g2441 ( 
.A(n_2385),
.B(n_287),
.C(n_288),
.Y(n_2441)
);

INVxp33_ASAP7_75t_L g2442 ( 
.A(n_2415),
.Y(n_2442)
);

NOR3xp33_ASAP7_75t_L g2443 ( 
.A(n_2389),
.B(n_2412),
.C(n_2393),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2396),
.A2(n_2407),
.B1(n_2181),
.B2(n_2115),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_L g2445 ( 
.A(n_2401),
.B(n_288),
.C(n_289),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2384),
.B(n_290),
.Y(n_2446)
);

NOR3xp33_ASAP7_75t_L g2447 ( 
.A(n_2379),
.B(n_291),
.C(n_292),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2392),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2401),
.B(n_292),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2392),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2401),
.B(n_293),
.Y(n_2451)
);

INVxp33_ASAP7_75t_SL g2452 ( 
.A(n_2405),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_SL g2453 ( 
.A1(n_2403),
.A2(n_2213),
.B1(n_2181),
.B2(n_2105),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2452),
.B(n_2022),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2436),
.Y(n_2455)
);

NOR2x1_ASAP7_75t_L g2456 ( 
.A(n_2421),
.B(n_293),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2429),
.B(n_2181),
.Y(n_2457)
);

AO21x1_ASAP7_75t_L g2458 ( 
.A1(n_2449),
.A2(n_2451),
.B(n_2432),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2420),
.B(n_294),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2417),
.Y(n_2460)
);

NOR3xp33_ASAP7_75t_SL g2461 ( 
.A(n_2446),
.B(n_294),
.C(n_297),
.Y(n_2461)
);

NOR2x1_ASAP7_75t_L g2462 ( 
.A(n_2416),
.B(n_297),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2428),
.Y(n_2463)
);

NAND4xp75_ASAP7_75t_L g2464 ( 
.A(n_2425),
.B(n_300),
.C(n_298),
.D(n_299),
.Y(n_2464)
);

NOR3xp33_ASAP7_75t_L g2465 ( 
.A(n_2419),
.B(n_298),
.C(n_299),
.Y(n_2465)
);

NOR2xp67_ASAP7_75t_L g2466 ( 
.A(n_2445),
.B(n_300),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2430),
.B(n_301),
.Y(n_2467)
);

NAND3x1_ASAP7_75t_L g2468 ( 
.A(n_2423),
.B(n_301),
.C(n_302),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2438),
.Y(n_2469)
);

NAND3xp33_ASAP7_75t_L g2470 ( 
.A(n_2447),
.B(n_303),
.C(n_305),
.Y(n_2470)
);

NOR3xp33_ASAP7_75t_L g2471 ( 
.A(n_2448),
.B(n_303),
.C(n_305),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2441),
.B(n_2450),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2434),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2426),
.B(n_306),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2431),
.B(n_306),
.C(n_307),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2427),
.B(n_307),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_SL g2477 ( 
.A(n_2418),
.B(n_308),
.C(n_309),
.Y(n_2477)
);

NOR2x1_ASAP7_75t_L g2478 ( 
.A(n_2435),
.B(n_308),
.Y(n_2478)
);

NOR2x1_ASAP7_75t_L g2479 ( 
.A(n_2433),
.B(n_310),
.Y(n_2479)
);

AND2x2_ASAP7_75t_SL g2480 ( 
.A(n_2437),
.B(n_311),
.Y(n_2480)
);

NOR4xp25_ASAP7_75t_L g2481 ( 
.A(n_2439),
.B(n_313),
.C(n_311),
.D(n_312),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2442),
.B(n_312),
.Y(n_2482)
);

NOR3x2_ASAP7_75t_L g2483 ( 
.A(n_2440),
.B(n_313),
.C(n_314),
.Y(n_2483)
);

XOR2x1_ASAP7_75t_L g2484 ( 
.A(n_2443),
.B(n_314),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2422),
.B(n_315),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2444),
.B(n_316),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2424),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2453),
.Y(n_2488)
);

AND3x4_ASAP7_75t_L g2489 ( 
.A(n_2430),
.B(n_316),
.C(n_318),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2452),
.B(n_318),
.Y(n_2490)
);

INVx2_ASAP7_75t_SL g2491 ( 
.A(n_2430),
.Y(n_2491)
);

INVx2_ASAP7_75t_SL g2492 ( 
.A(n_2430),
.Y(n_2492)
);

OAI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2416),
.A2(n_2099),
.B(n_319),
.Y(n_2493)
);

NOR2xp67_ASAP7_75t_SL g2494 ( 
.A(n_2429),
.B(n_320),
.Y(n_2494)
);

NAND4xp75_ASAP7_75t_L g2495 ( 
.A(n_2429),
.B(n_322),
.C(n_320),
.D(n_321),
.Y(n_2495)
);

NOR4xp75_ASAP7_75t_L g2496 ( 
.A(n_2429),
.B(n_323),
.C(n_321),
.D(n_322),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2429),
.B(n_323),
.C(n_324),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2452),
.B(n_324),
.Y(n_2498)
);

OAI22x1_ASAP7_75t_L g2499 ( 
.A1(n_2446),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2499)
);

AOI21xp33_ASAP7_75t_L g2500 ( 
.A1(n_2429),
.A2(n_325),
.B(n_326),
.Y(n_2500)
);

NOR3xp33_ASAP7_75t_L g2501 ( 
.A(n_2425),
.B(n_328),
.C(n_329),
.Y(n_2501)
);

NOR2xp67_ASAP7_75t_L g2502 ( 
.A(n_2416),
.B(n_328),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2417),
.Y(n_2503)
);

NAND2x1p5_ASAP7_75t_L g2504 ( 
.A(n_2429),
.B(n_330),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2436),
.Y(n_2505)
);

NOR2x1_ASAP7_75t_L g2506 ( 
.A(n_2421),
.B(n_330),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2421),
.B(n_331),
.Y(n_2507)
);

NOR3xp33_ASAP7_75t_L g2508 ( 
.A(n_2425),
.B(n_331),
.C(n_332),
.Y(n_2508)
);

AOI22x1_ASAP7_75t_L g2509 ( 
.A1(n_2425),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2509)
);

NOR2x1_ASAP7_75t_L g2510 ( 
.A(n_2421),
.B(n_333),
.Y(n_2510)
);

NOR2xp67_ASAP7_75t_L g2511 ( 
.A(n_2416),
.B(n_334),
.Y(n_2511)
);

NOR2x1_ASAP7_75t_L g2512 ( 
.A(n_2421),
.B(n_335),
.Y(n_2512)
);

NAND3x1_ASAP7_75t_L g2513 ( 
.A(n_2423),
.B(n_336),
.C(n_337),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2436),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_2425),
.B(n_336),
.C(n_337),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2472),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2484),
.B(n_338),
.Y(n_2517)
);

NAND4xp75_ASAP7_75t_L g2518 ( 
.A(n_2458),
.B(n_340),
.C(n_338),
.D(n_339),
.Y(n_2518)
);

OAI31xp33_ASAP7_75t_L g2519 ( 
.A1(n_2504),
.A2(n_342),
.A3(n_340),
.B(n_341),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2489),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2491),
.B(n_341),
.Y(n_2521)
);

NAND5xp2_ASAP7_75t_L g2522 ( 
.A(n_2477),
.B(n_2461),
.C(n_2463),
.D(n_2469),
.E(n_2485),
.Y(n_2522)
);

AOI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2494),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.C(n_346),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2496),
.Y(n_2524)
);

AOI221xp5_ASAP7_75t_L g2525 ( 
.A1(n_2472),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.C(n_351),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2492),
.B(n_349),
.Y(n_2526)
);

NAND3xp33_ASAP7_75t_L g2527 ( 
.A(n_2473),
.B(n_350),
.C(n_352),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2483),
.Y(n_2528)
);

NOR2x1_ASAP7_75t_L g2529 ( 
.A(n_2474),
.B(n_352),
.Y(n_2529)
);

NOR3xp33_ASAP7_75t_L g2530 ( 
.A(n_2498),
.B(n_353),
.C(n_354),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2467),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2487),
.A2(n_2181),
.B1(n_2099),
.B2(n_356),
.Y(n_2532)
);

OAI311xp33_ASAP7_75t_L g2533 ( 
.A1(n_2455),
.A2(n_353),
.A3(n_355),
.B1(n_357),
.C1(n_358),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2505),
.B(n_357),
.Y(n_2534)
);

NOR2x1_ASAP7_75t_L g2535 ( 
.A(n_2459),
.B(n_358),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2514),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_2457),
.B(n_359),
.Y(n_2537)
);

NOR2xp67_ASAP7_75t_L g2538 ( 
.A(n_2497),
.B(n_2475),
.Y(n_2538)
);

NAND2x1p5_ASAP7_75t_L g2539 ( 
.A(n_2456),
.B(n_359),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_SL g2540 ( 
.A(n_2481),
.B(n_360),
.C(n_361),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2460),
.A2(n_2214),
.B1(n_2211),
.B2(n_2185),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2506),
.Y(n_2542)
);

NAND2x1p5_ASAP7_75t_L g2543 ( 
.A(n_2507),
.B(n_360),
.Y(n_2543)
);

AND3x4_ASAP7_75t_L g2544 ( 
.A(n_2510),
.B(n_2512),
.C(n_2478),
.Y(n_2544)
);

AND4x1_ASAP7_75t_L g2545 ( 
.A(n_2482),
.B(n_361),
.C(n_362),
.D(n_363),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2503),
.B(n_362),
.Y(n_2546)
);

NAND3xp33_ASAP7_75t_SL g2547 ( 
.A(n_2465),
.B(n_2471),
.C(n_2501),
.Y(n_2547)
);

NAND4xp75_ASAP7_75t_L g2548 ( 
.A(n_2462),
.B(n_363),
.C(n_364),
.D(n_365),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2468),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2513),
.Y(n_2550)
);

AOI221xp5_ASAP7_75t_L g2551 ( 
.A1(n_2499),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.C(n_368),
.Y(n_2551)
);

NOR3xp33_ASAP7_75t_L g2552 ( 
.A(n_2490),
.B(n_368),
.C(n_369),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2495),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2464),
.Y(n_2554)
);

AOI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2500),
.A2(n_2486),
.B(n_2488),
.Y(n_2555)
);

AND3x1_ASAP7_75t_L g2556 ( 
.A(n_2508),
.B(n_369),
.C(n_370),
.Y(n_2556)
);

AOI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2515),
.A2(n_2181),
.B1(n_371),
.B2(n_372),
.Y(n_2557)
);

INVxp67_ASAP7_75t_L g2558 ( 
.A(n_2479),
.Y(n_2558)
);

NOR2x1_ASAP7_75t_L g2559 ( 
.A(n_2470),
.B(n_370),
.Y(n_2559)
);

NOR2x1_ASAP7_75t_L g2560 ( 
.A(n_2466),
.B(n_2502),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2476),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2509),
.Y(n_2562)
);

NAND4xp25_ASAP7_75t_L g2563 ( 
.A(n_2511),
.B(n_372),
.C(n_373),
.D(n_374),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2476),
.A2(n_2181),
.B1(n_375),
.B2(n_376),
.Y(n_2564)
);

NOR2x1_ASAP7_75t_L g2565 ( 
.A(n_2493),
.B(n_2454),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2480),
.A2(n_373),
.B(n_375),
.Y(n_2566)
);

XNOR2x1_ASAP7_75t_L g2567 ( 
.A(n_2484),
.B(n_376),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2504),
.Y(n_2568)
);

XNOR2xp5_ASAP7_75t_L g2569 ( 
.A(n_2484),
.B(n_377),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2491),
.B(n_378),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2484),
.B(n_378),
.Y(n_2571)
);

NAND4xp75_ASAP7_75t_L g2572 ( 
.A(n_2458),
.B(n_381),
.C(n_382),
.D(n_383),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2491),
.B(n_383),
.Y(n_2573)
);

NAND4xp75_ASAP7_75t_L g2574 ( 
.A(n_2458),
.B(n_384),
.C(n_385),
.D(n_386),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2498),
.A2(n_384),
.B(n_386),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2491),
.B(n_387),
.Y(n_2576)
);

NOR3xp33_ASAP7_75t_L g2577 ( 
.A(n_2498),
.B(n_387),
.C(n_388),
.Y(n_2577)
);

NAND2x1p5_ASAP7_75t_L g2578 ( 
.A(n_2494),
.B(n_389),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2516),
.B(n_389),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_R g2580 ( 
.A(n_2536),
.B(n_2516),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_R g2581 ( 
.A(n_2516),
.B(n_391),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2567),
.B(n_391),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_R g2583 ( 
.A(n_2562),
.B(n_2547),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2569),
.B(n_2520),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_R g2585 ( 
.A(n_2553),
.B(n_2540),
.Y(n_2585)
);

NAND3xp33_ASAP7_75t_L g2586 ( 
.A(n_2517),
.B(n_392),
.C(n_393),
.Y(n_2586)
);

NAND2xp33_ASAP7_75t_SL g2587 ( 
.A(n_2526),
.B(n_392),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_R g2588 ( 
.A(n_2542),
.B(n_393),
.Y(n_2588)
);

XOR2xp5_ASAP7_75t_L g2589 ( 
.A(n_2560),
.B(n_394),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_R g2590 ( 
.A(n_2568),
.B(n_394),
.Y(n_2590)
);

NOR3xp33_ASAP7_75t_SL g2591 ( 
.A(n_2522),
.B(n_395),
.C(n_396),
.Y(n_2591)
);

XNOR2x1_ASAP7_75t_L g2592 ( 
.A(n_2544),
.B(n_397),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_R g2593 ( 
.A(n_2524),
.B(n_398),
.Y(n_2593)
);

NAND2xp33_ASAP7_75t_SL g2594 ( 
.A(n_2534),
.B(n_2521),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2556),
.B(n_398),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_R g2596 ( 
.A(n_2570),
.B(n_399),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2571),
.B(n_400),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_R g2598 ( 
.A(n_2576),
.B(n_400),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2561),
.B(n_401),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2549),
.B(n_2550),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2528),
.B(n_401),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_SL g2602 ( 
.A(n_2537),
.B(n_402),
.Y(n_2602)
);

XNOR2x1_ASAP7_75t_L g2603 ( 
.A(n_2529),
.B(n_2535),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_R g2604 ( 
.A(n_2554),
.B(n_402),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2519),
.B(n_403),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_R g2606 ( 
.A(n_2531),
.B(n_404),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_R g2607 ( 
.A(n_2558),
.B(n_405),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_R g2608 ( 
.A(n_2573),
.B(n_406),
.Y(n_2608)
);

NAND3xp33_ASAP7_75t_L g2609 ( 
.A(n_2555),
.B(n_406),
.C(n_407),
.Y(n_2609)
);

NAND2xp33_ASAP7_75t_SL g2610 ( 
.A(n_2537),
.B(n_408),
.Y(n_2610)
);

NAND2xp33_ASAP7_75t_SL g2611 ( 
.A(n_2546),
.B(n_408),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_R g2612 ( 
.A(n_2573),
.B(n_409),
.Y(n_2612)
);

NAND2xp33_ASAP7_75t_SL g2613 ( 
.A(n_2546),
.B(n_410),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2545),
.B(n_410),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2563),
.B(n_2578),
.Y(n_2615)
);

NAND3xp33_ASAP7_75t_L g2616 ( 
.A(n_2525),
.B(n_411),
.C(n_412),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_R g2617 ( 
.A(n_2533),
.B(n_411),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_R g2618 ( 
.A(n_2539),
.B(n_412),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_R g2619 ( 
.A(n_2543),
.B(n_413),
.Y(n_2619)
);

NAND3xp33_ASAP7_75t_L g2620 ( 
.A(n_2552),
.B(n_414),
.C(n_415),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_R g2621 ( 
.A(n_2518),
.B(n_415),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_R g2622 ( 
.A(n_2572),
.B(n_416),
.Y(n_2622)
);

NAND3xp33_ASAP7_75t_L g2623 ( 
.A(n_2530),
.B(n_416),
.C(n_417),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2523),
.B(n_417),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2538),
.B(n_418),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_SL g2626 ( 
.A(n_2574),
.B(n_418),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_SL g2627 ( 
.A(n_2566),
.B(n_419),
.C(n_420),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_R g2628 ( 
.A(n_2548),
.B(n_421),
.Y(n_2628)
);

XNOR2xp5_ASAP7_75t_L g2629 ( 
.A(n_2565),
.B(n_422),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2551),
.B(n_424),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2527),
.B(n_424),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_R g2632 ( 
.A(n_2577),
.B(n_425),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2603),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2589),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2629),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2592),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2595),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2617),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2614),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2600),
.A2(n_2557),
.B1(n_2564),
.B2(n_2559),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2580),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2625),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2602),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2584),
.A2(n_2532),
.B1(n_2575),
.B2(n_2541),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2610),
.Y(n_2645)
);

OAI211xp5_ASAP7_75t_L g2646 ( 
.A1(n_2583),
.A2(n_426),
.B(n_427),
.C(n_428),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2591),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2599),
.Y(n_2648)
);

INVx1_ASAP7_75t_SL g2649 ( 
.A(n_2618),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2611),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2613),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2608),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2612),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2582),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2619),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2597),
.A2(n_428),
.B1(n_429),
.B2(n_431),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2579),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2601),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2587),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2593),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2615),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2590),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2609),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2607),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2588),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2627),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2605),
.B(n_433),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2604),
.Y(n_2668)
);

INVx1_ASAP7_75t_SL g2669 ( 
.A(n_2581),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2606),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2586),
.Y(n_2671)
);

AO22x2_ASAP7_75t_L g2672 ( 
.A1(n_2623),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2626),
.Y(n_2673)
);

XNOR2xp5_ASAP7_75t_L g2674 ( 
.A(n_2638),
.B(n_2594),
.Y(n_2674)
);

AO22x2_ASAP7_75t_L g2675 ( 
.A1(n_2643),
.A2(n_2620),
.B1(n_2630),
.B2(n_2616),
.Y(n_2675)
);

XNOR2x1_ASAP7_75t_L g2676 ( 
.A(n_2633),
.B(n_2585),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2668),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2665),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2645),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2642),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2650),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2651),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2660),
.A2(n_2631),
.B1(n_2628),
.B2(n_2622),
.Y(n_2683)
);

INVxp67_ASAP7_75t_L g2684 ( 
.A(n_2659),
.Y(n_2684)
);

XNOR2xp5_ASAP7_75t_L g2685 ( 
.A(n_2649),
.B(n_2624),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2655),
.Y(n_2686)
);

XNOR2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2640),
.B(n_2596),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2652),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2653),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2672),
.Y(n_2690)
);

AOI22x1_ASAP7_75t_L g2691 ( 
.A1(n_2641),
.A2(n_2598),
.B1(n_2621),
.B2(n_2632),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2672),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2662),
.Y(n_2693)
);

XOR2xp5_ASAP7_75t_L g2694 ( 
.A(n_2634),
.B(n_436),
.Y(n_2694)
);

OAI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2647),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.C(n_440),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_SL g2696 ( 
.A1(n_2664),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2670),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2666),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2661),
.A2(n_441),
.B1(n_442),
.B2(n_444),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2656),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2667),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2674),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2676),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2680),
.B(n_2669),
.Y(n_2704)
);

AOI22x1_ASAP7_75t_L g2705 ( 
.A1(n_2677),
.A2(n_2673),
.B1(n_2636),
.B2(n_2639),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2687),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2678),
.B(n_2684),
.Y(n_2707)
);

OAI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2679),
.A2(n_2635),
.B1(n_2637),
.B2(n_2654),
.Y(n_2708)
);

HB1xp67_ASAP7_75t_L g2709 ( 
.A(n_2690),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2681),
.A2(n_2658),
.B(n_2648),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2691),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2692),
.B(n_2682),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2694),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2701),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2698),
.Y(n_2715)
);

OR2x2_ASAP7_75t_L g2716 ( 
.A(n_2686),
.B(n_2693),
.Y(n_2716)
);

OAI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2685),
.A2(n_2657),
.B(n_2671),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2675),
.Y(n_2718)
);

NOR3xp33_ASAP7_75t_L g2719 ( 
.A(n_2697),
.B(n_2646),
.C(n_2644),
.Y(n_2719)
);

AO21x2_ASAP7_75t_L g2720 ( 
.A1(n_2688),
.A2(n_2663),
.B(n_445),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2683),
.B(n_2181),
.Y(n_2721)
);

INVx2_ASAP7_75t_SL g2722 ( 
.A(n_2716),
.Y(n_2722)
);

AO22x2_ASAP7_75t_L g2723 ( 
.A1(n_2718),
.A2(n_2689),
.B1(n_2700),
.B2(n_2675),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2709),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2703),
.B(n_2696),
.Y(n_2725)
);

XNOR2xp5_ASAP7_75t_L g2726 ( 
.A(n_2705),
.B(n_2699),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2715),
.B(n_2695),
.Y(n_2727)
);

NAND4xp25_ASAP7_75t_L g2728 ( 
.A(n_2707),
.B(n_444),
.C(n_445),
.D(n_446),
.Y(n_2728)
);

OAI22x1_ASAP7_75t_L g2729 ( 
.A1(n_2702),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_2729)
);

OAI22xp5_ASAP7_75t_SL g2730 ( 
.A1(n_2706),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2712),
.Y(n_2731)
);

OAI221xp5_ASAP7_75t_L g2732 ( 
.A1(n_2717),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.C(n_453),
.Y(n_2732)
);

NAND3xp33_ASAP7_75t_L g2733 ( 
.A(n_2710),
.B(n_450),
.C(n_452),
.Y(n_2733)
);

AOI211xp5_ASAP7_75t_SL g2734 ( 
.A1(n_2724),
.A2(n_2708),
.B(n_2714),
.C(n_2704),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2731),
.Y(n_2735)
);

BUFx2_ASAP7_75t_L g2736 ( 
.A(n_2722),
.Y(n_2736)
);

OA22x2_ASAP7_75t_L g2737 ( 
.A1(n_2729),
.A2(n_2711),
.B1(n_2713),
.B2(n_2721),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2723),
.Y(n_2738)
);

BUFx2_ASAP7_75t_L g2739 ( 
.A(n_2723),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2725),
.Y(n_2740)
);

OAI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2733),
.A2(n_2719),
.B1(n_2720),
.B2(n_456),
.Y(n_2741)
);

NAND3x1_ASAP7_75t_L g2742 ( 
.A(n_2738),
.B(n_2727),
.C(n_2726),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2739),
.A2(n_2732),
.B1(n_2730),
.B2(n_2728),
.Y(n_2743)
);

AOI211xp5_ASAP7_75t_L g2744 ( 
.A1(n_2735),
.A2(n_454),
.B(n_455),
.C(n_457),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2736),
.Y(n_2745)
);

OAI22xp33_ASAP7_75t_L g2746 ( 
.A1(n_2734),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_2746)
);

OAI322xp33_ASAP7_75t_L g2747 ( 
.A1(n_2745),
.A2(n_2740),
.A3(n_2737),
.B1(n_2741),
.B2(n_2743),
.C1(n_2746),
.C2(n_2742),
.Y(n_2747)
);

AOI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2744),
.A2(n_458),
.B(n_460),
.Y(n_2748)
);

XNOR2xp5_ASAP7_75t_L g2749 ( 
.A(n_2742),
.B(n_460),
.Y(n_2749)
);

XOR2xp5_ASAP7_75t_L g2750 ( 
.A(n_2745),
.B(n_461),
.Y(n_2750)
);

AOI21xp33_ASAP7_75t_L g2751 ( 
.A1(n_2749),
.A2(n_461),
.B(n_462),
.Y(n_2751)
);

OR2x6_ASAP7_75t_L g2752 ( 
.A(n_2751),
.B(n_2747),
.Y(n_2752)
);

AOI22xp33_ASAP7_75t_L g2753 ( 
.A1(n_2752),
.A2(n_2748),
.B1(n_2750),
.B2(n_464),
.Y(n_2753)
);

AOI221xp5_ASAP7_75t_L g2754 ( 
.A1(n_2753),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.C(n_465),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2754),
.A2(n_465),
.B(n_466),
.Y(n_2755)
);

AOI211xp5_ASAP7_75t_L g2756 ( 
.A1(n_2755),
.A2(n_467),
.B(n_468),
.C(n_469),
.Y(n_2756)
);


endmodule