module real_jpeg_24568_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_0),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_0),
.B(n_17),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_0),
.B(n_37),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_0),
.B(n_32),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_0),
.Y(n_256)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_37),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_32),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_2),
.B(n_45),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_2),
.B(n_43),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_26),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_51),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_2),
.B(n_298),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_37),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_4),
.B(n_32),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_6),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_17),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_6),
.B(n_32),
.Y(n_310)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_8),
.B(n_45),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_8),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_43),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_8),
.B(n_26),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_51),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_9),
.B(n_32),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_45),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_43),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_26),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_51),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_9),
.B(n_73),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_11),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_11),
.B(n_37),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_45),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_43),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_11),
.B(n_26),
.Y(n_311)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_13),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_13),
.B(n_51),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_13),
.B(n_37),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_14),
.B(n_37),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_32),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_14),
.B(n_45),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_14),
.B(n_43),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_14),
.B(n_26),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_14),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_14),
.B(n_73),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_16),
.B(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_16),
.B(n_26),
.Y(n_115)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_17),
.Y(n_165)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_17),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_86),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_21),
.A2(n_22),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_62),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_23),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.C(n_47),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_24),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g85 ( 
.A(n_25),
.B(n_31),
.C(n_34),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_30),
.A2(n_31),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_31),
.B(n_78),
.C(n_81),
.Y(n_93)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_32),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_65),
.C(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_34),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_36),
.B(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_40),
.B(n_47),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_324),
.SN(n_324)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_47),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_361),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_53),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_58),
.C(n_61),
.Y(n_91)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_56),
.B(n_150),
.Y(n_242)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_56),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.C(n_74),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_64),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_65),
.A2(n_66),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_65),
.B(n_302),
.C(n_303),
.Y(n_323)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_67),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_68),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_70),
.B(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_334),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_74),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_74),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_74),
.B(n_330),
.C(n_333),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_75),
.B(n_86),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.C(n_85),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_76),
.A2(n_77),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_79),
.B(n_82),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_98),
.C(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_82),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_84),
.B(n_85),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_93),
.C(n_94),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_104),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_88),
.SN(n_88)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_98),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_362),
.C(n_363),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_350),
.C(n_351),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_338),
.C(n_339),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_314),
.C(n_315),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_282),
.C(n_283),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_248),
.C(n_249),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_218),
.C(n_219),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_196),
.C(n_197),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_178),
.C(n_179),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_156),
.C(n_157),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.C(n_147),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_139),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_140),
.C(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_137),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.C(n_152),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_162),
.C(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_177),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_182),
.C(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_195),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_212),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_213),
.C(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_208),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_207),
.C(n_208),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_201),
.Y(n_206)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_206),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_208),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.CI(n_211),
.CON(n_208),
.SN(n_208)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_210),
.C(n_211),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.CI(n_216),
.CON(n_213),
.SN(n_213)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_234),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_223),
.C(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_230),
.C(n_233),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_225),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.CI(n_228),
.CON(n_225),
.SN(n_225)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_241),
.C(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_240),
.B(n_273),
.C(n_274),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_269),
.B2(n_281),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_270),
.C(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_254),
.C(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_262),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_258),
.C(n_261),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_310),
.C(n_311),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_278),
.CI(n_280),
.CON(n_275),
.SN(n_275)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_312),
.B2(n_313),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_304),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_304),
.C(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_295),
.C(n_296),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_299),
.B1(n_300),
.B2(n_303),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.C(n_308),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_318),
.C(n_337),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_325),
.B2(n_337),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_323),
.C(n_324),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g368 ( 
.A(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_332),
.B2(n_336),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_349),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_343),
.C(n_349),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_346),
.C(n_347),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_354),
.C(n_359),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_358),
.B2(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_364),
.Y(n_365)
);


endmodule