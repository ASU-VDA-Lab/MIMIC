module fake_jpeg_3222_n_260 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_20),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_20),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_63),
.Y(n_84)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_65),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_39),
.Y(n_105)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_32),
.B1(n_40),
.B2(n_33),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_83),
.B1(n_59),
.B2(n_39),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_26),
.C(n_36),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_105),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_SL g80 ( 
.A(n_57),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_39),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_18),
.B1(n_35),
.B2(n_27),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_34),
.B1(n_35),
.B2(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_103),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_22),
.B1(n_21),
.B2(n_39),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_1),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_43),
.B(n_65),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_90),
.B(n_89),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_63),
.B1(n_98),
.B2(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_115),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_116),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_122),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_39),
.B(n_2),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_3),
.B(n_4),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_44),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_134),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_60),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_138),
.B1(n_95),
.B2(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx16f_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_2),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_102),
.C(n_88),
.Y(n_139)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_94),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_100),
.B1(n_71),
.B2(n_75),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_146),
.B1(n_153),
.B2(n_159),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_106),
.B1(n_107),
.B2(n_134),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_156),
.B(n_164),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_74),
.A3(n_87),
.B1(n_76),
.B2(n_95),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_100),
.B1(n_71),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_89),
.B1(n_94),
.B2(n_76),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_89),
.B1(n_94),
.B2(n_9),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_162),
.B1(n_124),
.B2(n_128),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_109),
.A2(n_122),
.B(n_127),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_125),
.C(n_117),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_133),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_174),
.C(n_179),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_126),
.B(n_119),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_159),
.B(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_184),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_6),
.A3(n_7),
.B1(n_10),
.B2(n_11),
.C1(n_135),
.C2(n_120),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_108),
.B(n_118),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_140),
.B1(n_153),
.B2(n_152),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_188),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_147),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_11),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_147),
.A3(n_172),
.B1(n_168),
.B2(n_167),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_171),
.B(n_180),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_139),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_146),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_145),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_145),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_151),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_184),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_161),
.B1(n_148),
.B2(n_152),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_205),
.B1(n_180),
.B2(n_172),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_209),
.C(n_220),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_166),
.C(n_171),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_222),
.B1(n_190),
.B2(n_196),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_207),
.B(n_195),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_218),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_207),
.B1(n_205),
.B2(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_202),
.B1(n_193),
.B2(n_206),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_156),
.B(n_178),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_187),
.C(n_143),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_188),
.B1(n_155),
.B2(n_143),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_233),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_210),
.B1(n_214),
.B2(n_218),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_219),
.B(n_210),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_241),
.B(n_223),
.Y(n_243)
);

AOI31xp67_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_209),
.A3(n_222),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_189),
.C(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_232),
.B(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_149),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_235),
.B1(n_224),
.B2(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_244),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_143),
.C(n_11),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_226),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_223),
.B1(n_225),
.B2(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_230),
.C(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_248),
.B(n_203),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_203),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_244),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_247),
.C(n_245),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_251),
.B(n_112),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_255),
.B(n_124),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_257),
.Y(n_260)
);


endmodule