module fake_jpeg_30111_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_20),
.B(n_26),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_93),
.Y(n_162)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_15),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_15),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_103),
.Y(n_153)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_43),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_129),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_57),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_156),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_141),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_56),
.B(n_48),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_45),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_42),
.B1(n_31),
.B2(n_33),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_33),
.B1(n_44),
.B2(n_32),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_49),
.B1(n_91),
.B2(n_77),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_104),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_49),
.B1(n_23),
.B2(n_44),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_49),
.B1(n_23),
.B2(n_44),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_46),
.Y(n_173)
);

BUFx4f_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_67),
.B1(n_19),
.B2(n_95),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_170),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_178),
.Y(n_229)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_164),
.Y(n_176)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_68),
.B1(n_96),
.B2(n_58),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_182),
.A2(n_183),
.B1(n_210),
.B2(n_211),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_70),
.B1(n_63),
.B2(n_66),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_186),
.Y(n_231)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_188),
.Y(n_253)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_192),
.Y(n_255)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_122),
.A2(n_111),
.B1(n_152),
.B2(n_90),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_111),
.A2(n_95),
.B1(n_31),
.B2(n_42),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_31),
.B1(n_42),
.B2(n_24),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_108),
.A2(n_35),
.B(n_21),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_200),
.A2(n_38),
.B(n_28),
.Y(n_271)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_201),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_48),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_208),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_207),
.B(n_212),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_115),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_213),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_142),
.A2(n_71),
.B1(n_89),
.B2(n_80),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_60),
.B1(n_75),
.B2(n_78),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_216),
.Y(n_261)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_218),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_106),
.A2(n_102),
.B1(n_79),
.B2(n_24),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_147),
.B1(n_146),
.B2(n_107),
.Y(n_242)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_221),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_46),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_120),
.B(n_28),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_223),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_156),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_129),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_239),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_120),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_228),
.A2(n_6),
.B(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_230),
.B(n_228),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_190),
.B(n_124),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_232),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_125),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_242),
.A2(n_109),
.B1(n_154),
.B2(n_220),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_125),
.B(n_162),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_194),
.B(n_196),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_183),
.A2(n_144),
.B(n_25),
.C(n_21),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_246),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_204),
.B1(n_189),
.B2(n_195),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_180),
.B(n_144),
.C(n_52),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_162),
.C(n_124),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_254),
.C(n_260),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_131),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_197),
.C(n_198),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_176),
.B(n_131),
.C(n_134),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_191),
.B(n_35),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_25),
.C(n_38),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_184),
.B1(n_136),
.B2(n_170),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_274),
.A2(n_298),
.B1(n_311),
.B2(n_231),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_275),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_276),
.A2(n_231),
.B(n_245),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_277),
.B(n_279),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_211),
.B1(n_182),
.B2(n_154),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_287),
.B1(n_297),
.B2(n_309),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_292),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_282),
.A2(n_284),
.B1(n_290),
.B2(n_299),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_199),
.B1(n_218),
.B2(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_223),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_296),
.Y(n_328)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_227),
.A2(n_202),
.B1(n_23),
.B2(n_32),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_180),
.B1(n_32),
.B2(n_184),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_294),
.B(n_260),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_227),
.A2(n_15),
.B1(n_52),
.B2(n_3),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_1),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_248),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_248),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_230),
.B(n_5),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_302),
.Y(n_340)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_230),
.B(n_6),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g351 ( 
.A(n_303),
.B(n_13),
.CI(n_14),
.CON(n_351),
.SN(n_351)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_232),
.B(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_307),
.Y(n_341)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_308),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_248),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_7),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_314),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_242),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_226),
.Y(n_312)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_228),
.B(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_14),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_12),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_313),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_244),
.A2(n_13),
.B1(n_14),
.B2(n_250),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_297),
.B1(n_309),
.B2(n_305),
.Y(n_338)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_318),
.A2(n_327),
.B(n_335),
.Y(n_368)
);

BUFx24_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_319),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_264),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_334),
.C(n_315),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_251),
.B(n_246),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_347),
.B(n_335),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_336),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_270),
.C(n_268),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_293),
.A2(n_267),
.B(n_236),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_354),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_312),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_291),
.Y(n_367)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_303),
.A2(n_255),
.B(n_253),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_293),
.A2(n_255),
.B1(n_258),
.B2(n_235),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_349),
.A2(n_324),
.B1(n_282),
.B2(n_326),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_351),
.A2(n_238),
.B(n_234),
.Y(n_388)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_294),
.B(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_357),
.Y(n_374)
);

XNOR2x2_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_279),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_358),
.A2(n_365),
.B(n_376),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_360),
.A2(n_369),
.B1(n_372),
.B2(n_375),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_377),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_283),
.Y(n_364)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_259),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_324),
.A2(n_349),
.B1(n_338),
.B2(n_346),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_278),
.B1(n_307),
.B2(n_277),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_379),
.B1(n_384),
.B2(n_392),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_323),
.A2(n_299),
.B1(n_280),
.B2(n_283),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_344),
.B1(n_320),
.B2(n_329),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_267),
.B(n_236),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g378 ( 
.A(n_354),
.B(n_302),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_378),
.A2(n_330),
.B1(n_350),
.B2(n_237),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_337),
.A2(n_306),
.B1(n_301),
.B2(n_314),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_296),
.B1(n_300),
.B2(n_235),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_381),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_328),
.A2(n_245),
.B1(n_253),
.B2(n_249),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_231),
.Y(n_382)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_269),
.Y(n_383)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_337),
.A2(n_243),
.B1(n_238),
.B2(n_269),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_234),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_331),
.C(n_333),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_247),
.Y(n_387)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_247),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_341),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_389),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_322),
.A2(n_243),
.B(n_237),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_319),
.B(n_265),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_331),
.A2(n_333),
.B1(n_321),
.B2(n_343),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_385),
.C(n_377),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_348),
.C(n_357),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_356),
.C(n_342),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_400),
.C(n_420),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_363),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_399),
.B(n_405),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_342),
.C(n_330),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_389),
.A2(n_351),
.B1(n_321),
.B2(n_353),
.Y(n_402)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_351),
.B1(n_353),
.B2(n_352),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_403),
.A2(n_392),
.B1(n_387),
.B2(n_370),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_419),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_361),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_361),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_410),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_408),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_266),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_350),
.Y(n_415)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

AO22x2_ASAP7_75t_L g416 ( 
.A1(n_358),
.A2(n_319),
.B1(n_233),
.B2(n_265),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_370),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_359),
.B(n_233),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_418),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_419),
.A2(n_376),
.B(n_384),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_266),
.C(n_272),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_272),
.C(n_259),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_362),
.Y(n_439)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_401),
.A2(n_360),
.B1(n_369),
.B2(n_375),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_425),
.A2(n_429),
.B1(n_437),
.B2(n_441),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_415),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_427),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_418),
.Y(n_433)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_416),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_439),
.Y(n_464)
);

OA22x2_ASAP7_75t_L g437 ( 
.A1(n_423),
.A2(n_358),
.B1(n_379),
.B2(n_368),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_394),
.B(n_380),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_440),
.B(n_444),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_372),
.B1(n_381),
.B2(n_388),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_447),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_414),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_448),
.B(n_414),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_450),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_451),
.A2(n_413),
.B1(n_404),
.B2(n_409),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_396),
.C(n_398),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_453),
.C(n_454),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_411),
.C(n_395),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_411),
.C(n_397),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_422),
.C(n_400),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_457),
.C(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_407),
.C(n_412),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_407),
.C(n_412),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_409),
.C(n_421),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_437),
.C(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_463),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_446),
.Y(n_466)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_466),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_449),
.B(n_393),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_468),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_423),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_459),
.Y(n_484)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_430),
.B1(n_447),
.B2(n_435),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_483),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_490),
.Y(n_501)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_484),
.B(n_464),
.Y(n_496)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_473),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_486),
.Y(n_495)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_467),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_488),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_489),
.B(n_467),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_425),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_452),
.C(n_453),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_497),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_478),
.A2(n_427),
.B1(n_470),
.B2(n_461),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_503),
.B1(n_506),
.B2(n_416),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_502),
.Y(n_509)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_475),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_462),
.B(n_457),
.Y(n_499)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_499),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_478),
.A2(n_430),
.B1(n_472),
.B2(n_428),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_481),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_455),
.C(n_464),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_487),
.B(n_393),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_451),
.C(n_445),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_484),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_480),
.A2(n_427),
.B1(n_429),
.B2(n_428),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_513),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_477),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_514),
.C(n_517),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_477),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_498),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_516),
.Y(n_525)
);

NOR2x1_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_413),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_474),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_506),
.C(n_505),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_522),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_510),
.A2(n_504),
.B(n_495),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_524),
.B(n_438),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_501),
.C(n_494),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_501),
.C(n_493),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_523),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_491),
.C(n_431),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_511),
.C(n_515),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_531),
.Y(n_534)
);

XNOR2x1_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_516),
.Y(n_530)
);

AOI31xp33_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_432),
.A3(n_443),
.B(n_374),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_529),
.A2(n_525),
.B(n_433),
.Y(n_532)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_432),
.B(n_374),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_528),
.B(n_386),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_536),
.C(n_386),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

AOI211xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_534),
.B(n_373),
.C(n_390),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_373),
.B(n_390),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_386),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_14),
.B(n_259),
.Y(n_542)
);


endmodule