module fake_jpeg_2653_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_2),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_48),
.B(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_2),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.C(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_52),
.B1(n_41),
.B2(n_43),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_55),
.B1(n_47),
.B2(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_55),
.B1(n_50),
.B2(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_56),
.B1(n_58),
.B2(n_46),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_59),
.B1(n_60),
.B2(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_88),
.B1(n_66),
.B2(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_51),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_99),
.C(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_40),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_78),
.C(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_116),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_80),
.B(n_60),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_119),
.C(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_80),
.B(n_49),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_122),
.B(n_8),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_72),
.B(n_71),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_99),
.B1(n_102),
.B2(n_89),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_60),
.B(n_20),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_111),
.C(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_136),
.C(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_108),
.B1(n_113),
.B2(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_135),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_23),
.B(n_37),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_22),
.C(n_36),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_21),
.C(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_132),
.B1(n_129),
.B2(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.C(n_145),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_137),
.B(n_127),
.Y(n_147)
);

AOI31xp67_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_10),
.A3(n_13),
.B(n_14),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_9),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_140),
.B(n_12),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_152),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_149),
.B1(n_13),
.B2(n_15),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_10),
.B(n_16),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_18),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_24),
.C(n_25),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_26),
.B(n_27),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_28),
.B(n_33),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_38),
.Y(n_161)
);


endmodule