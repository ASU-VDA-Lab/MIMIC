module fake_jpeg_16241_n_211 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_211);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_46),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_1),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_22),
.Y(n_53)
);

XNOR2x1_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_59),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_22),
.B1(n_18),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_56),
.B1(n_61),
.B2(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_18),
.B1(n_28),
.B2(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_49),
.B1(n_29),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_69),
.B1(n_76),
.B2(n_34),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_2),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_2),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_31),
.B1(n_19),
.B2(n_24),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_34),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_88),
.Y(n_109)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_35),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_17),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_50),
.B1(n_48),
.B2(n_39),
.Y(n_90)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_91),
.B1(n_50),
.B2(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_100),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_27),
.C(n_48),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_27),
.C(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_7),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_108),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_68),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_83),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_131),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_139),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_90),
.B1(n_73),
.B2(n_71),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_149),
.B1(n_77),
.B2(n_119),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_87),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_79),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_60),
.B1(n_77),
.B2(n_86),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_112),
.C(n_108),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_146),
.C(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_149),
.B1(n_137),
.B2(n_144),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_123),
.B1(n_113),
.B2(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_131),
.B1(n_9),
.B2(n_10),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_99),
.B(n_75),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_143),
.B(n_132),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_141),
.C(n_129),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_176),
.C(n_152),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_129),
.B(n_147),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_172),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_179),
.B(n_8),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_182),
.B(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_155),
.B(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_152),
.B1(n_154),
.B2(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_162),
.C(n_165),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_119),
.B1(n_12),
.B2(n_13),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_111),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_174),
.C(n_150),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_188),
.B1(n_170),
.B2(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_9),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_193),
.A2(n_181),
.B1(n_186),
.B2(n_157),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_81),
.C(n_16),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_99),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_194),
.C(n_15),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_202),
.C(n_208),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_202),
.Y(n_211)
);


endmodule