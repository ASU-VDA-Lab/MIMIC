module fake_jpeg_942_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_7),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_4),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_61),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_52),
.Y(n_91)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_80),
.B1(n_79),
.B2(n_61),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_73),
.B(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_63),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

OR2x4_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_65),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_60),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_114),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_75),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_82),
.B(n_65),
.C(n_62),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_68),
.B(n_55),
.C(n_57),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_120),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_73),
.B1(n_56),
.B2(n_54),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_53),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_1),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_59),
.B1(n_62),
.B2(n_50),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_136),
.B1(n_67),
.B2(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_74),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_133),
.B(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_59),
.B1(n_64),
.B2(n_51),
.Y(n_136)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_58),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_148),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_112),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_150),
.C(n_66),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_159),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_115),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_67),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_2),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_60),
.B1(n_66),
.B2(n_5),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_2),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_3),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_146),
.B(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_168),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_172),
.B(n_22),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_6),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_12),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_178),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_153),
.B(n_138),
.C(n_137),
.D(n_149),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_28),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_31),
.C(n_46),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_181),
.C(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_30),
.C(n_45),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_169),
.C(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_23),
.C(n_44),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_33),
.C(n_43),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_13),
.B(n_15),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_198),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_166),
.B1(n_176),
.B2(n_175),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

AOI22x1_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_167),
.B1(n_173),
.B2(n_164),
.Y(n_197)
);

NOR4xp25_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_16),
.C(n_17),
.D(n_18),
.Y(n_203)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_193),
.C(n_194),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_196),
.B(n_192),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_202),
.B(n_199),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_207),
.B(n_36),
.C(n_19),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_20),
.B1(n_34),
.B2(n_37),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_38),
.Y(n_213)
);


endmodule