module real_aes_8123_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_0), .A2(n_229), .B1(n_609), .B2(n_610), .Y(n_791) );
XOR2x2_ASAP7_75t_L g454 ( .A(n_1), .B(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_2), .A2(n_168), .B1(n_313), .B2(n_336), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_3), .A2(n_56), .B1(n_458), .B2(n_699), .Y(n_825) );
INVx1_ASAP7_75t_L g563 ( .A(n_4), .Y(n_563) );
AOI222xp33_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_24), .B1(n_221), .B2(n_401), .C1(n_476), .C2(n_477), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_6), .A2(n_233), .B1(n_389), .B2(n_400), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_7), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_8), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_9), .A2(n_166), .B1(n_427), .B2(n_463), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_10), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_11), .B(n_459), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_12), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g388 ( .A1(n_13), .A2(n_96), .B1(n_313), .B2(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_14), .A2(n_149), .B1(n_389), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_15), .A2(n_68), .B1(n_465), .B2(n_467), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_16), .A2(n_482), .B1(n_520), .B2(n_521), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_16), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_17), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_18), .A2(n_202), .B1(n_519), .B2(n_783), .Y(n_782) );
XOR2x2_ASAP7_75t_L g285 ( .A(n_19), .B(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_20), .A2(n_71), .B1(n_377), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_21), .A2(n_86), .B1(n_477), .B2(n_492), .Y(n_701) );
INVx1_ASAP7_75t_L g828 ( .A(n_22), .Y(n_828) );
AO22x2_ASAP7_75t_L g292 ( .A1(n_23), .A2(n_77), .B1(n_293), .B2(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g809 ( .A(n_23), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g396 ( .A1(n_25), .A2(n_94), .B1(n_121), .B2(n_397), .C1(n_399), .C2(n_401), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_26), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_27), .A2(n_144), .B1(n_550), .B2(n_710), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_28), .A2(n_188), .B1(n_473), .B2(n_517), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_29), .A2(n_227), .B1(n_392), .B2(n_393), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g746 ( .A1(n_30), .A2(n_84), .B1(n_250), .B2(n_403), .C1(n_447), .C2(n_562), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_31), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_32), .A2(n_180), .B1(n_403), .B2(n_449), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_33), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_34), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_35), .A2(n_36), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_37), .A2(n_47), .B1(n_426), .B2(n_603), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_38), .A2(n_209), .B1(n_362), .B2(n_463), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_39), .A2(n_151), .B1(n_377), .B2(n_378), .Y(n_376) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_40), .A2(n_80), .B1(n_293), .B2(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g810 ( .A(n_40), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_41), .A2(n_127), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_42), .A2(n_199), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_43), .A2(n_114), .B1(n_392), .B2(n_465), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_44), .A2(n_45), .B1(n_346), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_46), .A2(n_257), .B1(n_399), .B2(n_401), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_48), .B(n_458), .Y(n_642) );
INVx1_ASAP7_75t_L g733 ( .A(n_49), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_50), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_51), .A2(n_228), .B1(n_368), .B2(n_370), .Y(n_367) );
AOI22xp5_ASAP7_75t_SL g817 ( .A1(n_52), .A2(n_253), .B1(n_818), .B2(n_820), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_53), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_54), .A2(n_201), .B1(n_549), .B2(n_610), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_55), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_57), .Y(n_621) );
XOR2x2_ASAP7_75t_L g691 ( .A(n_58), .B(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_59), .A2(n_246), .B1(n_399), .B2(n_401), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_60), .B(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_61), .A2(n_226), .B1(n_345), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_62), .A2(n_256), .B1(n_403), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_63), .A2(n_208), .B1(n_427), .B2(n_436), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_64), .B(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_65), .A2(n_252), .B1(n_312), .B2(n_335), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_66), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_67), .A2(n_155), .B1(n_342), .B2(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_69), .A2(n_181), .B1(n_728), .B2(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_70), .A2(n_142), .B1(n_305), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_72), .A2(n_120), .B1(n_447), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_73), .A2(n_150), .B1(n_505), .B2(n_555), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_74), .A2(n_92), .B1(n_517), .B2(n_519), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_75), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_76), .A2(n_259), .B1(n_319), .B2(n_328), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_78), .A2(n_137), .B1(n_371), .B2(n_436), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_79), .A2(n_167), .B1(n_313), .B2(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_81), .A2(n_212), .B1(n_471), .B2(n_550), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_82), .A2(n_255), .B1(n_508), .B2(n_576), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_83), .A2(n_207), .B1(n_553), .B2(n_755), .Y(n_823) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_85), .A2(n_272), .B(n_280), .C(n_811), .Y(n_271) );
INVx1_ASAP7_75t_L g278 ( .A(n_87), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_88), .B(n_318), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_89), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_90), .B(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_91), .A2(n_182), .B1(n_473), .B2(n_519), .Y(n_651) );
INVx1_ASAP7_75t_L g275 ( .A(n_93), .Y(n_275) );
INVx1_ASAP7_75t_L g839 ( .A(n_95), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_97), .A2(n_203), .B1(n_471), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_98), .A2(n_139), .B1(n_471), .B2(n_555), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_99), .A2(n_231), .B1(n_371), .B2(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_100), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_101), .A2(n_187), .B1(n_342), .B2(n_345), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_102), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_103), .A2(n_118), .B1(n_463), .B2(n_519), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_104), .A2(n_171), .B1(n_344), .B2(n_427), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_105), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_106), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_107), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_108), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_109), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_110), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_111), .A2(n_197), .B1(n_514), .B2(n_515), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_112), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_113), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_115), .A2(n_126), .B1(n_392), .B2(n_393), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_116), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_117), .A2(n_159), .B1(n_400), .B2(n_403), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_119), .A2(n_123), .B1(n_389), .B2(n_400), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_122), .A2(n_244), .B1(n_465), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_124), .A2(n_264), .B1(n_471), .B2(n_473), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_125), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_128), .A2(n_813), .B1(n_830), .B2(n_831), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_128), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_129), .A2(n_196), .B1(n_371), .B2(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_130), .A2(n_163), .B1(n_370), .B2(n_549), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_131), .A2(n_242), .B1(n_331), .B2(n_335), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_132), .A2(n_193), .B1(n_351), .B2(n_354), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_133), .A2(n_195), .B1(n_354), .B2(n_432), .Y(n_431) );
AOI22x1_ASAP7_75t_L g593 ( .A1(n_134), .A2(n_594), .B1(n_629), .B2(n_630), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_134), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g764 ( .A1(n_135), .A2(n_174), .B1(n_211), .B2(n_290), .C1(n_500), .C2(n_565), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_136), .A2(n_265), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_138), .A2(n_245), .B1(n_354), .B2(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g279 ( .A(n_140), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_141), .A2(n_234), .B1(n_305), .B2(n_310), .Y(n_304) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_143), .A2(n_204), .B1(n_363), .B2(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_145), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_146), .A2(n_161), .B1(n_215), .B2(n_290), .C1(n_449), .C2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_147), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_148), .A2(n_247), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_152), .A2(n_165), .B1(n_381), .B2(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_153), .A2(n_219), .B1(n_360), .B2(n_363), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_154), .A2(n_237), .B1(n_492), .B2(n_640), .Y(n_759) );
AND2x6_ASAP7_75t_L g274 ( .A(n_156), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_156), .Y(n_803) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_157), .A2(n_224), .B1(n_293), .B2(n_297), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_158), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_160), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_162), .A2(n_225), .B1(n_380), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_164), .B(n_319), .Y(n_387) );
INVx1_ASAP7_75t_L g652 ( .A(n_169), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_170), .A2(n_223), .B1(n_393), .B2(n_574), .Y(n_732) );
XNOR2xp5_ASAP7_75t_L g653 ( .A(n_172), .B(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_173), .A2(n_175), .B1(n_674), .B2(n_675), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_176), .A2(n_263), .B1(n_378), .B2(n_518), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_177), .A2(n_525), .B1(n_526), .B2(n_556), .Y(n_524) );
CKINVDCx14_ASAP7_75t_R g556 ( .A(n_177), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_178), .A2(n_217), .B1(n_609), .B2(n_610), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_179), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_183), .A2(n_222), .B1(n_465), .B2(n_576), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_184), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_185), .B(n_459), .Y(n_643) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_186), .A2(n_236), .B1(n_293), .B2(n_294), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_189), .A2(n_240), .B1(n_518), .B2(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_190), .B(n_699), .Y(n_698) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_191), .B(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_192), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_194), .A2(n_200), .B1(n_436), .B2(n_576), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_198), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_205), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_206), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_210), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_213), .A2(n_766), .B1(n_792), .B2(n_793), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_213), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_214), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_216), .A2(n_266), .B1(n_336), .B2(n_565), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_218), .A2(n_260), .B1(n_709), .B2(n_710), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_220), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_224), .B(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_230), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_232), .A2(n_239), .B1(n_360), .B2(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_235), .Y(n_419) );
INVx1_ASAP7_75t_L g806 ( .A(n_236), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_238), .A2(n_267), .B1(n_668), .B2(n_699), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_241), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_243), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_248), .A2(n_251), .B1(n_344), .B2(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_249), .Y(n_695) );
INVx1_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_258), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_261), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_262), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_268), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_269), .B(n_319), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_270), .A2(n_413), .B1(n_451), .B2(n_452), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_270), .Y(n_451) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_275), .Y(n_802) );
OA21x2_ASAP7_75t_L g837 ( .A1(n_276), .A2(n_801), .B(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_588), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_280) );
INVxp67_ASAP7_75t_L g796 ( .A(n_281), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_407), .B2(n_408), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AO22x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_373), .B1(n_405), .B2(n_406), .Y(n_284) );
INVx2_ASAP7_75t_L g405 ( .A(n_285), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_339), .Y(n_286) );
NOR2xp33_ASAP7_75t_SL g287 ( .A(n_288), .B(n_316), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_303), .B(n_304), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx4_ASAP7_75t_L g398 ( .A(n_290), .Y(n_398) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_290), .Y(n_476) );
BUFx3_ASAP7_75t_L g562 ( .A(n_290), .Y(n_562) );
INVx2_ASAP7_75t_L g637 ( .A(n_290), .Y(n_637) );
AND2x6_ASAP7_75t_L g290 ( .A(n_291), .B(n_298), .Y(n_290) );
AND2x4_ASAP7_75t_L g313 ( .A(n_291), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g543 ( .A(n_291), .Y(n_543) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_292), .B(n_300), .Y(n_309) );
INVx2_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_295), .Y(n_297) );
OR2x2_ASAP7_75t_L g324 ( .A(n_296), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g329 ( .A(n_296), .B(n_325), .Y(n_329) );
INVx2_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
INVx1_ASAP7_75t_L g338 ( .A(n_296), .Y(n_338) );
AND2x6_ASAP7_75t_L g344 ( .A(n_298), .B(n_323), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_298), .B(n_349), .Y(n_353) );
AND2x4_ASAP7_75t_L g362 ( .A(n_298), .B(n_329), .Y(n_362) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g322 ( .A(n_299), .B(n_302), .Y(n_322) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g348 ( .A(n_300), .B(n_315), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_300), .B(n_302), .Y(n_357) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g308 ( .A(n_302), .Y(n_308) );
INVx1_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
BUFx2_ASAP7_75t_L g450 ( .A(n_305), .Y(n_450) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx12f_ASAP7_75t_L g403 ( .A(n_306), .Y(n_403) );
INVx1_ASAP7_75t_L g662 ( .A(n_306), .Y(n_662) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_306), .Y(n_776) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g333 ( .A(n_308), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g332 ( .A(n_309), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g336 ( .A(n_309), .B(n_337), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_309), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g447 ( .A(n_313), .Y(n_447) );
BUFx2_ASAP7_75t_SL g477 ( .A(n_313), .Y(n_477) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_313), .Y(n_640) );
INVx1_ASAP7_75t_L g544 ( .A(n_314), .Y(n_544) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_326), .C(n_330), .Y(n_316) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_319), .Y(n_668) );
INVx5_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g458 ( .A(n_320), .Y(n_458) );
INVx2_ASAP7_75t_L g569 ( .A(n_320), .Y(n_569) );
INVx4_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x6_ASAP7_75t_L g328 ( .A(n_322), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g369 ( .A(n_322), .B(n_349), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_322), .B(n_329), .Y(n_386) );
INVx1_ASAP7_75t_L g441 ( .A(n_322), .Y(n_441) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g440 ( .A(n_324), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g349 ( .A(n_325), .B(n_334), .Y(n_349) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_328), .Y(n_459) );
INVx1_ASAP7_75t_SL g670 ( .A(n_328), .Y(n_670) );
AND2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_348), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_331), .Y(n_495) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_332), .Y(n_400) );
BUFx2_ASAP7_75t_L g449 ( .A(n_332), .Y(n_449) );
BUFx4f_ASAP7_75t_SL g565 ( .A(n_332), .Y(n_565) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_332), .Y(n_660) );
INVx1_ASAP7_75t_L g540 ( .A(n_334), .Y(n_540) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g389 ( .A(n_336), .Y(n_389) );
INVx1_ASAP7_75t_L g493 ( .A(n_336), .Y(n_493) );
BUFx2_ASAP7_75t_L g666 ( .A(n_336), .Y(n_666) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x6_ASAP7_75t_L g372 ( .A(n_338), .B(n_357), .Y(n_372) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_358), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_350), .Y(n_340) );
INVx1_ASAP7_75t_L g676 ( .A(n_342), .Y(n_676) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx5_ASAP7_75t_SL g434 ( .A(n_343), .Y(n_434) );
INVx4_ASAP7_75t_L g505 ( .A(n_343), .Y(n_505) );
INVx2_ASAP7_75t_L g603 ( .A(n_343), .Y(n_603) );
INVx1_ASAP7_75t_L g763 ( .A(n_343), .Y(n_763) );
INVx11_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx11_ASAP7_75t_L g472 ( .A(n_344), .Y(n_472) );
BUFx4f_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
BUFx3_ASAP7_75t_L g463 ( .A(n_347), .Y(n_463) );
BUFx3_ASAP7_75t_L g518 ( .A(n_347), .Y(n_518) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_348), .B(n_349), .Y(n_422) );
AND2x4_ASAP7_75t_L g355 ( .A(n_349), .B(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g580 ( .A(n_352), .Y(n_580) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_353), .Y(n_392) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
BUFx2_ASAP7_75t_SL g728 ( .A(n_353), .Y(n_728) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
INVx1_ASAP7_75t_L g468 ( .A(n_355), .Y(n_468) );
BUFx3_ASAP7_75t_L g519 ( .A(n_355), .Y(n_519) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_355), .Y(n_553) );
BUFx2_ASAP7_75t_L g574 ( .A(n_355), .Y(n_574) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_355), .Y(n_707) );
AND2x2_ASAP7_75t_L g576 ( .A(n_356), .B(n_540), .Y(n_576) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_367), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
INVx2_ASAP7_75t_L g515 ( .A(n_361), .Y(n_515) );
INVx3_ASAP7_75t_L g555 ( .A(n_361), .Y(n_555) );
INVx6_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
BUFx3_ASAP7_75t_L g473 ( .A(n_362), .Y(n_473) );
BUFx3_ASAP7_75t_L g710 ( .A(n_362), .Y(n_710) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
INVx2_ASAP7_75t_L g436 ( .A(n_365), .Y(n_436) );
INVx5_ASAP7_75t_L g550 ( .A(n_365), .Y(n_550) );
INVx4_ASAP7_75t_L g819 ( .A(n_365), .Y(n_819) );
INVx8_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_368), .Y(n_600) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
INVx2_ASAP7_75t_L g466 ( .A(n_369), .Y(n_466) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_369), .Y(n_508) );
BUFx3_ASAP7_75t_L g581 ( .A(n_369), .Y(n_581) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g381 ( .A(n_371), .Y(n_381) );
BUFx2_ASAP7_75t_L g610 ( .A(n_371), .Y(n_610) );
BUFx2_ASAP7_75t_L g820 ( .A(n_371), .Y(n_820) );
INVx6_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g511 ( .A(n_372), .Y(n_511) );
INVx1_ASAP7_75t_SL g678 ( .A(n_372), .Y(n_678) );
INVx3_ASAP7_75t_SL g406 ( .A(n_373), .Y(n_406) );
XOR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_404), .Y(n_373) );
NAND4xp75_ASAP7_75t_L g374 ( .A(n_375), .B(n_382), .C(n_390), .D(n_396), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_379), .Y(n_375) );
OA211x2_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_387), .C(n_388), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_384), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_528) );
BUFx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g489 ( .A(n_386), .Y(n_489) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .Y(n_390) );
INVxp67_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
INVx2_ASAP7_75t_L g497 ( .A(n_397), .Y(n_497) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g533 ( .A(n_398), .Y(n_533) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx4f_ASAP7_75t_SL g500 ( .A(n_403), .Y(n_500) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_480), .B1(n_586), .B2(n_587), .Y(n_410) );
INVx1_ASAP7_75t_L g587 ( .A(n_411), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_453), .B1(n_478), .B2(n_479), .Y(n_411) );
INVx1_ASAP7_75t_L g478 ( .A(n_412), .Y(n_478) );
INVx2_ASAP7_75t_SL g452 ( .A(n_413), .Y(n_452) );
AND4x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_430), .C(n_437), .D(n_448), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_423), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_419), .B2(n_420), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g605 ( .A1(n_417), .A2(n_420), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_605) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_428), .B2(n_429), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g514 ( .A(n_427), .Y(n_514) );
INVx3_ASAP7_75t_L g597 ( .A(n_427), .Y(n_597) );
BUFx3_ASAP7_75t_L g790 ( .A(n_427), .Y(n_790) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_435), .Y(n_430) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_442), .B1(n_443), .B2(n_445), .C(n_446), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
BUFx3_ASAP7_75t_L g716 ( .A(n_440), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_443), .A2(n_485), .B1(n_769), .B2(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g479 ( .A(n_453), .Y(n_479) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND4xp75_ASAP7_75t_L g455 ( .A(n_456), .B(n_461), .C(n_469), .D(n_475), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_460), .Y(n_456) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g709 ( .A(n_472), .Y(n_709) );
INVx2_ASAP7_75t_L g619 ( .A(n_476), .Y(n_619) );
INVx2_ASAP7_75t_SL g657 ( .A(n_476), .Y(n_657) );
INVx1_ASAP7_75t_L g586 ( .A(n_480), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_522), .B1(n_523), .B2(n_585), .Y(n_480) );
INVx1_ASAP7_75t_SL g585 ( .A(n_481), .Y(n_585) );
INVx1_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_502), .Y(n_482) );
NOR2xp33_ASAP7_75t_SL g483 ( .A(n_484), .B(n_494), .Y(n_483) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_487), .B1(n_488), .B2(n_490), .C(n_491), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_485), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g530 ( .A(n_486), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_488), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g615 ( .A(n_489), .Y(n_615) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI222xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_497), .B2(n_498), .C1(n_499), .C2(n_501), .Y(n_494) );
OAI222xp33_ASAP7_75t_L g616 ( .A1(n_499), .A2(n_617), .B1(n_618), .B2(n_619), .C1(n_620), .C2(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
OAI221xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B1(n_507), .B2(n_509), .C(n_510), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g682 ( .A(n_507), .Y(n_682) );
INVx4_ASAP7_75t_L g755 ( .A(n_507), .Y(n_755) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_516), .Y(n_512) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g784 ( .A(n_518), .Y(n_784) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AO22x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_557), .B1(n_583), .B2(n_584), .Y(n_523) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_545), .Y(n_526) );
NOR3xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .C(n_536), .Y(n_527) );
OAI21xp5_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g827 ( .A1(n_533), .A2(n_828), .B(n_829), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B1(n_541), .B2(n_542), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_538), .A2(n_627), .B1(n_778), .B2(n_779), .Y(n_777) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g625 ( .A(n_539), .Y(n_625) );
BUFx3_ASAP7_75t_L g723 ( .A(n_539), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_542), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_542), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g609 ( .A(n_550), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVx3_ASAP7_75t_SL g583 ( .A(n_557), .Y(n_583) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_582), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_559), .B(n_571), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B(n_564), .Y(n_560) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_561), .A2(n_719), .B(n_720), .Y(n_718) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .C(n_570), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g797 ( .A(n_588), .Y(n_797) );
AOI22xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_590), .B1(n_749), .B2(n_750), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B1(n_686), .B2(n_687), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_631), .B1(n_684), .B2(n_685), .Y(n_592) );
INVx1_ASAP7_75t_L g684 ( .A(n_593), .Y(n_684) );
INVx1_ASAP7_75t_L g630 ( .A(n_594), .Y(n_630) );
AND2x2_ASAP7_75t_SL g594 ( .A(n_595), .B(n_611), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_605), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_601), .C(n_602), .Y(n_596) );
INVx2_ASAP7_75t_L g674 ( .A(n_597), .Y(n_674) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .C(n_622), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g771 ( .A1(n_617), .A2(n_657), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_626), .B2(n_627), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g685 ( .A(n_631), .Y(n_685) );
OA22x2_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B1(n_653), .B2(n_683), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
XOR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_652), .Y(n_633) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_645), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_641), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B(n_639), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .C(n_644), .Y(n_641) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g683 ( .A(n_653), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_671), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_664), .Y(n_655) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_661), .C1(n_662), .C2(n_663), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_657), .A2(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g699 ( .A(n_670), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_679), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B1(n_735), .B2(n_748), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_711), .B2(n_734), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_702), .C(n_705), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .C(n_701), .Y(n_697) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx3_ASAP7_75t_L g787 ( .A(n_710), .Y(n_787) );
INVx2_ASAP7_75t_SL g734 ( .A(n_711), .Y(n_734) );
XOR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_733), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_725), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .C(n_721), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_730), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx2_ASAP7_75t_SL g748 ( .A(n_735), .Y(n_748) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_747), .Y(n_735) );
NAND4xp75_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .C(n_743), .D(n_746), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_SL g740 ( .A(n_741), .B(n_742), .Y(n_740) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OA22x2_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_765), .B1(n_794), .B2(n_795), .Y(n_750) );
INVx1_ASAP7_75t_L g795 ( .A(n_751), .Y(n_795) );
NAND4xp75_ASAP7_75t_L g752 ( .A(n_753), .B(n_757), .C(n_760), .D(n_764), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
AND2x2_ASAP7_75t_SL g757 ( .A(n_758), .B(n_759), .Y(n_757) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g794 ( .A(n_765), .Y(n_794) );
INVx2_ASAP7_75t_L g793 ( .A(n_766), .Y(n_793) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_780), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .C(n_777), .Y(n_767) );
BUFx4f_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_788), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
NOR2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_804), .Y(n_799) );
OR2x2_ASAP7_75t_SL g844 ( .A(n_800), .B(n_805), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_801), .Y(n_833) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_802), .B(n_836), .Y(n_838) );
CKINVDCx16_ASAP7_75t_R g836 ( .A(n_803), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
OAI322xp33_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_832), .A3(n_834), .B1(n_837), .B2(n_839), .C1(n_840), .C2(n_842), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_813), .Y(n_831) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_814), .B(n_839), .Y(n_841) );
NOR4xp75_ASAP7_75t_L g814 ( .A(n_815), .B(n_821), .C(n_824), .D(n_827), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_816), .B(n_817), .Y(n_815) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_825), .B(n_826), .Y(n_824) );
BUFx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
endmodule