module fake_jpeg_6341_n_97 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_3),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_4),
.C(n_5),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_30),
.B(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx12_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_16),
.B(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_21),
.Y(n_41)
);

NOR4xp25_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_51),
.C(n_53),
.D(n_6),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_17),
.B(n_20),
.C(n_13),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_43),
.B(n_22),
.C(n_16),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_17),
.B(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_15),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_50),
.B1(n_40),
.B2(n_53),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_15),
.C(n_22),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_7),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_49),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_42),
.B1(n_39),
.B2(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_68),
.B1(n_75),
.B2(n_59),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_48),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_77),
.B1(n_55),
.B2(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_82),
.B1(n_62),
.B2(n_64),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_67),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.C(n_84),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_54),
.B(n_40),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_54),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_79),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_77),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_84),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_69),
.C(n_68),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_92),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_88),
.A3(n_80),
.B1(n_87),
.B2(n_86),
.C1(n_46),
.C2(n_35),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_92),
.B(n_35),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_96),
.B(n_44),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_46),
.B(n_11),
.C(n_44),
.Y(n_96)
);


endmodule