module fake_jpeg_20924_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_82),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx12f_ASAP7_75t_SL g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_88),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_56),
.B1(n_49),
.B2(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_63),
.B1(n_54),
.B2(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_91),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_61),
.A3(n_74),
.B1(n_62),
.B2(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_72),
.Y(n_121)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_51),
.C(n_57),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_73),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_53),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_68),
.B(n_75),
.C(n_72),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_123),
.B(n_22),
.C(n_47),
.D(n_45),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_93),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_75),
.A3(n_64),
.B1(n_12),
.B2(n_25),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_128),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_0),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_133),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_65),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_136),
.A2(n_60),
.B(n_21),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_116),
.B1(n_124),
.B2(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_110),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_145),
.B(n_126),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_20),
.A3(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_132),
.A3(n_133),
.B1(n_10),
.B2(n_29),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_151),
.B(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_141),
.B1(n_150),
.B2(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_44),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_39),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_30),
.C(n_24),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_2),
.B(n_4),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule