module fake_netlist_6_3263_n_1139 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_265, n_113, n_39, n_63, n_223, n_270, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1139);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_270;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1139;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_874;
wire n_480;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1071;
wire n_1042;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_284;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_685;
wire n_832;
wire n_280;
wire n_287;
wire n_597;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_691;
wire n_901;
wire n_535;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_842;
wire n_720;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_940;
wire n_770;
wire n_795;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_844;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_910;
wire n_911;
wire n_947;
wire n_381;
wire n_486;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_719;
wire n_565;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_683;
wire n_620;
wire n_420;
wire n_527;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_792;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_831;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_301;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_27),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_26),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_155),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_48),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_138),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_208),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_102),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_130),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_110),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_70),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_147),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_96),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_184),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_93),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_120),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_165),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_119),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_251),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_115),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_143),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_249),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_107),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_170),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_78),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_187),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_91),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_80),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_0),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_189),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_10),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_156),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_230),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_40),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_69),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_256),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_169),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_43),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_86),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_202),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_219),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_47),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_237),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_259),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_203),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_227),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_97),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_238),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_252),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_101),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_106),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_103),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_222),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_234),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_34),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_239),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_273),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_24),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_75),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_108),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_253),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_161),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_141),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_135),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_232),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_95),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_20),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_49),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_254),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_114),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_152),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_99),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_261),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_8),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_157),
.Y(n_366)
);

BUFx8_ASAP7_75t_SL g367 ( 
.A(n_60),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_63),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_258),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_58),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_248),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_268),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_112),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_34),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_36),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_118),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_128),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_100),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_154),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_207),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_150),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_160),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_45),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_79),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_88),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_217),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_192),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_66),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_61),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_158),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_151),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_270),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_164),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_179),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_200),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_213),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_19),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_64),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_15),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_28),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_206),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_131),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_46),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_137),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_1),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_271),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_14),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_127),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_20),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_94),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_28),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_35),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_116),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_134),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_176),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_76),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_111),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_89),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_191),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_246),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_81),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_55),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_83),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_146),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_193),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_218),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_38),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_54),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_16),
.Y(n_431)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_26),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_247),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_243),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_229),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_105),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_185),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_223),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_233),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_262),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_267),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_68),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_82),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_266),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_37),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_209),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_52),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_27),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_142),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_196),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_126),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_77),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_73),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_144),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_21),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_221),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_19),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_125),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_8),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_98),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_24),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_41),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_257),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_92),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_153),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_298),
.B(n_0),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_395),
.B(n_1),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_276),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_326),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_326),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_389),
.B(n_2),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_395),
.B(n_2),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_368),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_368),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_307),
.B(n_3),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_325),
.B(n_3),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_339),
.B(n_4),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_409),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_409),
.B(n_4),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_312),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_298),
.B(n_5),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_5),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_305),
.B(n_6),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_303),
.B(n_309),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_432),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_377),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_279),
.B(n_6),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_278),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_305),
.B(n_7),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_309),
.B(n_7),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_314),
.B(n_39),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_438),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_335),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_446),
.B(n_9),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_314),
.B(n_9),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_315),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_335),
.B(n_11),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_337),
.B(n_11),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_327),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_337),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_355),
.B(n_407),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_367),
.Y(n_520)
);

BUFx12f_ASAP7_75t_L g521 ( 
.A(n_286),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_383),
.B(n_12),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_403),
.B(n_13),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_327),
.Y(n_524)
);

BUFx8_ASAP7_75t_SL g525 ( 
.A(n_423),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_358),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_401),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_281),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_345),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_275),
.B(n_13),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_277),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_327),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_327),
.Y(n_536)
);

BUFx12f_ASAP7_75t_L g537 ( 
.A(n_348),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_280),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_283),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_327),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_285),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_414),
.B(n_14),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_327),
.B(n_15),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_287),
.B(n_16),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_448),
.B(n_451),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_365),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_374),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_288),
.B(n_17),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_293),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_282),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_296),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_304),
.B(n_17),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_289),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_400),
.B(n_18),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_408),
.B(n_18),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_410),
.B(n_21),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_413),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_308),
.B(n_22),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_431),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_313),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_316),
.B(n_22),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_319),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_324),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_328),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_329),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_332),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_334),
.B(n_23),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_336),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_340),
.Y(n_573)
);

NOR2x1_ASAP7_75t_L g574 ( 
.A(n_341),
.B(n_42),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_290),
.Y(n_575)
);

CKINVDCx6p67_ASAP7_75t_R g576 ( 
.A(n_284),
.Y(n_576)
);

BUFx12f_ASAP7_75t_L g577 ( 
.A(n_291),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_545),
.A2(n_330),
.B1(n_363),
.B2(n_320),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_474),
.A2(n_378),
.B1(n_426),
.B2(n_375),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_467),
.A2(n_433),
.B1(n_343),
.B2(n_344),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_489),
.A2(n_461),
.B1(n_457),
.B2(n_455),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_470),
.A2(n_477),
.B1(n_510),
.B2(n_485),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_482),
.A2(n_483),
.B1(n_481),
.B2(n_522),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_528),
.B(n_564),
.Y(n_584)
);

AO22x2_ASAP7_75t_L g585 ( 
.A1(n_467),
.A2(n_419),
.B1(n_351),
.B2(n_352),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_475),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_471),
.B(n_292),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_342),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_550),
.B(n_357),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_537),
.B(n_546),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_554),
.A2(n_437),
.B1(n_453),
.B2(n_442),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_508),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_475),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_550),
.B(n_359),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_R g597 ( 
.A1(n_484),
.A2(n_436),
.B1(n_391),
.B2(n_396),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_516),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_531),
.B(n_294),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_488),
.A2(n_454),
.B1(n_397),
.B2(n_405),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_523),
.A2(n_466),
.B1(n_465),
.B2(n_464),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_295),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_488),
.A2(n_387),
.B1(n_411),
.B2(n_416),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_297),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_542),
.A2(n_463),
.B1(n_459),
.B2(n_452),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_520),
.B(n_418),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_468),
.A2(n_450),
.B1(n_447),
.B2(n_445),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_555),
.A2(n_441),
.B1(n_443),
.B2(n_440),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_475),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_299),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_493),
.A2(n_439),
.B1(n_435),
.B2(n_430),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_559),
.B(n_300),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_525),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_575),
.B(n_301),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_493),
.A2(n_429),
.B1(n_428),
.B2(n_427),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_553),
.B(n_425),
.Y(n_620)
);

OA22x2_ASAP7_75t_L g621 ( 
.A1(n_487),
.A2(n_424),
.B1(n_422),
.B2(n_421),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_496),
.B(n_302),
.Y(n_622)
);

AO22x2_ASAP7_75t_L g623 ( 
.A1(n_490),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_476),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_551),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_577),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_509),
.B(n_306),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_496),
.B(n_310),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_504),
.A2(n_369),
.B1(n_415),
.B2(n_412),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_504),
.A2(n_417),
.B1(n_404),
.B2(n_402),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_570),
.A2(n_399),
.B1(n_394),
.B2(n_393),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_507),
.B(n_311),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_507),
.B(n_25),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_497),
.A2(n_390),
.B1(n_388),
.B2(n_386),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_557),
.B(n_29),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_502),
.A2(n_385),
.B1(n_384),
.B2(n_382),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_519),
.B(n_317),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_556),
.A2(n_381),
.B1(n_380),
.B2(n_379),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_469),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_519),
.B(n_318),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_511),
.A2(n_376),
.B1(n_373),
.B2(n_372),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_557),
.B(n_321),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_563),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_500),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_SL g648 ( 
.A1(n_543),
.A2(n_371),
.B1(n_370),
.B2(n_366),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

OA22x2_ASAP7_75t_L g651 ( 
.A1(n_526),
.A2(n_364),
.B1(n_362),
.B2(n_361),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_472),
.B(n_473),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_552),
.A2(n_360),
.B1(n_356),
.B2(n_354),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_563),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_503),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_571),
.A2(n_501),
.B1(n_490),
.B2(n_513),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_513),
.A2(n_338),
.B1(n_350),
.B2(n_349),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_561),
.A2(n_353),
.B1(n_347),
.B2(n_346),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_514),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_491),
.A2(n_333),
.B1(n_331),
.B2(n_323),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_473),
.B(n_322),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_643),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_652),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_579),
.B(n_576),
.Y(n_666)
);

XOR2x2_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_514),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_649),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_650),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_622),
.B(n_563),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_574),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_596),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_604),
.B(n_530),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_612),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_656),
.A2(n_533),
.B(n_544),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_633),
.B(n_567),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_640),
.B(n_492),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_624),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_626),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_632),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_583),
.A2(n_533),
.B(n_544),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_629),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_651),
.A2(n_548),
.B(n_558),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_647),
.B(n_515),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_582),
.B(n_567),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_644),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_655),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_662),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_586),
.Y(n_692)
);

BUFx2_ASAP7_75t_R g693 ( 
.A(n_620),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_593),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_598),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_614),
.B(n_567),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_606),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_599),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_517),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_548),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_603),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_661),
.B(n_517),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_621),
.A2(n_558),
.B(n_572),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_588),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_608),
.Y(n_705)
);

XOR2xp5_ASAP7_75t_L g706 ( 
.A(n_592),
.B(n_44),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_625),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_584),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_587),
.Y(n_710)
);

INVx4_ASAP7_75t_SL g711 ( 
.A(n_636),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_590),
.Y(n_712)
);

XOR2xp5_ASAP7_75t_L g713 ( 
.A(n_610),
.B(n_50),
.Y(n_713)
);

XOR2x2_ASAP7_75t_L g714 ( 
.A(n_634),
.B(n_30),
.Y(n_714)
);

XOR2xp5_ASAP7_75t_L g715 ( 
.A(n_648),
.B(n_51),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_587),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_638),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_613),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_636),
.B(n_505),
.Y(n_719)
);

XNOR2xp5_ASAP7_75t_L g720 ( 
.A(n_591),
.B(n_31),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_602),
.Y(n_721)
);

XOR2xp5_ASAP7_75t_L g722 ( 
.A(n_630),
.B(n_53),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_595),
.B(n_524),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_607),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

INVxp33_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_580),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_627),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_585),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_517),
.Y(n_731)
);

INVxp33_ASAP7_75t_L g732 ( 
.A(n_615),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_585),
.Y(n_733)
);

XOR2xp5_ASAP7_75t_L g734 ( 
.A(n_631),
.B(n_56),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_591),
.B(n_32),
.Y(n_735)
);

XOR2xp5_ASAP7_75t_L g736 ( 
.A(n_639),
.B(n_57),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_601),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_635),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_618),
.B(n_562),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_601),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_605),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_605),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_618),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_657),
.B(n_573),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_712),
.B(n_637),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_718),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_723),
.B(n_642),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_723),
.B(n_653),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_664),
.B(n_658),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_683),
.A2(n_660),
.B(n_611),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_663),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_683),
.A2(n_505),
.B(n_540),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_707),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_664),
.B(n_518),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_700),
.B(n_623),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_676),
.B(n_702),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_700),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_738),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_676),
.B(n_518),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_689),
.B(n_732),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_708),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_668),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_699),
.B(n_518),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_687),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_670),
.B(n_518),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_678),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_739),
.B(n_623),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_681),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_690),
.Y(n_773)
);

OAI21xp33_ASAP7_75t_L g774 ( 
.A1(n_745),
.A2(n_532),
.B(n_527),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_691),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_677),
.B(n_505),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_678),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_669),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_744),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_703),
.B(n_659),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_673),
.B(n_505),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_717),
.B(n_646),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_719),
.B(n_659),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_725),
.B(n_704),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_693),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_566),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_741),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_710),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_685),
.A2(n_566),
.B(n_568),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_674),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_697),
.B(n_654),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_685),
.B(n_568),
.Y(n_793)
);

AND2x2_ASAP7_75t_SL g794 ( 
.A(n_719),
.B(n_478),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_726),
.B(n_479),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_679),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_688),
.B(n_534),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_680),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_684),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_692),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_728),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_665),
.B(n_696),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_730),
.B(n_512),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_512),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_737),
.Y(n_808)
);

AND2x2_ASAP7_75t_SL g809 ( 
.A(n_731),
.B(n_478),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_740),
.B(n_609),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_695),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_742),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_698),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_701),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_672),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_709),
.B(n_534),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_711),
.B(n_609),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_711),
.B(n_529),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_711),
.B(n_529),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_729),
.B(n_534),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_706),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_721),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_682),
.B(n_589),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_764),
.B(n_667),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_819),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_819),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_770),
.B(n_724),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_760),
.B(n_589),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_777),
.B(n_736),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_777),
.B(n_538),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_819),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_783),
.B(n_713),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_754),
.B(n_538),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_805),
.B(n_666),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_780),
.B(n_759),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_820),
.B(n_671),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_760),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_820),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_798),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_818),
.B(n_722),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_778),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_778),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_760),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_806),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_784),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_818),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_766),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_783),
.B(n_734),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_786),
.B(n_715),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_803),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_754),
.B(n_538),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_757),
.B(n_763),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_768),
.B(n_560),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_498),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_766),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_768),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_765),
.B(n_59),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_761),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_750),
.B(n_560),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_812),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_786),
.B(n_714),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_766),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_749),
.B(n_560),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_810),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_809),
.B(n_498),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_758),
.B(n_565),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_765),
.B(n_62),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_758),
.B(n_565),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_761),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_789),
.B(n_65),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_809),
.B(n_565),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_788),
.B(n_67),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_823),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_779),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_773),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_747),
.B(n_748),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_789),
.B(n_479),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_746),
.B(n_569),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_753),
.B(n_71),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_808),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_842),
.Y(n_883)
);

BUFx8_ASAP7_75t_SL g884 ( 
.A(n_841),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_866),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_878),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_842),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_828),
.A2(n_822),
.B1(n_751),
.B2(n_752),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_843),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_843),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_871),
.Y(n_891)
);

OR2x6_ASAP7_75t_SL g892 ( 
.A(n_830),
.B(n_822),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_875),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_847),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_848),
.Y(n_895)
);

INVx6_ASAP7_75t_L g896 ( 
.A(n_847),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_841),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_868),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

BUFx2_ASAP7_75t_R g900 ( 
.A(n_826),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_871),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_867),
.B(n_794),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_837),
.Y(n_903)
);

BUFx12f_ASAP7_75t_L g904 ( 
.A(n_829),
.Y(n_904)
);

BUFx4_ASAP7_75t_SL g905 ( 
.A(n_868),
.Y(n_905)
);

INVx8_ASAP7_75t_L g906 ( 
.A(n_847),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_836),
.A2(n_780),
.B1(n_794),
.B2(n_771),
.Y(n_907)
);

BUFx4_ASAP7_75t_SL g908 ( 
.A(n_870),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_840),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_852),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_862),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_860),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_827),
.Y(n_913)
);

INVx3_ASAP7_75t_SL g914 ( 
.A(n_829),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_832),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_863),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_846),
.B(n_790),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_825),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_877),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_857),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_858),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_836),
.A2(n_771),
.B1(n_755),
.B2(n_807),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_858),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_857),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_838),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_906),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_906),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_902),
.A2(n_836),
.B1(n_867),
.B2(n_850),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_897),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_883),
.Y(n_931)
);

INVx6_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_902),
.A2(n_859),
.B1(n_869),
.B2(n_881),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_894),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_922),
.B(n_924),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_893),
.Y(n_936)
);

INVx6_ASAP7_75t_L g937 ( 
.A(n_896),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_922),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_916),
.A2(n_849),
.B1(n_833),
.B2(n_835),
.Y(n_939)
);

BUFx8_ASAP7_75t_L g940 ( 
.A(n_885),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_889),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_904),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_907),
.A2(n_859),
.B1(n_869),
.B2(n_881),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_891),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_896),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_901),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_909),
.Y(n_947)
);

INVx6_ASAP7_75t_L g948 ( 
.A(n_896),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_883),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_886),
.B(n_919),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_910),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_921),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_888),
.A2(n_849),
.B1(n_833),
.B2(n_916),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_907),
.A2(n_793),
.B1(n_808),
.B2(n_873),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_917),
.A2(n_836),
.B1(n_839),
.B2(n_874),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_894),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_895),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_887),
.Y(n_959)
);

HB1xp67_ASAP7_75t_SL g960 ( 
.A(n_900),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_890),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_890),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_912),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_923),
.A2(n_880),
.B1(n_861),
.B2(n_865),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_952),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_939),
.A2(n_597),
.B1(n_923),
.B2(n_880),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_953),
.A2(n_892),
.B1(n_882),
.B2(n_876),
.Y(n_968)
);

BUFx4f_ASAP7_75t_SL g969 ( 
.A(n_940),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_931),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_939),
.A2(n_903),
.B1(n_808),
.B2(n_897),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_935),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_930),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_SL g974 ( 
.A1(n_929),
.A2(n_762),
.B1(n_720),
.B2(n_735),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_960),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_950),
.B(n_845),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_929),
.A2(n_823),
.B1(n_874),
.B2(n_824),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_951),
.B(n_772),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_936),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_943),
.A2(n_824),
.B1(n_903),
.B2(n_898),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_SL g981 ( 
.A1(n_943),
.A2(n_785),
.B(n_774),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_933),
.A2(n_911),
.B1(n_913),
.B2(n_915),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_960),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_930),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_933),
.A2(n_955),
.B1(n_956),
.B2(n_964),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_942),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_947),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_937),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_964),
.A2(n_915),
.B1(n_913),
.B2(n_821),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_941),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_955),
.A2(n_814),
.B1(n_802),
.B2(n_811),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_937),
.A2(n_762),
.B1(n_904),
.B2(n_792),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_963),
.A2(n_802),
.B1(n_811),
.B2(n_813),
.Y(n_993)
);

BUFx4f_ASAP7_75t_SL g994 ( 
.A(n_927),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_SL g995 ( 
.A1(n_932),
.A2(n_810),
.B1(n_782),
.B2(n_799),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_938),
.A2(n_814),
.B1(n_813),
.B2(n_773),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_L g997 ( 
.A1(n_935),
.A2(n_804),
.B(n_792),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_937),
.B(n_914),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_934),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_944),
.A2(n_920),
.B1(n_853),
.B2(n_855),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_948),
.A2(n_851),
.B1(n_864),
.B2(n_914),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_948),
.A2(n_796),
.B1(n_870),
.B2(n_787),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_974),
.A2(n_775),
.B1(n_884),
.B2(n_756),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_967),
.A2(n_800),
.B1(n_795),
.B2(n_946),
.Y(n_1004)
);

OA21x2_ASAP7_75t_L g1005 ( 
.A1(n_985),
.A2(n_776),
.B(n_834),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_967),
.A2(n_800),
.B1(n_795),
.B2(n_775),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_976),
.B(n_949),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_970),
.Y(n_1008)
);

OAI222xp33_ASAP7_75t_L g1009 ( 
.A1(n_980),
.A2(n_962),
.B1(n_961),
.B2(n_959),
.C1(n_954),
.C2(n_831),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_990),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_SL g1011 ( 
.A1(n_971),
.A2(n_932),
.B1(n_948),
.B2(n_934),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_972),
.B(n_945),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_977),
.A2(n_968),
.B1(n_995),
.B2(n_997),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_SL g1014 ( 
.A1(n_982),
.A2(n_932),
.B1(n_957),
.B2(n_934),
.Y(n_1014)
);

OAI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_981),
.A2(n_796),
.B1(n_791),
.B2(n_815),
.C(n_769),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_989),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_1002),
.B(n_816),
.C(n_797),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_SL g1018 ( 
.A1(n_992),
.A2(n_957),
.B(n_884),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_969),
.A2(n_957),
.B1(n_928),
.B2(n_927),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_978),
.A2(n_979),
.B1(n_973),
.B2(n_991),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_966),
.A2(n_756),
.B1(n_797),
.B2(n_854),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_969),
.A2(n_756),
.B1(n_854),
.B2(n_801),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_987),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1000),
.A2(n_945),
.B1(n_927),
.B2(n_928),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_975),
.A2(n_801),
.B1(n_815),
.B2(n_807),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_1000),
.A2(n_789),
.B1(n_817),
.B2(n_872),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_993),
.A2(n_983),
.B1(n_984),
.B2(n_996),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_SL g1028 ( 
.A1(n_999),
.A2(n_806),
.B1(n_998),
.B2(n_905),
.C(n_908),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_994),
.A2(n_928),
.B1(n_851),
.B2(n_864),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_986),
.A2(n_817),
.B1(n_872),
.B2(n_838),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1001),
.A2(n_844),
.B1(n_838),
.B2(n_857),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_988),
.A2(n_994),
.B1(n_926),
.B2(n_965),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_965),
.A2(n_844),
.B1(n_781),
.B2(n_926),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_974),
.A2(n_844),
.B1(n_925),
.B2(n_958),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_974),
.A2(n_952),
.B1(n_958),
.B2(n_921),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_974),
.A2(n_925),
.B1(n_767),
.B2(n_569),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_974),
.A2(n_569),
.B1(n_918),
.B2(n_895),
.Y(n_1037)
);

AOI222xp33_ASAP7_75t_L g1038 ( 
.A1(n_974),
.A2(n_535),
.B1(n_536),
.B2(n_33),
.C1(n_530),
.C2(n_918),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1010),
.B(n_33),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1038),
.A2(n_856),
.B(n_879),
.Y(n_1040)
);

OAI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_1004),
.A2(n_918),
.B1(n_895),
.B2(n_899),
.C(n_536),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1007),
.B(n_899),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1023),
.B(n_899),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1016),
.B(n_1023),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_1013),
.B(n_536),
.C(n_535),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1012),
.B(n_899),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1004),
.A2(n_921),
.B1(n_530),
.B2(n_535),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1008),
.B(n_72),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1006),
.B(n_74),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1006),
.A2(n_921),
.B1(n_495),
.B2(n_486),
.Y(n_1050)
);

OAI221xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1003),
.A2(n_1036),
.B1(n_1037),
.B2(n_1018),
.C(n_1020),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1014),
.B(n_85),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1011),
.B(n_87),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1005),
.B(n_90),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_1035),
.A2(n_104),
.B(n_109),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1015),
.A2(n_495),
.B(n_486),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1034),
.B(n_1032),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_1025),
.B(n_495),
.C(n_486),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1027),
.A2(n_113),
.B(n_117),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1005),
.B(n_121),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1005),
.B(n_122),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1024),
.B(n_123),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1017),
.B(n_124),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_L g1064 ( 
.A(n_1044),
.B(n_1009),
.Y(n_1064)
);

AOI221xp5_ASAP7_75t_L g1065 ( 
.A1(n_1051),
.A2(n_1028),
.B1(n_1022),
.B2(n_1021),
.C(n_1019),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_L g1066 ( 
.A(n_1051),
.B(n_1029),
.C(n_1030),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1043),
.B(n_1031),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1046),
.B(n_1026),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1059),
.A2(n_1033),
.B1(n_480),
.B2(n_479),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_129),
.B(n_132),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1057),
.B(n_136),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_1054),
.Y(n_1072)
);

NAND4xp75_ASAP7_75t_L g1073 ( 
.A(n_1061),
.B(n_139),
.C(n_140),
.D(n_145),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1045),
.A2(n_480),
.B1(n_149),
.B2(n_159),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1055),
.A2(n_480),
.B1(n_162),
.B2(n_163),
.Y(n_1075)
);

BUFx2_ASAP7_75t_SL g1076 ( 
.A(n_1071),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_1064),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1072),
.B(n_1061),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1067),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1070),
.B(n_1060),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_1042),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1070),
.Y(n_1082)
);

XNOR2xp5_ASAP7_75t_L g1083 ( 
.A(n_1065),
.B(n_1039),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1073),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1069),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1078),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1078),
.Y(n_1087)
);

XOR2x2_ASAP7_75t_L g1088 ( 
.A(n_1083),
.B(n_1066),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1079),
.B(n_1077),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1082),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_1081),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1081),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1092),
.Y(n_1093)
);

OA22x2_ASAP7_75t_L g1094 ( 
.A1(n_1089),
.A2(n_1084),
.B1(n_1076),
.B2(n_1080),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1086),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1091),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_1087),
.Y(n_1097)
);

OA22x2_ASAP7_75t_SL g1098 ( 
.A1(n_1088),
.A2(n_1084),
.B1(n_1085),
.B2(n_1082),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1090),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_1090),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1092),
.Y(n_1101)
);

OA22x2_ASAP7_75t_L g1102 ( 
.A1(n_1089),
.A2(n_1080),
.B1(n_1085),
.B2(n_1075),
.Y(n_1102)
);

OA22x2_ASAP7_75t_L g1103 ( 
.A1(n_1098),
.A2(n_1100),
.B1(n_1099),
.B2(n_1096),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_SL g1104 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1095),
.Y(n_1105)
);

OAI322xp33_ASAP7_75t_L g1106 ( 
.A1(n_1102),
.A2(n_1052),
.A3(n_1053),
.B1(n_1063),
.B2(n_1049),
.C1(n_1062),
.C2(n_1041),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1095),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1094),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_1103),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_1097),
.B1(n_1058),
.B2(n_1056),
.Y(n_1110)
);

NAND4xp25_ASAP7_75t_L g1111 ( 
.A(n_1104),
.B(n_1074),
.C(n_1040),
.D(n_1048),
.Y(n_1111)
);

AND4x1_ASAP7_75t_L g1112 ( 
.A(n_1105),
.B(n_1107),
.C(n_1106),
.D(n_1047),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_1106),
.A2(n_1050),
.B1(n_166),
.B2(n_167),
.Y(n_1113)
);

AND4x1_ASAP7_75t_L g1114 ( 
.A(n_1103),
.B(n_148),
.C(n_168),
.D(n_171),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1109),
.A2(n_173),
.B1(n_177),
.B2(n_181),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1110),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1113),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1114),
.A2(n_182),
.B(n_183),
.C(n_186),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1116),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_1111),
.B1(n_1112),
.B2(n_194),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1115),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1119),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1121),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_1120),
.B(n_1118),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_188),
.B1(n_190),
.B2(n_195),
.Y(n_1125)
);

NAND5xp2_ASAP7_75t_L g1126 ( 
.A(n_1123),
.B(n_197),
.C(n_198),
.D(n_199),
.E(n_201),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1125),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1127),
.A2(n_1122),
.B1(n_1126),
.B2(n_211),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1128),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1129),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_204),
.B1(n_210),
.B2(n_212),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1131),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1130),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1133),
.Y(n_1135)
);

AOI31xp33_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_1134),
.A3(n_1132),
.B(n_236),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1136),
.Y(n_1137)
);

AOI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_226),
.B1(n_231),
.B2(n_240),
.C(n_241),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1138),
.A2(n_272),
.B1(n_244),
.B2(n_245),
.Y(n_1139)
);


endmodule