module fake_jpeg_19342_n_319 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_32),
.B1(n_21),
.B2(n_13),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_44),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_53),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_43),
.B1(n_38),
.B2(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_37),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_19),
.B(n_11),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_45),
.B1(n_24),
.B2(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_15),
.B1(n_12),
.B2(n_21),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_34),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_61),
.Y(n_89)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_85),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_51),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_96),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_66),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_79),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_97),
.B(n_79),
.Y(n_113)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_22),
.B(n_11),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_50),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_79),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_63),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_83),
.B1(n_96),
.B2(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_123),
.B1(n_99),
.B2(n_69),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_105),
.B(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_88),
.C(n_69),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_113),
.B(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_124),
.B(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_12),
.Y(n_155)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_69),
.C(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_29),
.C(n_17),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_64),
.B1(n_78),
.B2(n_77),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_88),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_131),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_122),
.B1(n_121),
.B2(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_71),
.B1(n_97),
.B2(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_143),
.B1(n_144),
.B2(n_52),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_163),
.Y(n_174)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_150),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_152),
.B1(n_159),
.B2(n_129),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_95),
.B1(n_80),
.B2(n_75),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_75),
.B1(n_94),
.B2(n_63),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_113),
.B1(n_117),
.B2(n_114),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_65),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_65),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_94),
.B1(n_51),
.B2(n_57),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_160),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_111),
.A2(n_60),
.B1(n_12),
.B2(n_21),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_52),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_166),
.B(n_176),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_182),
.B1(n_194),
.B2(n_142),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_114),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_171),
.A2(n_20),
.B(n_16),
.Y(n_218)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_163),
.B1(n_135),
.B2(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_178),
.B1(n_144),
.B2(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_191),
.B1(n_137),
.B2(n_139),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_108),
.B1(n_110),
.B2(n_61),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_22),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_17),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_22),
.B1(n_19),
.B2(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_198),
.B(n_201),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_157),
.C(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_209),
.C(n_217),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_211),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_182),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_140),
.B1(n_134),
.B2(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_156),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_171),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_148),
.B1(n_132),
.B2(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_146),
.C(n_148),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_152),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_136),
.B1(n_153),
.B2(n_18),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_153),
.B1(n_18),
.B2(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_17),
.C(n_28),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_172),
.C(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_224),
.C(n_228),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_197),
.A3(n_241),
.B1(n_222),
.B2(n_226),
.C1(n_195),
.C2(n_240),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_185),
.C(n_192),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_171),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_226),
.A2(n_203),
.B(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_207),
.C(n_214),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_190),
.C(n_184),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_239),
.C(n_205),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_184),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_169),
.B(n_165),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_165),
.C(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_212),
.B1(n_206),
.B2(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_196),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_225),
.B1(n_235),
.B2(n_236),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_253),
.B1(n_254),
.B2(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_230),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_228),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_17),
.C(n_14),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_213),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_258),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_197),
.B1(n_183),
.B2(n_167),
.Y(n_259)
);

AOI22x1_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_220),
.B1(n_167),
.B2(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_270),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_229),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_248),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_220),
.C(n_17),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.C(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_260),
.C(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_245),
.C(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_281),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_257),
.B1(n_274),
.B2(n_244),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_8),
.B1(n_7),
.B2(n_2),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_254),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_249),
.B(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_27),
.C(n_14),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_14),
.B(n_27),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_14),
.C(n_20),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_10),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_0),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_9),
.B(n_8),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_292),
.B(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_9),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_293),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_20),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_295),
.A3(n_16),
.B1(n_1),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_0),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_7),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_0),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_0),
.B(n_1),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.Y(n_311)
);

NAND5xp2_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_16),
.C(n_20),
.D(n_2),
.E(n_3),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_308),
.C(n_1),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_307),
.B(n_289),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_312),
.A3(n_302),
.B(n_304),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_311),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_303),
.A3(n_16),
.B1(n_5),
.B2(n_6),
.C1(n_4),
.C2(n_1),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_4),
.C(n_5),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_4),
.C(n_6),
.Y(n_318)
);

AOI211xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_4),
.B(n_6),
.C(n_290),
.Y(n_319)
);


endmodule