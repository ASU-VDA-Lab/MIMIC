module real_aes_8208_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_156;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g459 ( .A1(n_0), .A2(n_139), .B(n_460), .C(n_463), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_1), .B(n_454), .Y(n_465) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g177 ( .A(n_3), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_4), .B(n_140), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_5), .A2(n_118), .B1(n_119), .B2(n_425), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_5), .Y(n_425) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_5), .A2(n_94), .B1(n_425), .B2(n_726), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_6), .A2(n_439), .B(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_7), .A2(n_146), .B(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_8), .A2(n_37), .B1(n_143), .B2(n_195), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_9), .B(n_146), .Y(n_163) );
AND2x6_ASAP7_75t_L g148 ( .A(n_10), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_11), .A2(n_148), .B(n_442), .C(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_38), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_12), .B(n_38), .Y(n_732) );
INVx1_ASAP7_75t_L g130 ( .A(n_13), .Y(n_130) );
INVx1_ASAP7_75t_L g169 ( .A(n_14), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_15), .B(n_136), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_16), .B(n_140), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_17), .B(n_126), .Y(n_125) );
AO32x2_ASAP7_75t_L g206 ( .A1(n_18), .A2(n_146), .A3(n_147), .B1(n_166), .B2(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_19), .B(n_143), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_20), .B(n_126), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_21), .A2(n_52), .B1(n_143), .B2(n_195), .Y(n_209) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_22), .A2(n_77), .B1(n_136), .B2(n_143), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_23), .B(n_143), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_24), .A2(n_147), .B(n_442), .C(n_444), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_25), .A2(n_147), .B(n_442), .C(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_26), .Y(n_134) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_27), .A2(n_35), .B1(n_116), .B2(n_715), .C1(n_717), .C2(n_718), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_27), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_28), .B(n_185), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_29), .A2(n_439), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_30), .B(n_185), .Y(n_222) );
INVx2_ASAP7_75t_L g138 ( .A(n_31), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_32), .A2(n_474), .B(n_475), .C(n_479), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_33), .B(n_143), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_34), .B(n_185), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_36), .B(n_191), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_39), .B(n_438), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_40), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_41), .B(n_140), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_42), .B(n_439), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_43), .A2(n_474), .B(n_479), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_44), .B(n_143), .Y(n_156) );
INVx1_ASAP7_75t_L g461 ( .A(n_45), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_46), .A2(n_87), .B1(n_195), .B2(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g500 ( .A(n_47), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_48), .B(n_143), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_49), .B(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_50), .B(n_439), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_51), .B(n_161), .Y(n_160) );
AOI22xp33_ASAP7_75t_SL g142 ( .A1(n_53), .A2(n_57), .B1(n_136), .B2(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_54), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_55), .B(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_56), .B(n_143), .Y(n_242) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_59), .B(n_439), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_60), .B(n_454), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_61), .A2(n_161), .B(n_172), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_62), .B(n_143), .Y(n_178) );
INVx1_ASAP7_75t_L g129 ( .A(n_63), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_64), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_65), .B(n_140), .Y(n_477) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_66), .A2(n_146), .A3(n_147), .B1(n_200), .B2(n_204), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_67), .B(n_141), .Y(n_511) );
INVx1_ASAP7_75t_L g241 ( .A(n_68), .Y(n_241) );
INVx1_ASAP7_75t_L g217 ( .A(n_69), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_70), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_71), .B(n_446), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_72), .A2(n_442), .B(n_479), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_73), .B(n_136), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_74), .Y(n_487) );
INVx1_ASAP7_75t_L g736 ( .A(n_75), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_76), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_78), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_79), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_80), .B(n_136), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g100 ( .A1(n_81), .A2(n_101), .B1(n_728), .B2(n_737), .Y(n_100) );
INVx2_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_83), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_84), .B(n_133), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_85), .B(n_136), .Y(n_157) );
OR2x2_ASAP7_75t_L g110 ( .A(n_86), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g428 ( .A(n_86), .B(n_112), .Y(n_428) );
INVx2_ASAP7_75t_L g714 ( .A(n_86), .Y(n_714) );
NAND3xp33_ASAP7_75t_SL g733 ( .A(n_86), .B(n_113), .C(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_88), .A2(n_99), .B1(n_136), .B2(n_137), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_89), .B(n_439), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_90), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_91), .Y(n_107) );
INVxp67_ASAP7_75t_L g490 ( .A(n_92), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_93), .B(n_136), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_94), .Y(n_726) );
INVx1_ASAP7_75t_L g507 ( .A(n_95), .Y(n_507) );
INVx1_ASAP7_75t_L g536 ( .A(n_96), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_97), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g502 ( .A(n_98), .B(n_185), .Y(n_502) );
AOI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_115), .B1(n_721), .B2(n_722), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g721 ( .A(n_104), .Y(n_721) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_106), .A2(n_723), .B(n_727), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g727 ( .A(n_109), .Y(n_727) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_111), .B(n_714), .Y(n_720) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g713 ( .A(n_112), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_426), .B1(n_429), .B2(n_711), .Y(n_116) );
INVx1_ASAP7_75t_L g716 ( .A(n_117), .Y(n_716) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g724 ( .A(n_119), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_359), .Y(n_119) );
NOR5xp2_ASAP7_75t_L g120 ( .A(n_121), .B(n_272), .C(n_318), .D(n_331), .E(n_343), .Y(n_120) );
OAI211xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_180), .B(n_226), .C(n_253), .Y(n_121) );
INVx1_ASAP7_75t_SL g354 ( .A(n_122), .Y(n_354) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_150), .Y(n_122) );
AND2x2_ASAP7_75t_L g278 ( .A(n_123), .B(n_151), .Y(n_278) );
AND2x2_ASAP7_75t_L g306 ( .A(n_123), .B(n_252), .Y(n_306) );
AND2x2_ASAP7_75t_L g314 ( .A(n_123), .B(n_257), .Y(n_314) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g244 ( .A(n_124), .B(n_152), .Y(n_244) );
INVx2_ASAP7_75t_L g256 ( .A(n_124), .Y(n_256) );
AND2x2_ASAP7_75t_L g381 ( .A(n_124), .B(n_323), .Y(n_381) );
OR2x2_ASAP7_75t_L g383 ( .A(n_124), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_131), .Y(n_124) );
INVx1_ASAP7_75t_L g250 ( .A(n_125), .Y(n_250) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
INVx1_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_127), .B(n_128), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
NAND3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_145), .C(n_147), .Y(n_131) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_132), .A2(n_145), .B(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .B1(n_139), .B2(n_142), .Y(n_132) );
INVx2_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_133), .A2(n_141), .B1(n_201), .B2(n_203), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_133), .A2(n_139), .B1(n_208), .B2(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g462 ( .A(n_133), .Y(n_462) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx3_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
INVx1_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
AND2x2_ASAP7_75t_L g440 ( .A(n_134), .B(n_162), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_134), .Y(n_443) );
INVx2_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_139), .A2(n_159), .B(n_160), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_139), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_140), .A2(n_156), .B(n_157), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_SL g215 ( .A1(n_140), .A2(n_216), .B(n_217), .C(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_140), .A2(n_238), .B(n_239), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_140), .B(n_490), .Y(n_489) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_143), .Y(n_538) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
BUFx3_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
AND2x6_ASAP7_75t_L g442 ( .A(n_144), .B(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g454 ( .A(n_145), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_145), .B(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_145), .A2(n_506), .B(n_513), .Y(n_505) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_145), .A2(n_533), .B(n_540), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_145), .B(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_146), .A2(n_154), .B(n_163), .Y(n_153) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_146), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_146), .A2(n_518), .B(n_519), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_147), .A2(n_237), .B(n_240), .Y(n_236) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_148), .A2(n_155), .B(n_158), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_148), .A2(n_168), .B(n_175), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_148), .A2(n_187), .B(n_192), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_148), .A2(n_215), .B(n_219), .Y(n_214) );
AND2x4_ASAP7_75t_L g439 ( .A(n_148), .B(n_440), .Y(n_439) );
INVx4_ASAP7_75t_SL g464 ( .A(n_148), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_148), .B(n_440), .Y(n_508) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g294 ( .A(n_151), .B(n_266), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_151), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g408 ( .A(n_151), .B(n_248), .Y(n_408) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_164), .Y(n_151) );
AND2x2_ASAP7_75t_L g251 ( .A(n_152), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g298 ( .A(n_152), .Y(n_298) );
AND2x2_ASAP7_75t_L g323 ( .A(n_152), .B(n_235), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_152), .B(n_356), .Y(n_393) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g257 ( .A(n_153), .B(n_235), .Y(n_257) );
AND2x2_ASAP7_75t_L g271 ( .A(n_153), .B(n_234), .Y(n_271) );
AND2x2_ASAP7_75t_L g288 ( .A(n_153), .B(n_164), .Y(n_288) );
AND2x2_ASAP7_75t_L g345 ( .A(n_153), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_153), .B(n_252), .Y(n_358) );
AND2x2_ASAP7_75t_L g410 ( .A(n_153), .B(n_335), .Y(n_410) );
INVx2_ASAP7_75t_L g176 ( .A(n_161), .Y(n_176) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g233 ( .A(n_164), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g252 ( .A(n_164), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_164), .B(n_235), .Y(n_329) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_179), .Y(n_164) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_165), .A2(n_236), .B(n_243), .Y(n_235) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_166), .B(n_514), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_172), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_170), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_170), .A2(n_521), .B(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_172), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_173), .A2(n_220), .B(n_221), .Y(n_219) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g446 ( .A(n_174), .Y(n_446) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_176), .A2(n_196), .B(n_241), .C(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_176), .A2(n_445), .B(n_447), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_210), .B(n_223), .Y(n_180) );
INVx1_ASAP7_75t_SL g342 ( .A(n_181), .Y(n_342) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_198), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_183), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
INVx1_ASAP7_75t_L g262 ( .A(n_184), .Y(n_262) );
AND2x2_ASAP7_75t_L g283 ( .A(n_184), .B(n_205), .Y(n_283) );
AND2x2_ASAP7_75t_L g317 ( .A(n_184), .B(n_206), .Y(n_317) );
OR2x2_ASAP7_75t_L g336 ( .A(n_184), .B(n_212), .Y(n_336) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_184), .Y(n_350) );
AND2x2_ASAP7_75t_L g363 ( .A(n_184), .B(n_364), .Y(n_363) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_197), .Y(n_184) );
INVx2_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_185), .A2(n_214), .B(n_222), .Y(n_213) );
INVx1_ASAP7_75t_L g452 ( .A(n_185), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_185), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_185), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_198), .A2(n_285), .B1(n_286), .B2(n_295), .Y(n_284) );
AND2x2_ASAP7_75t_L g368 ( .A(n_198), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
INVx1_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_199), .Y(n_266) );
INVx1_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
AND2x2_ASAP7_75t_L g292 ( .A(n_199), .B(n_206), .Y(n_292) );
INVx2_ASAP7_75t_L g463 ( .A(n_202), .Y(n_463) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_202), .Y(n_478) );
INVx1_ASAP7_75t_L g449 ( .A(n_204), .Y(n_449) );
OR2x2_ASAP7_75t_L g246 ( .A(n_205), .B(n_231), .Y(n_246) );
AND2x2_ASAP7_75t_L g276 ( .A(n_205), .B(n_277), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_205), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g224 ( .A(n_206), .B(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g333 ( .A(n_206), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_210), .B(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g311 ( .A(n_211), .B(n_277), .Y(n_311) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g223 ( .A(n_212), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g282 ( .A(n_212), .Y(n_282) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
OR2x2_ASAP7_75t_L g261 ( .A(n_213), .B(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_213), .Y(n_316) );
AOI32xp33_ASAP7_75t_L g353 ( .A1(n_223), .A2(n_283), .A3(n_354), .B1(n_355), .B2(n_357), .Y(n_353) );
AND2x2_ASAP7_75t_L g279 ( .A(n_224), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_224), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_224), .B(n_311), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_224), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_232), .B1(n_245), .B2(n_247), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g332 ( .A(n_228), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_229), .B(n_231), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_254), .B1(n_258), .B2(n_268), .Y(n_253) );
AND2x2_ASAP7_75t_L g275 ( .A(n_230), .B(n_276), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_230), .A2(n_244), .B(n_292), .C(n_327), .Y(n_326) );
OAI332xp33_ASAP7_75t_L g331 ( .A1(n_230), .A2(n_332), .A3(n_334), .B1(n_336), .B2(n_337), .B3(n_339), .C1(n_340), .C2(n_342), .Y(n_331) );
INVx2_ASAP7_75t_L g372 ( .A(n_230), .Y(n_372) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_231), .Y(n_290) );
INVx1_ASAP7_75t_L g365 ( .A(n_231), .Y(n_365) );
AND2x2_ASAP7_75t_L g419 ( .A(n_231), .B(n_283), .Y(n_419) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_244), .Y(n_232) );
AND2x2_ASAP7_75t_L g299 ( .A(n_234), .B(n_249), .Y(n_299) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g347 ( .A(n_235), .B(n_249), .Y(n_347) );
INVx1_ASAP7_75t_L g356 ( .A(n_235), .Y(n_356) );
INVx1_ASAP7_75t_L g330 ( .A(n_244), .Y(n_330) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g414 ( .A(n_246), .B(n_266), .Y(n_414) );
INVx1_ASAP7_75t_SL g325 ( .A(n_247), .Y(n_325) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
AND2x2_ASAP7_75t_L g352 ( .A(n_248), .B(n_310), .Y(n_352) );
INVx1_ASAP7_75t_L g371 ( .A(n_248), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_248), .B(n_338), .Y(n_373) );
INVx1_ASAP7_75t_L g270 ( .A(n_249), .Y(n_270) );
AND2x2_ASAP7_75t_L g274 ( .A(n_251), .B(n_255), .Y(n_274) );
AND2x2_ASAP7_75t_L g341 ( .A(n_251), .B(n_299), .Y(n_341) );
INVx2_ASAP7_75t_L g384 ( .A(n_251), .Y(n_384) );
INVx2_ASAP7_75t_L g267 ( .A(n_252), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_252), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_256), .B(n_329), .Y(n_335) );
OR2x2_ASAP7_75t_L g399 ( .A(n_256), .B(n_358), .Y(n_399) );
INVx1_ASAP7_75t_L g423 ( .A(n_256), .Y(n_423) );
INVx1_ASAP7_75t_L g379 ( .A(n_257), .Y(n_379) );
AND2x2_ASAP7_75t_L g424 ( .A(n_257), .B(n_267), .Y(n_424) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_261), .A2(n_287), .B1(n_289), .B2(n_293), .Y(n_286) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI322xp33_ASAP7_75t_SL g370 ( .A1(n_264), .A2(n_371), .A3(n_372), .B1(n_373), .B2(n_374), .C1(n_377), .C2(n_379), .Y(n_370) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
AND2x2_ASAP7_75t_L g367 ( .A(n_265), .B(n_283), .Y(n_367) );
OR2x2_ASAP7_75t_L g401 ( .A(n_265), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_265), .B(n_336), .Y(n_404) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g349 ( .A(n_266), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g405 ( .A(n_266), .B(n_336), .Y(n_405) );
INVx3_ASAP7_75t_L g338 ( .A(n_267), .Y(n_338) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g394 ( .A(n_269), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g273 ( .A1(n_271), .A2(n_274), .B1(n_275), .B2(n_278), .C1(n_279), .C2(n_281), .Y(n_273) );
INVx1_ASAP7_75t_L g304 ( .A(n_271), .Y(n_304) );
NAND3xp33_ASAP7_75t_SL g272 ( .A(n_273), .B(n_284), .C(n_301), .Y(n_272) );
AND2x2_ASAP7_75t_L g389 ( .A(n_276), .B(n_290), .Y(n_389) );
BUFx2_ASAP7_75t_L g280 ( .A(n_277), .Y(n_280) );
INVx1_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_278), .A2(n_314), .B1(n_367), .B2(n_368), .C(n_370), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_280), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
AND2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_288), .B(n_299), .Y(n_300) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_290), .A2(n_296), .B(n_300), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_290), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g387 ( .A(n_292), .B(n_369), .Y(n_387) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_299), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g416 ( .A(n_299), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .B1(n_308), .B2(n_311), .C(n_312), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_303), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g412 ( .A(n_311), .B(n_317), .Y(n_412) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OAI31xp33_ASAP7_75t_SL g380 ( .A1(n_315), .A2(n_354), .A3(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_317), .B(n_321), .Y(n_420) );
OAI221xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_322), .B1(n_324), .B2(n_325), .C(n_326), .Y(n_318) );
INVx1_ASAP7_75t_L g324 ( .A(n_320), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_323), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g339 ( .A(n_332), .Y(n_339) );
INVx2_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g361 ( .A(n_338), .B(n_347), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_338), .A2(n_355), .B(n_412), .C(n_413), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g343 ( .A1(n_339), .A2(n_344), .B1(n_348), .B2(n_351), .C(n_353), .Y(n_343) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_342), .A2(n_407), .B(n_409), .C(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_345), .A2(n_396), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_395) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NOR4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_385), .C(n_406), .D(n_417), .Y(n_359) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B(n_366), .C(n_380), .Y(n_360) );
INVx1_ASAP7_75t_SL g415 ( .A(n_367), .Y(n_415) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_376), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_383), .A2(n_392), .B1(n_404), .B2(n_405), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_390), .C(n_395), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI31xp33_ASAP7_75t_L g417 ( .A1(n_388), .A2(n_418), .A3(n_420), .B(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_428), .A2(n_430), .B1(n_713), .B2(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_431), .B(n_647), .Y(n_430) );
NOR5xp2_ASAP7_75t_L g431 ( .A(n_432), .B(n_578), .C(n_607), .D(n_627), .E(n_634), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_466), .B(n_523), .C(n_565), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_434), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_649) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_453), .Y(n_434) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_435), .Y(n_526) );
AND2x4_ASAP7_75t_L g558 ( .A(n_435), .B(n_559), .Y(n_558) );
INVx5_ASAP7_75t_L g576 ( .A(n_435), .Y(n_576) );
AND2x2_ASAP7_75t_L g585 ( .A(n_435), .B(n_577), .Y(n_585) );
AND2x2_ASAP7_75t_L g597 ( .A(n_435), .B(n_470), .Y(n_597) );
AND2x2_ASAP7_75t_L g693 ( .A(n_435), .B(n_561), .Y(n_693) );
OR2x6_ASAP7_75t_L g435 ( .A(n_436), .B(n_450), .Y(n_435) );
AOI21xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_441), .B(n_449), .Y(n_436) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx5_ASAP7_75t_L g458 ( .A(n_442), .Y(n_458) );
INVx2_ASAP7_75t_L g448 ( .A(n_446), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_448), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_448), .A2(n_478), .B(n_500), .C(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g559 ( .A(n_453), .Y(n_559) );
AND2x2_ASAP7_75t_L g577 ( .A(n_453), .B(n_532), .Y(n_577) );
AND2x2_ASAP7_75t_L g596 ( .A(n_453), .B(n_531), .Y(n_596) );
AND2x2_ASAP7_75t_L g636 ( .A(n_453), .B(n_576), .Y(n_636) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_465), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B(n_459), .C(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g474 ( .A(n_458), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_458), .A2(n_464), .B(n_487), .C(n_488), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g479 ( .A(n_464), .Y(n_479) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_492), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_469), .A2(n_503), .A3(n_550), .B1(n_558), .B2(n_612), .C1(n_696), .C2(n_699), .Y(n_695) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_482), .Y(n_469) );
INVx5_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
AND2x2_ASAP7_75t_L g544 ( .A(n_470), .B(n_530), .Y(n_544) );
BUFx2_ASAP7_75t_L g622 ( .A(n_470), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_470), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g699 ( .A(n_470), .B(n_606), .Y(n_699) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_482), .B(n_494), .Y(n_553) );
INVx1_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_482), .B(n_515), .Y(n_593) );
AND2x2_ASAP7_75t_L g694 ( .A(n_482), .B(n_612), .Y(n_694) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g548 ( .A(n_483), .B(n_494), .Y(n_548) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_483), .Y(n_556) );
OR2x2_ASAP7_75t_L g563 ( .A(n_483), .B(n_515), .Y(n_563) );
AND2x2_ASAP7_75t_L g573 ( .A(n_483), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_483), .B(n_505), .Y(n_602) );
INVxp67_ASAP7_75t_L g626 ( .A(n_483), .Y(n_626) );
AND2x2_ASAP7_75t_L g633 ( .A(n_483), .B(n_503), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_483), .B(n_515), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_483), .B(n_504), .Y(n_659) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B(n_491), .Y(n_483) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_494), .B(n_516), .Y(n_603) );
OR2x2_ASAP7_75t_L g625 ( .A(n_494), .B(n_504), .Y(n_625) );
AND2x2_ASAP7_75t_L g638 ( .A(n_494), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_494), .B(n_593), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_494), .A2(n_649), .B(n_654), .C(n_663), .Y(n_648) );
AND2x2_ASAP7_75t_L g709 ( .A(n_494), .B(n_515), .Y(n_709) );
INVx5_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_495), .B(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_495), .B(n_557), .Y(n_569) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
OR2x2_ASAP7_75t_L g582 ( .A(n_495), .B(n_504), .Y(n_582) );
AND2x2_ASAP7_75t_SL g587 ( .A(n_495), .B(n_573), .Y(n_587) );
AND2x2_ASAP7_75t_L g612 ( .A(n_495), .B(n_504), .Y(n_612) );
AND2x2_ASAP7_75t_L g632 ( .A(n_495), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g670 ( .A(n_495), .B(n_503), .Y(n_670) );
OR2x2_ASAP7_75t_L g673 ( .A(n_495), .B(n_659), .Y(n_673) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_504), .A2(n_617), .B(n_620), .C(n_626), .Y(n_616) );
INVx5_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_505), .B(n_515), .Y(n_547) );
AND2x2_ASAP7_75t_L g551 ( .A(n_505), .B(n_516), .Y(n_551) );
OR2x2_ASAP7_75t_L g557 ( .A(n_505), .B(n_515), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_SL g574 ( .A(n_515), .Y(n_574) );
OR2x2_ASAP7_75t_L g702 ( .A(n_515), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_542), .B(n_545), .C(n_554), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI31xp33_ASAP7_75t_L g627 ( .A1(n_525), .A2(n_628), .A3(n_630), .B(n_631), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_526), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_527), .B(n_558), .Y(n_564) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_528), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g584 ( .A(n_528), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_528), .B(n_559), .Y(n_589) );
AND2x2_ASAP7_75t_L g599 ( .A(n_528), .B(n_558), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_528), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g619 ( .A(n_528), .B(n_576), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_528), .B(n_596), .Y(n_624) );
OR2x2_ASAP7_75t_L g643 ( .A(n_528), .B(n_530), .Y(n_643) );
OR2x2_ASAP7_75t_L g645 ( .A(n_528), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_528), .Y(n_692) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g592 ( .A(n_530), .B(n_559), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_530), .B(n_576), .Y(n_615) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g561 ( .A(n_532), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g652 ( .A(n_544), .B(n_576), .Y(n_652) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_544), .A2(n_558), .A3(n_596), .B1(n_655), .B2(n_656), .C1(n_657), .C2(n_660), .Y(n_654) );
INVx1_ASAP7_75t_L g662 ( .A(n_544), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx1_ASAP7_75t_SL g656 ( .A(n_546), .Y(n_656) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
OR2x2_ASAP7_75t_L g608 ( .A(n_547), .B(n_553), .Y(n_608) );
INVx1_ASAP7_75t_L g639 ( .A(n_547), .Y(n_639) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI32xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .A3(n_560), .B1(n_562), .B2(n_564), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI21xp33_ASAP7_75t_SL g594 ( .A1(n_557), .A2(n_572), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g609 ( .A(n_558), .Y(n_609) );
AND2x4_ASAP7_75t_L g606 ( .A(n_559), .B(n_576), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_559), .B(n_642), .Y(n_641) );
AOI322xp5_ASAP7_75t_L g671 ( .A1(n_560), .A2(n_587), .A3(n_606), .B1(n_639), .B2(n_672), .C1(n_674), .C2(n_675), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_560), .A2(n_637), .B1(n_701), .B2(n_702), .C(n_704), .Y(n_700) );
AND2x2_ASAP7_75t_L g588 ( .A(n_561), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g568 ( .A(n_563), .Y(n_568) );
OR2x2_ASAP7_75t_L g640 ( .A(n_563), .B(n_625), .Y(n_640) );
OAI31xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .A3(n_570), .B(n_575), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_566), .A2(n_599), .B1(n_600), .B2(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g611 ( .A(n_568), .B(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_570), .A2(n_611), .B1(n_664), .B2(n_667), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g653 ( .A(n_573), .B(n_622), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_573), .B(n_612), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_574), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g687 ( .A(n_574), .B(n_625), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_575), .A2(n_670), .B1(n_683), .B2(n_686), .Y(n_682) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g591 ( .A(n_576), .Y(n_591) );
AND2x2_ASAP7_75t_L g674 ( .A(n_576), .B(n_596), .Y(n_674) );
OR2x2_ASAP7_75t_L g676 ( .A(n_576), .B(n_643), .Y(n_676) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_576), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_577), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_577), .B(n_622), .Y(n_630) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_586), .C(n_598), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_590), .B2(n_593), .C(n_594), .Y(n_586) );
INVxp67_ASAP7_75t_L g698 ( .A(n_589), .Y(n_698) );
INVx1_ASAP7_75t_L g665 ( .A(n_590), .Y(n_665) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g629 ( .A(n_591), .B(n_596), .Y(n_629) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_592), .B(n_619), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g661 ( .A(n_596), .Y(n_661) );
AND2x2_ASAP7_75t_L g667 ( .A(n_596), .B(n_622), .Y(n_667) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g655 ( .A(n_603), .Y(n_655) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_606), .B(n_642), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_610), .B2(n_613), .C(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g703 ( .A(n_612), .Y(n_703) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g621 ( .A(n_615), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_619), .B(n_678), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B(n_625), .Y(n_620) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_623), .A2(n_669), .B(n_671), .C(n_677), .Y(n_668) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g680 ( .A(n_625), .Y(n_680) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_640), .B2(n_641), .C1(n_644), .C2(n_645), .Y(n_634) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g710 ( .A(n_641), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_642), .B(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_642), .A2(n_689), .B1(n_691), .B2(n_694), .Y(n_688) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
NOR4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_668), .C(n_681), .D(n_700), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_650), .B(n_680), .Y(n_690) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g657 ( .A(n_655), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_658), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_688), .C(n_695), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx2_ASAP7_75t_L g697 ( .A(n_693), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_710), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx12_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_731), .Y(n_737) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
endmodule