module real_aes_15559_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1402 ( .A1(n_0), .A2(n_72), .B1(n_609), .B2(n_614), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_0), .A2(n_224), .B1(n_546), .B2(n_697), .Y(n_1412) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_1), .A2(n_5), .B1(n_1132), .B2(n_1135), .Y(n_1174) );
INVx1_ASAP7_75t_L g1002 ( .A(n_2), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_2), .A2(n_95), .B1(n_546), .B2(n_738), .Y(n_1019) );
INVx1_ASAP7_75t_L g1353 ( .A(n_3), .Y(n_1353) );
INVx1_ASAP7_75t_L g1406 ( .A(n_4), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_6), .A2(n_110), .B1(n_675), .B2(n_678), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_6), .A2(n_114), .B1(n_545), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_7), .A2(n_73), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_7), .A2(n_52), .B1(n_639), .B2(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g264 ( .A(n_8), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_8), .B(n_274), .Y(n_296) );
AND2x2_ASAP7_75t_L g513 ( .A(n_8), .B(n_198), .Y(n_513) );
AND2x2_ASAP7_75t_L g531 ( .A(n_8), .B(n_417), .Y(n_531) );
INVx1_ASAP7_75t_L g298 ( .A(n_9), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g1400 ( .A1(n_10), .A2(n_126), .B1(n_606), .B2(n_1397), .C(n_1401), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_10), .A2(n_60), .B1(n_546), .B2(n_861), .Y(n_1414) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_11), .A2(n_137), .B1(n_625), .B2(n_673), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_11), .A2(n_16), .B1(n_534), .B2(n_541), .C(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_12), .A2(n_118), .B1(n_474), .B2(n_478), .Y(n_473) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_12), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_13), .A2(n_131), .B1(n_738), .B2(n_741), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_13), .A2(n_229), .B1(n_474), .B2(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_14), .Y(n_1088) );
INVx2_ASAP7_75t_L g1128 ( .A(n_15), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_15), .B(n_99), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_15), .B(n_1134), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_16), .A2(n_33), .B1(n_490), .B2(n_620), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g1394 ( .A(n_17), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_18), .A2(n_215), .B1(n_478), .B2(n_488), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_18), .A2(n_118), .B1(n_534), .B2(n_536), .C(n_540), .Y(n_533) );
INVx1_ASAP7_75t_L g670 ( .A(n_19), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_20), .A2(n_183), .B1(n_492), .B2(n_499), .Y(n_684) );
INVx1_ASAP7_75t_L g700 ( .A(n_20), .Y(n_700) );
INVx1_ASAP7_75t_L g1093 ( .A(n_21), .Y(n_1093) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_22), .A2(n_205), .B1(n_1132), .B2(n_1135), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_23), .A2(n_207), .B1(n_518), .B2(n_522), .Y(n_517) );
XOR2x2_ASAP7_75t_L g278 ( .A(n_24), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_25), .A2(n_71), .B1(n_474), .B2(n_1004), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_25), .A2(n_247), .B1(n_535), .B2(n_541), .C(n_859), .Y(n_1018) );
INVx1_ASAP7_75t_L g732 ( .A(n_26), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_26), .A2(n_214), .B1(n_518), .B2(n_522), .Y(n_761) );
INVx1_ASAP7_75t_L g1022 ( .A(n_27), .Y(n_1022) );
INVx1_ASAP7_75t_L g1042 ( .A(n_28), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_28), .A2(n_147), .B1(n_492), .B2(n_781), .Y(n_1059) );
INVx1_ASAP7_75t_L g1021 ( .A(n_29), .Y(n_1021) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_30), .A2(n_55), .B1(n_557), .B2(n_657), .C(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1067 ( .A(n_30), .Y(n_1067) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_31), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_32), .A2(n_247), .B1(n_474), .B2(n_1004), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_32), .A2(n_71), .B1(n_543), .B2(n_1028), .Y(n_1027) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_33), .A2(n_656), .B(n_704), .C(n_711), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_34), .A2(n_234), .B1(n_1125), .B2(n_1145), .Y(n_1144) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_35), .B(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_35), .A2(n_138), .B1(n_478), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_36), .A2(n_138), .B1(n_529), .B2(n_740), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_36), .A2(n_218), .B1(n_478), .B2(n_490), .Y(n_884) );
INVx1_ASAP7_75t_L g1344 ( .A(n_37), .Y(n_1344) );
INVx1_ASAP7_75t_L g324 ( .A(n_38), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_39), .A2(n_57), .B1(n_518), .B2(n_599), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_39), .A2(n_691), .B(n_692), .C(n_698), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_40), .A2(n_219), .B1(n_1132), .B2(n_1135), .Y(n_1148) );
INVx1_ASAP7_75t_L g985 ( .A(n_41), .Y(n_985) );
AO22x1_ASAP7_75t_L g1124 ( .A1(n_41), .A2(n_59), .B1(n_1125), .B2(n_1129), .Y(n_1124) );
XOR2x2_ASAP7_75t_L g450 ( .A(n_42), .B(n_451), .Y(n_450) );
XNOR2x2_ASAP7_75t_L g664 ( .A(n_43), .B(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_44), .A2(n_116), .B1(n_617), .B2(n_618), .Y(n_616) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_44), .Y(n_654) );
INVx1_ASAP7_75t_L g808 ( .A(n_45), .Y(n_808) );
INVx1_ASAP7_75t_L g338 ( .A(n_46), .Y(n_338) );
INVx1_ASAP7_75t_L g345 ( .A(n_46), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_47), .A2(n_122), .B1(n_1307), .B2(n_1309), .Y(n_1306) );
OAI22xp33_ASAP7_75t_L g1337 ( .A1(n_47), .A2(n_122), .B1(n_266), .B2(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g841 ( .A(n_48), .Y(n_841) );
INVx1_ASAP7_75t_L g992 ( .A(n_49), .Y(n_992) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_50), .A2(n_152), .B1(n_492), .B2(n_499), .Y(n_491) );
INVx1_ASAP7_75t_L g549 ( .A(n_50), .Y(n_549) );
INVxp67_ASAP7_75t_SL g1033 ( .A(n_51), .Y(n_1033) );
AND4x1_ASAP7_75t_L g1069 ( .A(n_51), .B(n_1035), .C(n_1038), .D(n_1057), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_52), .A2(n_123), .B1(n_609), .B2(n_613), .Y(n_612) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_53), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_53), .A2(n_117), .B1(n_483), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_54), .A2(n_114), .B1(n_678), .B2(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_54), .A2(n_110), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g1068 ( .A(n_55), .Y(n_1068) );
INVx1_ASAP7_75t_L g257 ( .A(n_56), .Y(n_257) );
INVx2_ASAP7_75t_L g331 ( .A(n_58), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_60), .A2(n_68), .B1(n_620), .B2(n_1397), .C(n_1398), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_61), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g767 ( .A(n_61), .Y(n_767) );
INVx1_ASAP7_75t_L g623 ( .A(n_62), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_63), .A2(n_78), .B1(n_797), .B2(n_799), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_63), .A2(n_203), .B1(n_738), .B2(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g1389 ( .A(n_64), .Y(n_1389) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_65), .A2(n_156), .B1(n_1125), .B2(n_1129), .Y(n_1149) );
INVx1_ASAP7_75t_L g1388 ( .A(n_66), .Y(n_1388) );
AO221x2_ASAP7_75t_L g1175 ( .A1(n_67), .A2(n_189), .B1(n_1132), .B2(n_1135), .C(n_1176), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g1410 ( .A1(n_68), .A2(n_126), .B1(n_535), .B2(n_537), .C(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g892 ( .A(n_69), .Y(n_892) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_70), .A2(n_160), .B1(n_478), .B2(n_604), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g1110 ( .A1(n_70), .A2(n_209), .B1(n_697), .B2(n_1028), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g1415 ( .A1(n_72), .A2(n_74), .B1(n_537), .B2(n_579), .C(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g651 ( .A(n_73), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g1399 ( .A1(n_74), .A2(n_224), .B1(n_609), .B2(n_614), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_75), .A2(n_179), .B1(n_518), .B2(n_522), .Y(n_1037) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_75), .A2(n_691), .B(n_1040), .C(n_1043), .Y(n_1039) );
INVx1_ASAP7_75t_L g594 ( .A(n_76), .Y(n_594) );
OAI222xp33_ASAP7_75t_L g643 ( .A1(n_76), .A2(n_112), .B1(n_644), .B2(n_645), .C1(n_652), .C2(n_657), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_77), .A2(n_360), .B(n_385), .C(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g439 ( .A(n_77), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g827 ( .A1(n_78), .A2(n_577), .B(n_744), .Y(n_827) );
OAI22xp5_ASAP7_75t_SL g856 ( .A1(n_79), .A2(n_92), .B1(n_284), .B2(n_305), .Y(n_856) );
OAI21xp33_ASAP7_75t_L g869 ( .A1(n_79), .A2(n_870), .B(n_873), .Y(n_869) );
INVx1_ASAP7_75t_L g464 ( .A(n_80), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_80), .A2(n_86), .B1(n_557), .B2(n_561), .C(n_565), .Y(n_556) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_81), .A2(n_83), .B1(n_499), .B2(n_780), .Y(n_809) );
INVx1_ASAP7_75t_L g819 ( .A(n_81), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_82), .A2(n_233), .B1(n_620), .B2(n_795), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_82), .A2(n_150), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g820 ( .A(n_83), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_84), .A2(n_240), .B1(n_1028), .B2(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_84), .A2(n_104), .B1(n_483), .B2(n_1063), .Y(n_1064) );
INVx1_ASAP7_75t_L g1350 ( .A(n_85), .Y(n_1350) );
INVx1_ASAP7_75t_L g455 ( .A(n_86), .Y(n_455) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_87), .Y(n_259) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_87), .B(n_257), .Y(n_1126) );
INVx1_ASAP7_75t_L g927 ( .A(n_88), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g950 ( .A1(n_88), .A2(n_190), .B1(n_606), .B2(n_951), .C(n_953), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_89), .A2(n_248), .B1(n_775), .B2(n_947), .Y(n_1083) );
AOI21xp33_ASAP7_75t_L g1107 ( .A1(n_89), .A2(n_579), .B(n_1108), .Y(n_1107) );
CKINVDCx5p33_ASAP7_75t_R g1392 ( .A(n_90), .Y(n_1392) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_91), .A2(n_846), .B(n_847), .C(n_849), .Y(n_845) );
INVxp33_ASAP7_75t_SL g874 ( .A(n_91), .Y(n_874) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_92), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_93), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_94), .Y(n_588) );
INVx1_ASAP7_75t_L g1010 ( .A(n_95), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_96), .A2(n_230), .B1(n_499), .B2(n_780), .Y(n_1094) );
INVx1_ASAP7_75t_L g1101 ( .A(n_96), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_97), .A2(n_206), .B1(n_976), .B2(n_979), .Y(n_975) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_97), .Y(n_982) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_98), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_98), .A2(n_182), .B1(n_778), .B2(n_955), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_99), .B(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1134 ( .A(n_99), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_100), .Y(n_1036) );
INVx1_ASAP7_75t_L g396 ( .A(n_101), .Y(n_396) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_101), .A2(n_289), .B(n_430), .C(n_435), .Y(n_429) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_102), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_102), .A2(n_227), .B1(n_772), .B2(n_773), .Y(n_771) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_103), .A2(n_561), .B(n_734), .C(n_745), .Y(n_733) );
INVx1_ASAP7_75t_L g765 ( .A(n_103), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_104), .A2(n_192), .B1(n_579), .B2(n_814), .C(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g998 ( .A(n_105), .Y(n_998) );
AOI21xp33_ASAP7_75t_L g1026 ( .A1(n_105), .A2(n_579), .B(n_859), .Y(n_1026) );
INVx2_ASAP7_75t_L g330 ( .A(n_106), .Y(n_330) );
INVx1_ASAP7_75t_L g369 ( .A(n_106), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_106), .B(n_331), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_107), .A2(n_187), .B1(n_1125), .B2(n_1129), .Y(n_1173) );
INVx1_ASAP7_75t_L g936 ( .A(n_108), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_109), .A2(n_128), .B1(n_905), .B2(n_906), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_109), .A2(n_175), .B1(n_614), .B2(n_955), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_111), .A2(n_200), .B1(n_522), .B2(n_994), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g1016 ( .A1(n_111), .A2(n_527), .B(n_1017), .C(n_1020), .Y(n_1016) );
INVx1_ASAP7_75t_L g592 ( .A(n_112), .Y(n_592) );
INVx1_ASAP7_75t_L g730 ( .A(n_113), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g779 ( .A1(n_113), .A2(n_242), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g1361 ( .A(n_115), .Y(n_1361) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_116), .A2(n_237), .B1(n_632), .B2(n_635), .C(n_637), .Y(n_631) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_117), .Y(n_735) );
INVx1_ASAP7_75t_L g283 ( .A(n_119), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_120), .A2(n_203), .B1(n_799), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g823 ( .A(n_120), .Y(n_823) );
INVx1_ASAP7_75t_L g323 ( .A(n_121), .Y(n_323) );
INVx1_ASAP7_75t_L g647 ( .A(n_123), .Y(n_647) );
INVxp67_ASAP7_75t_SL g1080 ( .A(n_124), .Y(n_1080) );
OAI211xp5_ASAP7_75t_L g1096 ( .A1(n_124), .A2(n_527), .B(n_1097), .C(n_1100), .Y(n_1096) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_125), .A2(n_223), .B1(n_775), .B2(n_947), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_125), .A2(n_248), .B1(n_546), .B2(n_829), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_127), .A2(n_1385), .B1(n_1421), .B2(n_1422), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1421 ( .A(n_127), .Y(n_1421) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_128), .A2(n_225), .B1(n_946), .B2(n_947), .Y(n_945) );
AO22x1_ASAP7_75t_L g1131 ( .A1(n_129), .A2(n_202), .B1(n_1132), .B2(n_1135), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_130), .A2(n_235), .B1(n_480), .B2(n_483), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_130), .A2(n_164), .B1(n_543), .B2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_131), .A2(n_153), .B1(n_474), .B2(n_770), .Y(n_769) );
BUFx3_ASAP7_75t_L g336 ( .A(n_132), .Y(n_336) );
INVx1_ASAP7_75t_L g1077 ( .A(n_133), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_133), .A2(n_134), .B1(n_658), .B2(n_756), .C(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1078 ( .A(n_134), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_135), .A2(n_209), .B1(n_478), .B2(n_617), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_135), .A2(n_160), .B1(n_535), .B2(n_541), .C(n_859), .Y(n_1098) );
INVx1_ASAP7_75t_L g1342 ( .A(n_136), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_137), .B(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g784 ( .A(n_139), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_140), .A2(n_151), .B1(n_1132), .B2(n_1135), .Y(n_1154) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_141), .A2(n_518), .B(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_142), .A2(n_150), .B1(n_618), .B2(n_795), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g813 ( .A1(n_142), .A2(n_233), .B1(n_541), .B2(n_754), .C(n_814), .Y(n_813) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_143), .Y(n_271) );
INVx1_ASAP7_75t_L g1407 ( .A(n_144), .Y(n_1407) );
INVx1_ASAP7_75t_L g1348 ( .A(n_145), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_146), .A2(n_175), .B1(n_906), .B2(n_923), .C(n_925), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_146), .A2(n_184), .B1(n_474), .B2(n_478), .C(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g1041 ( .A(n_147), .Y(n_1041) );
INVx1_ASAP7_75t_L g1314 ( .A(n_148), .Y(n_1314) );
OAI21xp5_ASAP7_75t_SL g1418 ( .A1(n_149), .A2(n_994), .B(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g553 ( .A(n_152), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_153), .A2(n_229), .B1(n_541), .B2(n_752), .C(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g626 ( .A(n_154), .Y(n_626) );
INVx1_ASAP7_75t_L g789 ( .A(n_155), .Y(n_789) );
OAI221xp5_ASAP7_75t_SL g821 ( .A1(n_155), .A2(n_231), .B1(n_557), .B2(n_657), .C(n_822), .Y(n_821) );
XOR2x2_ASAP7_75t_L g723 ( .A(n_156), .B(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_157), .A2(n_217), .B1(n_1125), .B2(n_1129), .Y(n_1139) );
INVx1_ASAP7_75t_L g597 ( .A(n_158), .Y(n_597) );
INVx1_ASAP7_75t_L g311 ( .A(n_159), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_161), .A2(n_177), .B1(n_401), .B2(n_404), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_161), .A2(n_177), .B1(n_413), .B2(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g287 ( .A(n_162), .Y(n_287) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_163), .A2(n_744), .B(n_859), .Y(n_866) );
INVx1_ASAP7_75t_L g882 ( .A(n_163), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_164), .A2(n_245), .B1(n_480), .B2(n_483), .Y(n_479) );
OAI211xp5_ASAP7_75t_SL g1310 ( .A1(n_165), .A2(n_385), .B(n_1311), .C(n_1313), .Y(n_1310) );
INVx1_ASAP7_75t_L g1331 ( .A(n_165), .Y(n_1331) );
INVxp67_ASAP7_75t_SL g1051 ( .A(n_166), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_166), .A2(n_191), .B1(n_490), .B2(n_770), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_167), .A2(n_212), .B1(n_1125), .B2(n_1129), .Y(n_1153) );
OAI22xp33_ASAP7_75t_L g1316 ( .A1(n_168), .A2(n_236), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_168), .A2(n_236), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_169), .Y(n_270) );
INVx1_ASAP7_75t_L g390 ( .A(n_170), .Y(n_390) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_171), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g760 ( .A(n_172), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_173), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_174), .A2(n_226), .B1(n_529), .B2(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g883 ( .A(n_174), .Y(n_883) );
INVx1_ASAP7_75t_L g302 ( .A(n_176), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_178), .B(n_1073), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_178), .A2(n_1090), .B1(n_1091), .B2(n_1111), .Y(n_1089) );
INVx1_ASAP7_75t_L g1113 ( .A(n_178), .Y(n_1113) );
AO22x1_ASAP7_75t_L g1169 ( .A1(n_180), .A2(n_204), .B1(n_1125), .B2(n_1170), .Y(n_1169) );
CKINVDCx16_ASAP7_75t_R g1177 ( .A(n_181), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1044 ( .A1(n_182), .A2(n_191), .B1(n_637), .B2(n_752), .C(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g699 ( .A(n_183), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_184), .A2(n_190), .B1(n_908), .B2(n_910), .C(n_911), .Y(n_907) );
INVx1_ASAP7_75t_L g312 ( .A(n_185), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_186), .A2(n_199), .B1(n_376), .B2(n_380), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_186), .A2(n_199), .B1(n_421), .B2(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g669 ( .A(n_188), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_192), .A2(n_240), .B1(n_483), .B2(n_1063), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g939 ( .A(n_193), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_193), .A2(n_195), .B1(n_968), .B2(n_970), .C(n_972), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_194), .A2(n_237), .B1(n_604), .B2(n_606), .Y(n_603) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_194), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_195), .A2(n_208), .B1(n_914), .B2(n_919), .C(n_920), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_196), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_197), .A2(n_222), .B1(n_1132), .B2(n_1135), .Y(n_1143) );
BUFx3_ASAP7_75t_L g274 ( .A(n_198), .Y(n_274) );
INVx1_ASAP7_75t_L g417 ( .A(n_198), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_201), .Y(n_1179) );
XOR2x2_ASAP7_75t_L g1303 ( .A(n_205), .B(n_1304), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_205), .A2(n_1383), .B1(n_1423), .B2(n_1425), .Y(n_1382) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_206), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_207), .A2(n_527), .B(n_532), .C(n_548), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_208), .A2(n_211), .B1(n_958), .B2(n_961), .Y(n_957) );
INVx1_ASAP7_75t_L g1355 ( .A(n_210), .Y(n_1355) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_211), .Y(n_941) );
INVx2_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
INVx1_ASAP7_75t_L g320 ( .A(n_213), .Y(n_320) );
INVx1_ASAP7_75t_L g368 ( .A(n_213), .Y(n_368) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_215), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_216), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g858 ( .A(n_218), .B(n_859), .Y(n_858) );
AO22x1_ASAP7_75t_L g1171 ( .A1(n_220), .A2(n_238), .B1(n_1132), .B2(n_1135), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_221), .Y(n_792) );
OAI211xp5_ASAP7_75t_SL g811 ( .A1(n_221), .A2(n_691), .B(n_812), .C(n_818), .Y(n_811) );
INVx1_ASAP7_75t_L g1105 ( .A(n_223), .Y(n_1105) );
INVx1_ASAP7_75t_L g926 ( .A(n_225), .Y(n_926) );
INVxp67_ASAP7_75t_SL g888 ( .A(n_226), .Y(n_888) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_227), .A2(n_743), .B(n_744), .Y(n_742) );
OAI22xp33_ASAP7_75t_SL g1012 ( .A1(n_228), .A2(n_239), .B1(n_457), .B2(n_1013), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1023 ( .A1(n_228), .A2(n_239), .B1(n_557), .B2(n_658), .C(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1102 ( .A(n_230), .Y(n_1102) );
INVx1_ASAP7_75t_L g790 ( .A(n_231), .Y(n_790) );
XNOR2xp5_ASAP7_75t_L g989 ( .A(n_232), .B(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g662 ( .A(n_234), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g573 ( .A1(n_235), .A2(n_245), .B1(n_574), .B2(n_575), .C(n_579), .Y(n_573) );
INVx1_ASAP7_75t_L g1315 ( .A(n_241), .Y(n_1315) );
OAI211xp5_ASAP7_75t_L g1322 ( .A1(n_241), .A2(n_1323), .B(n_1326), .C(n_1327), .Y(n_1322) );
INVx1_ASAP7_75t_L g728 ( .A(n_242), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_243), .Y(n_850) );
INVx1_ASAP7_75t_L g1358 ( .A(n_244), .Y(n_1358) );
INVx1_ASAP7_75t_L g865 ( .A(n_246), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_275), .B(n_1116), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_260), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_254), .B(n_263), .Y(n_1381) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_256), .B(n_259), .Y(n_1424) );
INVx1_ASAP7_75t_L g1426 ( .A(n_256), .Y(n_1426) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_259), .B(n_1426), .Y(n_1429) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g446 ( .A(n_263), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g321 ( .A(n_264), .B(n_274), .Y(n_321) );
AND2x4_ASAP7_75t_L g580 ( .A(n_264), .B(n_273), .Y(n_580) );
INVx1_ASAP7_75t_L g413 ( .A(n_265), .Y(n_413) );
AND2x4_ASAP7_75t_SL g1380 ( .A(n_265), .B(n_1381), .Y(n_1380) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x6_ASAP7_75t_L g266 ( .A(n_267), .B(n_272), .Y(n_266) );
OR2x6_ASAP7_75t_L g422 ( .A(n_267), .B(n_416), .Y(n_422) );
INVxp67_ASAP7_75t_L g710 ( .A(n_267), .Y(n_710) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_268), .Y(n_568) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g286 ( .A(n_270), .Y(n_286) );
NAND2x1_ASAP7_75t_L g291 ( .A(n_270), .B(n_271), .Y(n_291) );
INVx2_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
AND2x2_ASAP7_75t_L g418 ( .A(n_270), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g434 ( .A(n_270), .B(n_271), .Y(n_434) );
INVx1_ASAP7_75t_L g444 ( .A(n_270), .Y(n_444) );
OR2x2_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_271), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g419 ( .A(n_271), .Y(n_419) );
BUFx2_ASAP7_75t_L g438 ( .A(n_271), .Y(n_438) );
INVx1_ASAP7_75t_L g515 ( .A(n_271), .Y(n_515) );
AND2x2_ASAP7_75t_L g530 ( .A(n_271), .B(n_309), .Y(n_530) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g432 ( .A(n_273), .Y(n_432) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx2_ASAP7_75t_L g428 ( .A(n_274), .Y(n_428) );
AND2x4_ASAP7_75t_L g442 ( .A(n_274), .B(n_443), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_719), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_583), .B1(n_584), .B2(n_718), .Y(n_276) );
INVx1_ASAP7_75t_L g718 ( .A(n_277), .Y(n_718) );
OA22x2_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_449), .B1(n_450), .B2(n_582), .Y(n_277) );
INVx1_ASAP7_75t_L g582 ( .A(n_278), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_374), .C(n_411), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_325), .Y(n_280) );
OAI33xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_292), .A3(n_297), .B1(n_310), .B2(n_313), .B3(n_322), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_287), .B2(n_288), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_283), .A2(n_311), .B1(n_348), .B2(n_353), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_284), .A2(n_303), .B1(n_323), .B2(n_324), .Y(n_322) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g650 ( .A(n_285), .Y(n_650) );
BUFx3_ASAP7_75t_L g909 ( .A(n_285), .Y(n_909) );
INVx2_ASAP7_75t_L g1372 ( .A(n_285), .Y(n_1372) );
AND2x2_ASAP7_75t_L g514 ( .A(n_286), .B(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_286), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_287), .A2(n_312), .B1(n_358), .B2(n_360), .Y(n_357) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_289), .A2(n_299), .B1(n_311), .B2(n_312), .Y(n_310) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx4f_ASAP7_75t_L g646 ( .A(n_290), .Y(n_646) );
BUFx4f_ASAP7_75t_L g736 ( .A(n_290), .Y(n_736) );
INVx4_ASAP7_75t_L g848 ( .A(n_290), .Y(n_848) );
OR2x6_ASAP7_75t_L g920 ( .A(n_290), .B(n_921), .Y(n_920) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g826 ( .A(n_291), .Y(n_826) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_293), .A2(n_646), .B1(n_909), .B2(n_926), .C(n_927), .Y(n_925) );
INVx2_ASAP7_75t_L g1363 ( .A(n_293), .Y(n_1363) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g661 ( .A(n_294), .Y(n_661) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_294), .B(n_949), .Y(n_1398) );
BUFx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g472 ( .A(n_295), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_295), .B(n_513), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_302), .B2(n_303), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_298), .A2(n_323), .B1(n_333), .B2(n_339), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_299), .A2(n_1051), .B1(n_1052), .B2(n_1053), .C(n_1054), .Y(n_1050) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_301), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_302), .A2(n_324), .B1(n_371), .B2(n_373), .Y(n_370) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g571 ( .A(n_306), .Y(n_571) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_306), .Y(n_656) );
INVx2_ASAP7_75t_SL g749 ( .A(n_306), .Y(n_749) );
INVx8_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g924 ( .A(n_307), .Y(n_924) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1375 ( .A(n_316), .B(n_321), .Y(n_1375) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_318), .Y(n_410) );
OR2x2_ASAP7_75t_L g497 ( .A(n_318), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_SL g912 ( .A(n_318), .B(n_321), .Y(n_912) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g448 ( .A(n_319), .Y(n_448) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g541 ( .A(n_321), .Y(n_541) );
INVx1_ASAP7_75t_SL g637 ( .A(n_321), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_321), .B(n_858), .C(n_860), .D(n_862), .Y(n_857) );
INVx4_ASAP7_75t_L g1411 ( .A(n_321), .Y(n_1411) );
OAI33xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_332), .A3(n_347), .B1(n_357), .B2(n_362), .B3(n_370), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_SL g996 ( .A1(n_327), .A2(n_997), .B1(n_1005), .B2(n_1006), .Y(n_996) );
BUFx4f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g879 ( .A(n_328), .Y(n_879) );
BUFx2_ASAP7_75t_L g953 ( .A(n_329), .Y(n_953) );
NAND2xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_330), .Y(n_408) );
INVx1_ASAP7_75t_L g463 ( .A(n_330), .Y(n_463) );
AND3x4_ASAP7_75t_L g471 ( .A(n_330), .B(n_394), .C(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
BUFx3_ASAP7_75t_L g394 ( .A(n_331), .Y(n_394) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
BUFx4f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x4_ASAP7_75t_L g378 ( .A(n_335), .B(n_379), .Y(n_378) );
OR2x4_ASAP7_75t_L g403 ( .A(n_335), .B(n_366), .Y(n_403) );
INVx2_ASAP7_75t_L g494 ( .A(n_335), .Y(n_494) );
BUFx3_ASAP7_75t_L g1343 ( .A(n_335), .Y(n_1343) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_336), .Y(n_346) );
INVx2_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_336), .B(n_345), .Y(n_356) );
AND2x4_ASAP7_75t_L g387 ( .A(n_336), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g477 ( .A(n_337), .Y(n_477) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_L g351 ( .A(n_338), .Y(n_351) );
INVx2_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g521 ( .A(n_342), .B(n_497), .Y(n_521) );
INVx4_ASAP7_75t_L g1312 ( .A(n_342), .Y(n_1312) );
INVx3_ASAP7_75t_L g1346 ( .A(n_342), .Y(n_1346) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx3_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
BUFx2_ASAP7_75t_L g973 ( .A(n_343), .Y(n_973) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
BUFx2_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g388 ( .A(n_345), .Y(n_388) );
BUFx2_ASAP7_75t_L g395 ( .A(n_346), .Y(n_395) );
INVx2_ASAP7_75t_L g459 ( .A(n_346), .Y(n_459) );
AND2x4_ASAP7_75t_L g484 ( .A(n_346), .B(n_469), .Y(n_484) );
INVx1_ASAP7_75t_L g1063 ( .A(n_348), .Y(n_1063) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
AND2x4_ASAP7_75t_L g405 ( .A(n_349), .B(n_379), .Y(n_405) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_349), .Y(n_609) );
INVx2_ASAP7_75t_L g1007 ( .A(n_349), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx8_ASAP7_75t_L g482 ( .A(n_350), .Y(n_482) );
INVx2_ASAP7_75t_L g677 ( .A(n_350), .Y(n_677) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_350), .Y(n_682) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g476 ( .A(n_352), .B(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g373 ( .A(n_354), .Y(n_373) );
CKINVDCx8_ASAP7_75t_R g1009 ( .A(n_354), .Y(n_1009) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g510 ( .A(n_355), .Y(n_510) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g383 ( .A(n_356), .Y(n_383) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI33xp33_ASAP7_75t_L g1060 ( .A1(n_363), .A2(n_471), .A3(n_1061), .B1(n_1062), .B2(n_1064), .B3(n_1065), .Y(n_1060) );
BUFx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g486 ( .A(n_364), .Y(n_486) );
BUFx2_ASAP7_75t_L g615 ( .A(n_364), .Y(n_615) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_364), .Y(n_1086) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g803 ( .A(n_365), .Y(n_803) );
NAND3x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .C(n_369), .Y(n_365) );
INVx1_ASAP7_75t_L g379 ( .A(n_366), .Y(n_379) );
OR2x6_ASAP7_75t_L g382 ( .A(n_366), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g386 ( .A(n_366), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g462 ( .A(n_366), .B(n_463), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g949 ( .A(n_366), .B(n_369), .Y(n_949) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g461 ( .A(n_368), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_368), .B(n_531), .Y(n_935) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_373), .A2(n_881), .B1(n_882), .B2(n_883), .C(n_884), .Y(n_880) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_384), .A3(n_400), .B(n_406), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g1317 ( .A(n_378), .Y(n_1317) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g1319 ( .A(n_382), .Y(n_1319) );
INVx1_ASAP7_75t_L g1001 ( .A(n_383), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_383), .Y(n_1354) );
CKINVDCx8_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g478 ( .A(n_387), .Y(n_478) );
BUFx2_ASAP7_75t_L g505 ( .A(n_387), .Y(n_505) );
INVx2_ASAP7_75t_L g607 ( .A(n_387), .Y(n_607) );
BUFx2_ASAP7_75t_L g620 ( .A(n_387), .Y(n_620) );
BUFx2_ASAP7_75t_L g770 ( .A(n_387), .Y(n_770) );
AND2x2_ASAP7_75t_L g962 ( .A(n_387), .B(n_960), .Y(n_962) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_387), .Y(n_1004) );
INVx1_ASAP7_75t_L g469 ( .A(n_388), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_396), .B2(n_397), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_390), .A2(n_436), .B1(n_439), .B2(n_440), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_391), .A2(n_397), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
BUFx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
AND2x4_ASAP7_75t_L g398 ( .A(n_393), .B(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g1308 ( .A(n_403), .Y(n_1308) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g1309 ( .A(n_405), .Y(n_1309) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_406), .Y(n_1320) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI31xp33_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_420), .A3(n_429), .B(n_445), .Y(n_411) );
INVx3_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g1338 ( .A(n_415), .Y(n_1338) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_418), .Y(n_539) );
INVx2_ASAP7_75t_L g578 ( .A(n_418), .Y(n_578) );
BUFx3_ASAP7_75t_L g859 ( .A(n_418), .Y(n_859) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g1333 ( .A(n_422), .Y(n_1333) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g1336 ( .A(n_427), .Y(n_1336) );
AND2x4_ASAP7_75t_L g437 ( .A(n_428), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_428), .B(n_438), .Y(n_1328) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g1326 ( .A(n_431), .Y(n_1326) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_433), .Y(n_535) );
AND2x6_ASAP7_75t_L g547 ( .A(n_433), .B(n_513), .Y(n_547) );
AND2x4_ASAP7_75t_SL g560 ( .A(n_433), .B(n_531), .Y(n_560) );
BUFx3_ASAP7_75t_L g574 ( .A(n_433), .Y(n_574) );
BUFx3_ASAP7_75t_L g754 ( .A(n_433), .Y(n_754) );
BUFx3_ASAP7_75t_L g863 ( .A(n_433), .Y(n_863) );
INVx1_ASAP7_75t_L g1046 ( .A(n_433), .Y(n_1046) );
BUFx3_ASAP7_75t_L g1416 ( .A(n_433), .Y(n_1416) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g634 ( .A(n_434), .Y(n_634) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g563 ( .A(n_438), .Y(n_563) );
BUFx2_ASAP7_75t_L g851 ( .A(n_438), .Y(n_851) );
INVx1_ASAP7_75t_L g918 ( .A(n_438), .Y(n_918) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g1330 ( .A(n_442), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_443), .B(n_513), .Y(n_520) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI31xp33_ASAP7_75t_L g1321 ( .A1(n_445), .A2(n_1322), .A3(n_1332), .B(n_1337), .Y(n_1321) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g519 ( .A(n_448), .B(n_520), .Y(n_519) );
INVxp67_ASAP7_75t_L g524 ( .A(n_448), .Y(n_524) );
INVx1_ASAP7_75t_L g896 ( .A(n_448), .Y(n_896) );
OR2x2_ASAP7_75t_L g919 ( .A(n_448), .B(n_520), .Y(n_919) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_506), .C(n_525), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_491), .C(n_502), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_470), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_464), .B2(n_465), .Y(n_454) );
AOI221x1_ASAP7_75t_L g877 ( .A1(n_456), .A2(n_465), .B1(n_841), .B2(n_850), .C(n_878), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_456), .A2(n_465), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g593 ( .A(n_458), .B(n_460), .Y(n_593) );
AND2x2_ASAP7_75t_L g766 ( .A(n_458), .B(n_460), .Y(n_766) );
AND2x6_ASAP7_75t_L g969 ( .A(n_458), .B(n_462), .Y(n_969) );
AND2x4_ASAP7_75t_SL g1393 ( .A(n_458), .B(n_460), .Y(n_1393) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g465 ( .A(n_460), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g504 ( .A(n_460), .B(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_SL g1014 ( .A(n_460), .B(n_466), .Y(n_1014) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OR2x2_ASAP7_75t_L g511 ( .A(n_461), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g930 ( .A(n_461), .Y(n_930) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_462), .B(n_476), .Y(n_523) );
AND2x2_ASAP7_75t_L g971 ( .A(n_462), .B(n_468), .Y(n_971) );
INVx1_ASAP7_75t_L g974 ( .A(n_462), .Y(n_974) );
AO22x1_ASAP7_75t_L g591 ( .A1(n_465), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_465), .A2(n_593), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_465), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_465), .A2(n_766), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_465), .A2(n_766), .B1(n_1067), .B2(n_1068), .Y(n_1066) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI33xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .A3(n_479), .B1(n_485), .B2(n_486), .B3(n_487), .Y(n_470) );
BUFx3_ASAP7_75t_L g602 ( .A(n_471), .Y(n_602) );
AOI33xp33_ASAP7_75t_L g768 ( .A1(n_471), .A2(n_486), .A3(n_769), .B1(n_771), .B2(n_774), .B3(n_777), .Y(n_768) );
AOI33xp33_ASAP7_75t_L g1081 ( .A1(n_471), .A2(n_1082), .A3(n_1083), .B1(n_1084), .B2(n_1085), .B3(n_1086), .Y(n_1081) );
INVx1_ASAP7_75t_L g1401 ( .A(n_471), .Y(n_1401) );
INVx2_ASAP7_75t_SL g581 ( .A(n_472), .Y(n_581) );
INVx1_ASAP7_75t_L g715 ( .A(n_472), .Y(n_715) );
BUFx2_ASAP7_75t_L g795 ( .A(n_474), .Y(n_795) );
INVx8_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g617 ( .A(n_475), .Y(n_617) );
INVx2_ASAP7_75t_L g625 ( .A(n_475), .Y(n_625) );
INVx2_ASAP7_75t_L g1397 ( .A(n_475), .Y(n_1397) );
INVx8_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g490 ( .A(n_476), .Y(n_490) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_476), .Y(n_890) );
BUFx3_ASAP7_75t_L g956 ( .A(n_476), .Y(n_956) );
AND2x2_ASAP7_75t_L g959 ( .A(n_476), .B(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g500 ( .A(n_482), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g802 ( .A(n_482), .Y(n_802) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx5_ASAP7_75t_L g611 ( .A(n_484), .Y(n_611) );
BUFx12f_ASAP7_75t_L g614 ( .A(n_484), .Y(n_614) );
BUFx3_ASAP7_75t_L g678 ( .A(n_484), .Y(n_678) );
BUFx2_ASAP7_75t_L g947 ( .A(n_484), .Y(n_947) );
AND2x4_ASAP7_75t_L g980 ( .A(n_484), .B(n_978), .Y(n_980) );
AOI33xp33_ASAP7_75t_L g671 ( .A1(n_486), .A2(n_602), .A3(n_672), .B1(n_674), .B2(n_679), .B3(n_683), .Y(n_671) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g605 ( .A(n_490), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_492), .B(n_894), .Y(n_893) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
OR2x2_ASAP7_75t_L g780 ( .A(n_493), .B(n_495), .Y(n_780) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g871 ( .A(n_496), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g501 ( .A(n_497), .Y(n_501) );
OR2x2_ASAP7_75t_L g509 ( .A(n_497), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g960 ( .A(n_498), .Y(n_960) );
INVx1_ASAP7_75t_L g978 ( .A(n_498), .Y(n_978) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_500), .A2(n_623), .B1(n_624), .B2(n_626), .Y(n_622) );
INVx2_ASAP7_75t_L g781 ( .A(n_500), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_500), .A2(n_624), .B1(n_1021), .B2(n_1022), .Y(n_1029) );
AND2x4_ASAP7_75t_L g624 ( .A(n_501), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_501), .B(n_625), .Y(n_1420) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND5x1_ASAP7_75t_L g837 ( .A(n_503), .B(n_838), .C(n_877), .D(n_891), .E(n_897), .Y(n_837) );
AND4x1_ASAP7_75t_L g1057 ( .A(n_503), .B(n_1058), .C(n_1060), .D(n_1066), .Y(n_1057) );
NAND3xp33_ASAP7_75t_SL g1390 ( .A(n_503), .B(n_1391), .C(n_1395), .Y(n_1390) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g600 ( .A(n_504), .Y(n_600) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_504), .Y(n_685) );
BUFx2_ASAP7_75t_L g673 ( .A(n_505), .Y(n_673) );
AOI21xp33_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_516), .B(n_517), .Y(n_506) );
AOI211x1_ASAP7_75t_L g587 ( .A1(n_507), .A2(n_588), .B(n_589), .C(n_621), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_507), .A2(n_687), .B(n_688), .Y(n_686) );
AOI21xp33_ASAP7_75t_SL g759 ( .A1(n_507), .A2(n_760), .B(n_761), .Y(n_759) );
AOI211x1_ASAP7_75t_L g785 ( .A1(n_507), .A2(n_786), .B(n_787), .C(n_805), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g991 ( .A1(n_507), .A2(n_992), .B(n_993), .Y(n_991) );
AOI21xp33_ASAP7_75t_L g1035 ( .A1(n_507), .A2(n_1036), .B(n_1037), .Y(n_1035) );
NAND2xp33_ASAP7_75t_L g1087 ( .A(n_507), .B(n_1088), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1386 ( .A1(n_507), .A2(n_1387), .B1(n_1388), .B2(n_1389), .C(n_1390), .Y(n_1386) );
INVx8_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g875 ( .A(n_509), .Y(n_875) );
BUFx3_ASAP7_75t_L g887 ( .A(n_510), .Y(n_887) );
INVx1_ASAP7_75t_L g931 ( .A(n_512), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g564 ( .A(n_513), .Y(n_564) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_513), .B(n_851), .Y(n_1417) );
INVx3_ASAP7_75t_L g544 ( .A(n_514), .Y(n_544) );
AND2x2_ASAP7_75t_L g552 ( .A(n_514), .B(n_531), .Y(n_552) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_514), .Y(n_740) );
INVx2_ASAP7_75t_L g807 ( .A(n_518), .Y(n_807) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
AND2x4_ASAP7_75t_L g994 ( .A(n_519), .B(n_521), .Y(n_994) );
INVx2_ASAP7_75t_L g876 ( .A(n_521), .Y(n_876) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
OR2x6_ASAP7_75t_L g599 ( .A(n_523), .B(n_524), .Y(n_599) );
INVx2_ASAP7_75t_L g966 ( .A(n_523), .Y(n_966) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_556), .B(n_581), .Y(n_525) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_R g642 ( .A(n_528), .B(n_597), .Y(n_642) );
INVx3_ASAP7_75t_L g691 ( .A(n_528), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_528), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
BUFx2_ASAP7_75t_L g741 ( .A(n_529), .Y(n_741) );
INVx1_ASAP7_75t_L g831 ( .A(n_529), .Y(n_831) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g546 ( .A(n_530), .Y(n_546) );
INVx2_ASAP7_75t_L g817 ( .A(n_530), .Y(n_817) );
AND2x4_ASAP7_75t_L g555 ( .A(n_531), .B(n_539), .Y(n_555) );
BUFx2_ASAP7_75t_L g855 ( .A(n_531), .Y(n_855) );
AND2x2_ASAP7_75t_L g984 ( .A(n_531), .B(n_539), .Y(n_984) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_531), .B(n_816), .Y(n_1409) );
AOI21xp5_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_542), .B(n_547), .Y(n_532) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g695 ( .A(n_537), .Y(n_695) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_539), .Y(n_636) );
HB1xp67_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g639 ( .A(n_544), .Y(n_639) );
INVx2_ASAP7_75t_L g697 ( .A(n_544), .Y(n_697) );
INVx1_ASAP7_75t_L g861 ( .A(n_544), .Y(n_861) );
INVx2_ASAP7_75t_L g1048 ( .A(n_544), .Y(n_1048) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_SL g641 ( .A(n_546), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_547), .A2(n_631), .B(n_638), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_547), .A2(n_693), .B(n_696), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_547), .A2(n_554), .B(n_728), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_547), .A2(n_813), .B(n_815), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_547), .A2(n_1018), .B(n_1019), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1043 ( .A1(n_547), .A2(n_1044), .B(n_1047), .Y(n_1043) );
AOI21xp5_ASAP7_75t_L g1097 ( .A1(n_547), .A2(n_1098), .B(n_1099), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_547), .A2(n_1388), .B1(n_1409), .B2(n_1410), .C(n_1412), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_553), .B2(n_554), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_550), .A2(n_555), .B1(n_623), .B2(n_626), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_550), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_552), .Y(n_731) );
AND2x4_ASAP7_75t_L g895 ( .A(n_552), .B(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_554), .A2(n_731), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_554), .A2(n_731), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g702 ( .A(n_555), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_555), .A2(n_731), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_555), .A2(n_731), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_555), .A2(n_731), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g644 ( .A(n_558), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_558), .A2(n_562), .B1(n_669), .B2(n_670), .Y(n_711) );
INVx2_ASAP7_75t_L g756 ( .A(n_558), .Y(n_756) );
INVx4_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g842 ( .A(n_560), .Y(n_842) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g658 ( .A(n_562), .Y(n_658) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g844 ( .A(n_564), .Y(n_844) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_572), .C(n_573), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_566), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx4_ASAP7_75t_L g846 ( .A(n_568), .Y(n_846) );
INVx3_ASAP7_75t_L g1367 ( .A(n_568), .Y(n_1367) );
INVx1_ASAP7_75t_L g905 ( .A(n_570), .Y(n_905) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_570), .Y(n_1052) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g743 ( .A(n_576), .Y(n_743) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_577), .Y(n_707) );
INVx1_ASAP7_75t_L g753 ( .A(n_577), .Y(n_753) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g814 ( .A(n_578), .Y(n_814) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_580), .A2(n_646), .B1(n_647), .B2(n_648), .C(n_651), .Y(n_645) );
INVx2_ASAP7_75t_L g708 ( .A(n_580), .Y(n_708) );
INVx3_ASAP7_75t_L g744 ( .A(n_580), .Y(n_744) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_663), .B1(n_716), .B2(n_717), .Y(n_584) );
INVx2_ASAP7_75t_L g717 ( .A(n_585), .Y(n_717) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_662), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_627), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_601), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_595), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_600), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_598), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_598), .B(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_598), .B(n_1080), .Y(n_1079) );
INVx5_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx3_ASAP7_75t_L g1387 ( .A(n_599), .Y(n_1387) );
INVx1_ASAP7_75t_L g782 ( .A(n_600), .Y(n_782) );
NAND4xp25_ASAP7_75t_SL g787 ( .A(n_600), .B(n_788), .C(n_791), .D(n_793), .Y(n_787) );
NAND4xp25_ASAP7_75t_SL g1075 ( .A(n_600), .B(n_1076), .C(n_1079), .D(n_1081), .Y(n_1075) );
AOI33xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .A3(n_608), .B1(n_612), .B2(n_615), .B3(n_616), .Y(n_601) );
AOI33xp33_ASAP7_75t_L g793 ( .A1(n_602), .A2(n_794), .A3(n_796), .B1(n_800), .B2(n_803), .B3(n_804), .Y(n_793) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g778 ( .A(n_607), .Y(n_778) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_R g773 ( .A(n_611), .Y(n_773) );
INVx1_ASAP7_75t_L g799 ( .A(n_611), .Y(n_799) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_643), .B(n_659), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_629), .B(n_630), .C(n_642), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g706 ( .A(n_633), .Y(n_706) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_SL g910 ( .A(n_646), .Y(n_910) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx4_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx5_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx6_ASAP7_75t_L g1368 ( .A(n_656), .Y(n_1368) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_659), .A2(n_1016), .B(n_1023), .Y(n_1015) );
OAI21xp5_ASAP7_75t_L g1095 ( .A1(n_659), .A2(n_1096), .B(n_1103), .Y(n_1095) );
AOI21xp5_ASAP7_75t_L g1403 ( .A1(n_659), .A2(n_1404), .B(n_1418), .Y(n_1403) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g832 ( .A(n_660), .Y(n_832) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g1056 ( .A(n_661), .Y(n_1056) );
INVx1_ASAP7_75t_L g716 ( .A(n_663), .Y(n_716) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_686), .C(n_689), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_684), .C(n_685), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g798 ( .A(n_677), .Y(n_798) );
INVx3_ASAP7_75t_L g872 ( .A(n_677), .Y(n_872) );
INVx1_ASAP7_75t_L g946 ( .A(n_677), .Y(n_946) );
OR2x6_ASAP7_75t_SL g976 ( .A(n_677), .B(n_977), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_677), .A2(n_998), .B1(n_999), .B2(n_1002), .C(n_1003), .Y(n_997) );
INVx8_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g886 ( .A1(n_681), .A2(n_865), .B1(n_887), .B2(n_888), .C(n_889), .Y(n_886) );
BUFx3_ASAP7_75t_L g1349 ( .A(n_681), .Y(n_1349) );
INVx5_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_682), .Y(n_772) );
INVx2_ASAP7_75t_SL g776 ( .A(n_682), .Y(n_776) );
INVx2_ASAP7_75t_SL g881 ( .A(n_682), .Y(n_881) );
INVx3_ASAP7_75t_L g952 ( .A(n_682), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g995 ( .A(n_685), .B(n_996), .C(n_1012), .Y(n_995) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_703), .B(n_712), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_709), .Y(n_704) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g758 ( .A(n_714), .Y(n_758) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_714), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_714), .A2(n_944), .B(n_963), .C(n_981), .Y(n_943) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_1030), .B2(n_1115), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_833), .Y(n_721) );
XNOR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_783), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_759), .C(n_762), .Y(n_724) );
OAI31xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_733), .A3(n_755), .B(n_757), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
OAI211xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_737), .C(n_742), .Y(n_734) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_740), .Y(n_829) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_748), .B2(n_750), .C(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g906 ( .A(n_746), .Y(n_906) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_779), .C(n_782), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_768), .Y(n_763) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
XNOR2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g885 ( .A(n_803), .Y(n_885) );
INVx2_ASAP7_75t_L g1005 ( .A(n_803), .Y(n_1005) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_803), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B(n_809), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g1092 ( .A1(n_807), .A2(n_1093), .B(n_1094), .Y(n_1092) );
OAI21xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_821), .B(n_832), .Y(n_810) );
AND2x4_ASAP7_75t_L g933 ( .A(n_816), .B(n_934), .Y(n_933) );
INVx3_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g1028 ( .A(n_817), .Y(n_1028) );
OAI211xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B(n_827), .C(n_828), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g864 ( .A1(n_824), .A2(n_865), .B(n_866), .C(n_867), .Y(n_864) );
INVx5_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
OR2x2_ASAP7_75t_L g938 ( .A(n_826), .B(n_935), .Y(n_938) );
BUFx3_ASAP7_75t_L g1325 ( .A(n_826), .Y(n_1325) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_987), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B1(n_899), .B2(n_986), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_868), .B(n_869), .Y(n_838) );
NAND4xp25_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .C(n_857), .D(n_864), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
AOI222xp33_ASAP7_75t_L g1413 ( .A1(n_842), .A2(n_1392), .B1(n_1394), .B2(n_1414), .C1(n_1415), .C2(n_1417), .Y(n_1413) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_855), .B2(n_856), .Y(n_843) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g1025 ( .A(n_848), .Y(n_1025) );
INVx2_ASAP7_75t_L g1106 ( .A(n_848), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_852), .B2(n_853), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_852), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1109 ( .A(n_859), .Y(n_1109) );
INVx2_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_871), .A2(n_1406), .B1(n_1407), .B2(n_1420), .Y(n_1419) );
OAI22xp5_ASAP7_75t_SL g878 ( .A1(n_879), .A2(n_880), .B1(n_885), .B2(n_886), .Y(n_878) );
OAI33xp33_ASAP7_75t_L g1340 ( .A1(n_879), .A2(n_1341), .A3(n_1347), .B1(n_1351), .B2(n_1356), .B3(n_1357), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g942 ( .A(n_894), .Y(n_942) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AND2x4_ASAP7_75t_L g983 ( .A(n_896), .B(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g986 ( .A(n_899), .Y(n_986) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
XNOR2x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_985), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_943), .Y(n_901) );
NAND3xp33_ASAP7_75t_SL g902 ( .A(n_903), .B(n_928), .C(n_940), .Y(n_902) );
AOI211xp5_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_907), .B(n_913), .C(n_922), .Y(n_903) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_917), .Y(n_914) );
INVx1_ASAP7_75t_L g921 ( .A(n_915), .Y(n_921) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI222xp33_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_932), .B1(n_933), .B2(n_936), .C1(n_937), .C2(n_939), .Y(n_928) );
AND2x4_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AOI211xp5_ASAP7_75t_L g963 ( .A1(n_936), .A2(n_964), .B(n_967), .C(n_975), .Y(n_963) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_948), .B1(n_950), .B2(n_954), .C(n_957), .Y(n_944) );
INVx2_ASAP7_75t_L g1352 ( .A(n_951), .Y(n_1352) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
BUFx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx4_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OR2x6_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .Y(n_972) );
INVx1_ASAP7_75t_L g1360 ( .A(n_973), .Y(n_1360) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx3_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
AND4x1_ASAP7_75t_L g990 ( .A(n_991), .B(n_995), .C(n_1015), .D(n_1029), .Y(n_990) );
INVx3_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1006) );
OAI211xp5_ASAP7_75t_L g1024 ( .A1(n_1008), .A2(n_1025), .B(n_1026), .C(n_1027), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1009), .A2(n_1348), .B1(n_1349), .B2(n_1350), .Y(n_1347) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1391 ( .A1(n_1014), .A2(n_1392), .B1(n_1393), .B2(n_1394), .Y(n_1391) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_1025), .A2(n_1344), .B1(n_1361), .B2(n_1370), .Y(n_1373) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1030), .Y(n_1115) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
OAI22x1_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1070), .B1(n_1071), .B2(n_1114), .Y(n_1031) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1032), .Y(n_1114) );
AO21x2_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .B(n_1069), .Y(n_1032) );
NAND3xp33_ASAP7_75t_SL g1034 ( .A(n_1035), .B(n_1038), .C(n_1057), .Y(n_1034) );
OAI21xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1049), .B(n_1056), .Y(n_1038) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1046), .Y(n_1055) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NAND2x1p5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1089), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1087), .Y(n_1073) );
INVxp67_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
NOR2xp33_ASAP7_75t_SL g1111 ( .A(n_1075), .B(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1087), .B(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1095), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B(n_1107), .C(n_1110), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_1106), .A2(n_1348), .B1(n_1353), .B2(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1300), .B1(n_1302), .B2(n_1377), .C(n_1382), .Y(n_1116) );
AOI221xp5_ASAP7_75t_SL g1117 ( .A1(n_1118), .A2(n_1181), .B1(n_1238), .B2(n_1240), .C(n_1267), .Y(n_1117) );
A2O1A1Ixp33_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1155), .B(n_1166), .C(n_1175), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1150), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1140), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1122), .B(n_1147), .Y(n_1192) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1122), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1122), .B(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1137), .Y(n_1122) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1123), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1123), .B(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1123), .B(n_1160), .Y(n_1189) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1131), .Y(n_1123) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1125), .Y(n_1178) );
AND2x6_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1126), .B(n_1130), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_1126), .B(n_1133), .Y(n_1132) );
AND2x6_ASAP7_75t_L g1135 ( .A(n_1126), .B(n_1136), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1126), .B(n_1130), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1126), .B(n_1130), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1126), .B(n_1133), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1128), .B(n_1134), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1180 ( .A(n_1129), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1427 ( .A(n_1133), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1137), .B(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1137), .Y(n_1165) );
AND3x1_ASAP7_75t_L g1210 ( .A(n_1137), .B(n_1141), .C(n_1162), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1137), .B(n_1160), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1137), .B(n_1141), .Y(n_1219) );
OAI32xp33_ASAP7_75t_L g1296 ( .A1(n_1137), .A2(n_1211), .A3(n_1221), .B1(n_1297), .B2(n_1299), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1140), .B(n_1226), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1140), .B(n_1161), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1146), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1141), .B(n_1164), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1141), .B(n_1233), .Y(n_1279) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_1142), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1142), .B(n_1164), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1142), .B(n_1192), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1142), .B(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1142), .B(n_1226), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1146), .B(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1146), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1146), .B(n_1212), .Y(n_1211) );
NOR2xp33_ASAP7_75t_L g1214 ( .A(n_1146), .B(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1146), .B(n_1207), .Y(n_1266) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1147), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1147), .B(n_1152), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1147), .B(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1147), .B(n_1172), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1147), .B(n_1152), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1147), .B(n_1189), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1147), .B(n_1160), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1147), .B(n_1218), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1147), .B(n_1168), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
INVx2_ASAP7_75t_L g1183 ( .A(n_1150), .Y(n_1183) );
A2O1A1Ixp33_ASAP7_75t_L g1186 ( .A1(n_1150), .A2(n_1187), .B(n_1188), .C(n_1190), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1150), .B(n_1201), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1150), .B(n_1284), .Y(n_1283) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1151), .B(n_1172), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1151), .B(n_1201), .Y(n_1274) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1152), .B(n_1172), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1152), .B(n_1208), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1152), .B(n_1172), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1154), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1157), .B1(n_1159), .B2(n_1163), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1157), .B(n_1185), .Y(n_1184) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1158), .B(n_1226), .Y(n_1233) );
O2A1O1Ixp33_ASAP7_75t_SL g1235 ( .A1(n_1158), .A2(n_1162), .B(n_1236), .C(n_1237), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1158), .B(n_1159), .Y(n_1269) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1159), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1161), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_1160), .A2(n_1194), .B1(n_1198), .B2(n_1200), .C(n_1203), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1160), .B(n_1162), .Y(n_1199) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1161), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1161), .B(n_1164), .Y(n_1243) );
OAI332xp33_ASAP7_75t_L g1203 ( .A1(n_1162), .A2(n_1168), .A3(n_1172), .B1(n_1204), .B2(n_1206), .B3(n_1207), .C1(n_1209), .C2(n_1211), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1162), .B(n_1165), .Y(n_1226) );
O2A1O1Ixp33_ASAP7_75t_L g1248 ( .A1(n_1163), .A2(n_1249), .B(n_1251), .C(n_1252), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_1165), .A2(n_1242), .B1(n_1244), .B2(n_1246), .Y(n_1241) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1172), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1168), .B(n_1196), .Y(n_1195) );
CKINVDCx6p67_ASAP7_75t_R g1201 ( .A(n_1168), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_1168), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1168), .B(n_1172), .Y(n_1254) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1171), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1169), .B(n_1171), .Y(n_1187) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1172), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1172), .B(n_1201), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1172), .B(n_1247), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1172), .B(n_1201), .Y(n_1280) );
AND2x4_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1175), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_1175), .Y(n_1239) );
OAI22xp5_ASAP7_75t_SL g1176 ( .A1(n_1177), .A2(n_1178), .B1(n_1179), .B2(n_1180), .Y(n_1176) );
NAND5xp2_ASAP7_75t_SL g1181 ( .A(n_1182), .B(n_1186), .C(n_1193), .D(n_1213), .E(n_1228), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1183), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1185), .Y(n_1236) );
OAI211xp5_ASAP7_75t_SL g1240 ( .A1(n_1187), .A2(n_1241), .B(n_1248), .C(n_1257), .Y(n_1240) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1189), .Y(n_1299) );
OAI21xp5_ASAP7_75t_L g1281 ( .A1(n_1190), .A2(n_1206), .B(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1195), .B(n_1230), .Y(n_1293) );
CKINVDCx6p67_ASAP7_75t_R g1196 ( .A(n_1197), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1197), .B(n_1205), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_1197), .A2(n_1214), .B1(n_1216), .B2(n_1218), .C(n_1220), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1197), .A2(n_1258), .B1(n_1263), .B2(n_1266), .Y(n_1257) );
O2A1O1Ixp33_ASAP7_75t_L g1294 ( .A1(n_1197), .A2(n_1256), .B(n_1295), .C(n_1296), .Y(n_1294) );
A2O1A1Ixp33_ASAP7_75t_L g1277 ( .A1(n_1198), .A2(n_1205), .B(n_1278), .C(n_1280), .Y(n_1277) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_1200), .A2(n_1212), .B1(n_1269), .B2(n_1270), .C(n_1275), .Y(n_1268) );
NOR2xp33_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
NOR2xp33_ASAP7_75t_L g1216 ( .A(n_1201), .B(n_1217), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1201), .B(n_1224), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1201), .B(n_1207), .Y(n_1292) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1202), .Y(n_1224) );
AOI21xp33_ASAP7_75t_L g1275 ( .A1(n_1202), .A2(n_1253), .B(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1207), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1207), .B(n_1298), .Y(n_1297) );
A2O1A1Ixp33_ASAP7_75t_L g1252 ( .A1(n_1209), .A2(n_1253), .B(n_1254), .C(n_1255), .Y(n_1252) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1212), .Y(n_1222) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1217), .Y(n_1251) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
OAI211xp5_ASAP7_75t_SL g1220 ( .A1(n_1221), .A2(n_1222), .B(n_1223), .C(n_1227), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1225), .Y(n_1223) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1226), .Y(n_1286) );
O2A1O1Ixp33_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1232), .B(n_1234), .C(n_1235), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NAND3xp33_ASAP7_75t_SL g1288 ( .A(n_1233), .B(n_1289), .C(n_1290), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1237), .B(n_1264), .Y(n_1263) );
INVx3_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
AOI21xp33_ASAP7_75t_L g1270 ( .A1(n_1239), .A2(n_1271), .B(n_1273), .Y(n_1270) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVxp67_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVxp67_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1262), .Y(n_1285) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NAND5xp2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1277), .C(n_1281), .D(n_1287), .E(n_1294), .Y(n_1267) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1280), .Y(n_1289) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1284), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
AOI21xp5_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1292), .B(n_1293), .Y(n_1287) );
INVxp67_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
BUFx2_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
NAND3xp33_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1321), .C(n_1339), .Y(n_1304) );
OAI31xp33_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1310), .A3(n_1316), .B(n_1320), .Y(n_1305) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_1314), .A2(n_1328), .B1(n_1329), .B2(n_1331), .Y(n_1327) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx2_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx2_ASAP7_75t_SL g1335 ( .A(n_1336), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1362), .Y(n_1339) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1343), .B1(n_1344), .B2(n_1345), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1364 ( .A1(n_1342), .A2(n_1358), .B1(n_1365), .B2(n_1368), .Y(n_1364) );
OAI22xp33_ASAP7_75t_L g1357 ( .A1(n_1343), .A2(n_1358), .B1(n_1359), .B2(n_1361), .Y(n_1357) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_1350), .A2(n_1355), .B1(n_1365), .B2(n_1368), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1353), .B1(n_1354), .B2(n_1355), .Y(n_1351) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
OAI33xp33_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1364), .A3(n_1369), .B1(n_1373), .B2(n_1374), .B3(n_1376), .Y(n_1362) );
INVx2_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_1367), .Y(n_1366) );
INVx4_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
BUFx2_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
CKINVDCx5p33_ASAP7_75t_R g1374 ( .A(n_1375), .Y(n_1374) );
CKINVDCx20_ASAP7_75t_R g1377 ( .A(n_1378), .Y(n_1377) );
CKINVDCx20_ASAP7_75t_R g1378 ( .A(n_1379), .Y(n_1378) );
INVx3_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVxp33_ASAP7_75t_SL g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1385), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1403), .Y(n_1385) );
AOI22xp5_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1399), .B1(n_1400), .B2(n_1402), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1408), .C(n_1413), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
OAI21xp5_ASAP7_75t_L g1425 ( .A1(n_1426), .A2(n_1427), .B(n_1428), .Y(n_1425) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
endmodule