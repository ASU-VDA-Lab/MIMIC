module fake_netlist_6_4003_n_1800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1800;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_47),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

INVx4_ASAP7_75t_R g167 ( 
.A(n_58),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_42),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_3),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_70),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_129),
.Y(n_177)
);

BUFx8_ASAP7_75t_SL g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_83),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_41),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_86),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_11),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_27),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_62),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_115),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_53),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_138),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_24),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_66),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_48),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_99),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_100),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_97),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_112),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_87),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_47),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_21),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_75),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_30),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_67),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_54),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_98),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_41),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_71),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_52),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_61),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_95),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_65),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_22),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_43),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_1),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_35),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_121),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_11),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_73),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_59),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_27),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_7),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_96),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_84),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_69),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_156),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_24),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_144),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_74),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_56),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_82),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_92),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_0),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_93),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_13),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_131),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_57),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_32),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_107),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_151),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_147),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_109),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_135),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_63),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_158),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_32),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_31),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_72),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_5),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_42),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_128),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_142),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_19),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_88),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_14),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_113),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_153),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_94),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_9),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_118),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_111),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_4),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_26),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_90),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_51),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_46),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_125),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_8),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_37),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_20),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_40),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_36),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_137),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_226),
.B(n_0),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_315),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_226),
.B(n_2),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_236),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_175),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_236),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_310),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_168),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_169),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_272),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_172),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_236),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_209),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_176),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_R g351 ( 
.A(n_194),
.B(n_2),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_284),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_177),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_179),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_183),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_187),
.B(n_6),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_185),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_186),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_191),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_192),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_175),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_166),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_166),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_196),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_182),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_170),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_170),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_197),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_182),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_198),
.B(n_210),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_173),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_199),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_200),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_205),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_202),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_232),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_204),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_198),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_242),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_210),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_R g390 ( 
.A(n_206),
.B(n_208),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_231),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_213),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_173),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_211),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_213),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_181),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_231),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_217),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_246),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_181),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_216),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_219),
.B(n_64),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_217),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_227),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_227),
.Y(n_406)
);

BUFx2_ASAP7_75t_SL g407 ( 
.A(n_184),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_241),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_184),
.B(n_8),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_246),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_221),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_241),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_165),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_253),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_180),
.Y(n_415)
);

BUFx6f_ASAP7_75t_SL g416 ( 
.A(n_205),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_189),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_228),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_261),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_232),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_261),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_347),
.B(n_195),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_234),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_380),
.B(n_234),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_343),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_396),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_203),
.B(n_195),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_333),
.B(n_205),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_348),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_354),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_339),
.B(n_203),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_251),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_407),
.B(n_262),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_360),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_339),
.B(n_285),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_366),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_368),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_368),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_353),
.B(n_285),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_374),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_378),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_339),
.B(n_189),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_400),
.B(n_218),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_237),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_218),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_335),
.B(n_265),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_392),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_392),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

CKINVDCx8_ASAP7_75t_R g496 ( 
.A(n_437),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_349),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_443),
.B(n_334),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_475),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_489),
.B(n_344),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_220),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_346),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_421),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_462),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_459),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

AND3x2_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_355),
.C(n_224),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

CKINVDCx11_ASAP7_75t_R g516 ( 
.A(n_437),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_350),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_428),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_489),
.B(n_356),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_363),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_365),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_489),
.B(n_373),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_377),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_438),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_489),
.B(n_381),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_382),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_429),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_474),
.A2(n_345),
.B1(n_418),
.B2(n_357),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_434),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_423),
.A2(n_351),
.B1(n_430),
.B2(n_171),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

BUFx6f_ASAP7_75t_SL g545 ( 
.A(n_488),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_489),
.B(n_384),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_476),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_489),
.B(n_493),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_386),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_438),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_429),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_434),
.B(n_415),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_220),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_432),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_479),
.B(n_224),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_489),
.B(n_394),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_489),
.B(n_402),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_463),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_488),
.A2(n_361),
.B1(n_304),
.B2(n_187),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_379),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_463),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_488),
.B(n_413),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_479),
.B(n_233),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_426),
.B(n_379),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_436),
.B(n_404),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_436),
.B(n_405),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_423),
.B(n_408),
.Y(n_576)
);

NOR3xp33_ASAP7_75t_L g577 ( 
.A(n_437),
.B(n_273),
.C(n_361),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_436),
.B(n_362),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_483),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_430),
.A2(n_291),
.B1(n_279),
.B2(n_275),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_439),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_488),
.B(n_277),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_487),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_488),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_479),
.B(n_364),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_491),
.A2(n_225),
.B1(n_290),
.B2(n_289),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_442),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_481),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_481),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_432),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_488),
.A2(n_304),
.B1(n_302),
.B2(n_325),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_491),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_488),
.A2(n_411),
.B1(n_399),
.B2(n_367),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_488),
.B(n_336),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_481),
.B(n_370),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_481),
.B(n_233),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_432),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_433),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_481),
.B(n_398),
.C(n_188),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_431),
.A2(n_238),
.B(n_235),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_442),
.Y(n_607)
);

OA22x2_ASAP7_75t_L g608 ( 
.A1(n_485),
.A2(n_295),
.B1(n_264),
.B2(n_263),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_239),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_488),
.A2(n_286),
.B1(n_302),
.B2(n_325),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_433),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_485),
.B(n_403),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_488),
.B(n_265),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_485),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_439),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_244),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_485),
.B(n_286),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_439),
.B(n_405),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_492),
.A2(n_250),
.B1(n_278),
.B2(n_249),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_485),
.A2(n_264),
.B1(n_303),
.B2(n_253),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_458),
.B(n_265),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_485),
.B(n_229),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_468),
.B(n_235),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_468),
.B(n_492),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_442),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_442),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_468),
.A2(n_301),
.B1(n_308),
.B2(n_259),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_433),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_433),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_468),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_494),
.B(n_383),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_435),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_435),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_494),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_442),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_435),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_442),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_435),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_468),
.B(n_238),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_450),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_442),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_341),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_549),
.B(n_477),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_508),
.B(n_616),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_608),
.A2(n_574),
.B1(n_575),
.B2(n_505),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_576),
.B(n_383),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_576),
.B(n_383),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_585),
.B(n_265),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_477),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_526),
.B(n_383),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_631),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_517),
.A2(n_287),
.B1(n_248),
.B2(n_255),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_625),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_586),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_585),
.B(n_265),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_585),
.B(n_312),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_528),
.A2(n_291),
.B1(n_247),
.B2(n_257),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_506),
.B(n_416),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_498),
.B(n_494),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_586),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_505),
.B(n_280),
.Y(n_662)
);

NOR2x1p5_ASAP7_75t_L g663 ( 
.A(n_555),
.B(n_174),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_604),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_592),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_477),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_543),
.B(n_416),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_538),
.B(n_416),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_523),
.B(n_477),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_523),
.B(n_477),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_524),
.B(n_431),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_524),
.B(n_431),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_570),
.B(n_312),
.Y(n_675)
);

AOI22x1_ASAP7_75t_L g676 ( 
.A1(n_615),
.A2(n_323),
.B1(n_247),
.B2(n_257),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_629),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_600),
.B(n_312),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_589),
.A2(n_319),
.B1(n_259),
.B2(n_260),
.C(n_263),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_547),
.B(n_431),
.Y(n_680)
);

AND2x2_ASAP7_75t_SL g681 ( 
.A(n_614),
.B(n_596),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_629),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_630),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_547),
.B(n_431),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_552),
.B(n_431),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_619),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_498),
.B(n_416),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_509),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_574),
.B(n_495),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_583),
.B(n_312),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_552),
.B(n_478),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_619),
.B(n_406),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_566),
.B(n_193),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_591),
.B(n_478),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_581),
.A2(n_495),
.B(n_295),
.C(n_301),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_499),
.B(n_229),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_630),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_513),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_591),
.B(n_478),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_633),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_633),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_598),
.B(n_478),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_563),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_566),
.A2(n_495),
.B(n_260),
.C(n_276),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_513),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_613),
.B(n_478),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_592),
.B(n_312),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_541),
.Y(n_710)
);

AND2x6_ASAP7_75t_SL g711 ( 
.A(n_588),
.B(n_268),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_567),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_566),
.A2(n_303),
.B(n_322),
.C(n_308),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_634),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_593),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_566),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_613),
.B(n_478),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_593),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_635),
.B(n_478),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_497),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_478),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_497),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_496),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_501),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_599),
.B(n_454),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_519),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_572),
.B(n_579),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_573),
.B(n_268),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_609),
.B(n_558),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_573),
.B(n_201),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_608),
.A2(n_451),
.B1(n_328),
.B2(n_276),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_519),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_540),
.B(n_212),
.C(n_207),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_573),
.B(n_406),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_580),
.B(n_584),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_573),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_505),
.A2(n_292),
.B1(n_281),
.B2(n_282),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_505),
.A2(n_293),
.B1(n_283),
.B2(n_288),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_480),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_558),
.B(n_480),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_634),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_601),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_578),
.B(n_223),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_601),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_505),
.B(n_480),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_605),
.B(n_230),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_565),
.A2(n_309),
.B1(n_332),
.B2(n_326),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_637),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_617),
.B(n_480),
.Y(n_752)
);

INVx8_ASAP7_75t_L g753 ( 
.A(n_560),
.Y(n_753)
);

AOI22x1_ASAP7_75t_SL g754 ( 
.A1(n_516),
.A2(n_258),
.B1(n_256),
.B2(n_254),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_632),
.B(n_480),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_548),
.A2(n_298),
.B1(n_294),
.B2(n_296),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_594),
.B(n_480),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_597),
.B(n_480),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_597),
.B(n_451),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_620),
.B(n_240),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_577),
.B(n_297),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_597),
.B(n_451),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_608),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_516),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_612),
.A2(n_623),
.B1(n_618),
.B2(n_571),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_453),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_610),
.A2(n_323),
.B1(n_320),
.B2(n_266),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_638),
.B(n_453),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_500),
.B(n_510),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_618),
.B(n_412),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_504),
.B(n_451),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_614),
.A2(n_622),
.B(n_618),
.C(n_628),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_504),
.B(n_442),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_500),
.B(n_453),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_504),
.B(n_215),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_641),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_639),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_500),
.B(n_453),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_502),
.A2(n_427),
.B(n_425),
.Y(n_779)
);

AND2x6_ASAP7_75t_L g780 ( 
.A(n_545),
.B(n_266),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_503),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_520),
.B(n_454),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_504),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_503),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_510),
.B(n_469),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_529),
.B(n_537),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_512),
.B(n_267),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_512),
.B(n_267),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_621),
.A2(n_279),
.B(n_269),
.C(n_332),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_514),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_624),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_507),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_624),
.B(n_458),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_507),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_512),
.B(n_269),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_511),
.Y(n_796)
);

BUFx8_ASAP7_75t_L g797 ( 
.A(n_496),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_560),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_546),
.B(n_243),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_645),
.A2(n_562),
.B(n_561),
.C(n_320),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_748),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_654),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_748),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_660),
.B(n_412),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_661),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_658),
.A2(n_275),
.B(n_316),
.C(n_314),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_682),
.B(n_245),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_729),
.A2(n_515),
.B(n_512),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_724),
.B(n_700),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_689),
.B(n_229),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_688),
.B(n_252),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_743),
.B(n_270),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_763),
.A2(n_305),
.B(n_309),
.C(n_314),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_689),
.B(n_515),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_707),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_691),
.B(n_560),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_678),
.A2(n_518),
.B(n_515),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_720),
.B(n_560),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_748),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_722),
.B(n_560),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_748),
.B(n_518),
.Y(n_821)
);

AO21x1_ASAP7_75t_L g822 ( 
.A1(n_759),
.A2(n_606),
.B(n_316),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_726),
.B(n_560),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_643),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_664),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_644),
.A2(n_536),
.B(n_518),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_665),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_667),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_652),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_732),
.B(n_571),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_687),
.B(n_571),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_723),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_757),
.A2(n_758),
.B(n_752),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_659),
.B(n_571),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_739),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_690),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_659),
.B(n_571),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_745),
.B(n_414),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_670),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_651),
.B(n_571),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_668),
.A2(n_525),
.B(n_521),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_677),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_650),
.A2(n_556),
.B(n_550),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_766),
.A2(n_556),
.B(n_550),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_414),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_716),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_705),
.B(n_602),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_661),
.B(n_550),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_734),
.B(n_271),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_712),
.B(n_602),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_789),
.A2(n_326),
.B(n_318),
.C(n_305),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_706),
.A2(n_318),
.B(n_622),
.C(n_222),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_768),
.A2(n_556),
.B(n_636),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_744),
.B(n_299),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_744),
.B(n_300),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_759),
.A2(n_556),
.B(n_636),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_694),
.B(n_602),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_715),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_762),
.A2(n_556),
.B(n_636),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_697),
.A2(n_522),
.B(n_603),
.C(n_595),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_661),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_602),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_736),
.B(n_602),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_718),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_669),
.A2(n_642),
.B(n_607),
.C(n_525),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_663),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_725),
.A2(n_640),
.B1(n_624),
.B2(n_602),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_735),
.B(n_624),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_760),
.B(n_306),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_666),
.B(n_640),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_683),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_797),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_666),
.B(n_640),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_681),
.A2(n_771),
.B(n_672),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_698),
.B(n_627),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_765),
.A2(n_646),
.B1(n_681),
.B2(n_786),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_760),
.B(n_311),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_646),
.B(n_647),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_684),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_710),
.B(n_454),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_769),
.A2(n_535),
.B(n_607),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_728),
.B(n_322),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_770),
.B(n_455),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_647),
.B(n_525),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_648),
.B(n_624),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_648),
.B(n_455),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_740),
.A2(n_535),
.B(n_607),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_671),
.A2(n_531),
.B(n_534),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_753),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_741),
.A2(n_534),
.B(n_531),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_673),
.A2(n_534),
.B(n_531),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_773),
.A2(n_533),
.B(n_539),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_695),
.B(n_455),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_674),
.A2(n_557),
.B(n_542),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_669),
.B(n_640),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_799),
.B(n_640),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_680),
.A2(n_557),
.B(n_542),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_716),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_799),
.B(n_640),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_728),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_685),
.A2(n_542),
.B(n_554),
.Y(n_901)
);

AO21x1_ASAP7_75t_L g902 ( 
.A1(n_649),
.A2(n_328),
.B(n_603),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_798),
.A2(n_545),
.B1(n_554),
.B2(n_590),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_686),
.A2(n_554),
.B(n_557),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_655),
.B(n_624),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_655),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_699),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_719),
.A2(n_544),
.B(n_527),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_695),
.B(n_313),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_750),
.B(n_568),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_728),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_679),
.A2(n_321),
.B(n_324),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_653),
.B(n_456),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_702),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_649),
.A2(n_544),
.B(n_527),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_776),
.B(n_568),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_755),
.A2(n_590),
.B(n_569),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_753),
.B(n_458),
.Y(n_919)
);

NAND2xp33_ASAP7_75t_L g920 ( 
.A(n_753),
.B(n_780),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_656),
.A2(n_590),
.B(n_569),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_730),
.B(n_317),
.Y(n_922)
);

O2A1O1Ixp5_ASAP7_75t_L g923 ( 
.A1(n_692),
.A2(n_551),
.B(n_564),
.C(n_559),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_656),
.A2(n_569),
.B(n_564),
.Y(n_924)
);

OR2x2_ASAP7_75t_SL g925 ( 
.A(n_711),
.B(n_167),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_790),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_747),
.B(n_456),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_784),
.B(n_530),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_657),
.A2(n_559),
.B(n_553),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_796),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_657),
.A2(n_553),
.B(n_551),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_774),
.A2(n_539),
.B(n_533),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_778),
.A2(n_530),
.B(n_447),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_703),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_747),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_777),
.B(n_484),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_675),
.A2(n_420),
.B(n_425),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_714),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_785),
.A2(n_447),
.B(n_448),
.Y(n_939)
);

INVx3_ASAP7_75t_SL g940 ( 
.A(n_761),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_713),
.B(n_329),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_782),
.A2(n_545),
.B1(n_458),
.B2(n_486),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_781),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_675),
.A2(n_448),
.B(n_449),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_737),
.B(n_484),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_792),
.B(n_794),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_756),
.B(n_709),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_742),
.B(n_484),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_780),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_772),
.A2(n_469),
.B(n_464),
.C(n_467),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_754),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_783),
.A2(n_448),
.B(n_449),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_709),
.B(n_330),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_738),
.B(n_486),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_797),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_751),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_733),
.B(n_791),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_767),
.B(n_456),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_692),
.A2(n_779),
.B(n_746),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_L g960 ( 
.A(n_749),
.B(n_464),
.C(n_467),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_693),
.A2(n_449),
.B(n_447),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_696),
.B(n_486),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_701),
.B(n_704),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_708),
.A2(n_449),
.B(n_444),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_767),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_662),
.B(n_464),
.C(n_467),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_878),
.B(n_731),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_955),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_854),
.A2(n_721),
.B(n_717),
.C(n_788),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_876),
.A2(n_767),
.B1(n_731),
.B2(n_676),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_896),
.A2(n_793),
.B(n_775),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_814),
.A2(n_775),
.B(n_788),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_899),
.A2(n_795),
.B(n_787),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_835),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_949),
.A2(n_780),
.B(n_440),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_832),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_927),
.B(n_780),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_880),
.B(n_804),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_935),
.B(n_469),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_815),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_854),
.B(n_490),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_949),
.A2(n_440),
.B(n_445),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_872),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_856),
.A2(n_419),
.B(n_425),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_869),
.A2(n_490),
.B(n_471),
.C(n_472),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_836),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_801),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_855),
.A2(n_469),
.B(n_764),
.C(n_472),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_855),
.B(n_490),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_877),
.A2(n_490),
.B(n_472),
.C(n_471),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_809),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_893),
.B(n_471),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_877),
.A2(n_446),
.B(n_441),
.C(n_444),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_815),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_825),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_935),
.B(n_9),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_963),
.A2(n_441),
.B(n_445),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_863),
.B(n_473),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_883),
.B(n_446),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_886),
.B(n_419),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_914),
.B(n_473),
.Y(n_1001)
);

NOR2x1p5_ASAP7_75t_L g1002 ( 
.A(n_829),
.B(n_473),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_801),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_802),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_914),
.B(n_10),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_926),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_926),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_846),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_868),
.A2(n_419),
.B(n_420),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_824),
.B(n_470),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_839),
.B(n_419),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_824),
.B(n_14),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_866),
.B(n_805),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_965),
.A2(n_470),
.B1(n_466),
.B2(n_461),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_909),
.B(n_470),
.C(n_466),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_801),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_833),
.A2(n_862),
.B(n_870),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_909),
.A2(n_458),
.B1(n_466),
.B2(n_461),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_873),
.A2(n_419),
.B(n_420),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_922),
.B(n_15),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_827),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_846),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_900),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_922),
.B(n_470),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_947),
.A2(n_466),
.B(n_461),
.C(n_460),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_898),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_828),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_801),
.B(n_461),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_959),
.A2(n_826),
.B(n_816),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_947),
.A2(n_460),
.B1(n_457),
.B2(n_450),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_895),
.A2(n_460),
.B1(n_457),
.B2(n_450),
.Y(n_1031)
);

AO32x2_ASAP7_75t_L g1032 ( 
.A1(n_903),
.A2(n_19),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_950),
.A2(n_460),
.B1(n_457),
.B2(n_450),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_941),
.A2(n_457),
.B(n_425),
.C(n_427),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_803),
.B(n_420),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_958),
.B(n_427),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_920),
.A2(n_843),
.B(n_859),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_874),
.A2(n_420),
.B1(n_425),
.B2(n_427),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_842),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_871),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_863),
.B(n_425),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_941),
.A2(n_427),
.B(n_458),
.C(n_33),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_845),
.B(n_427),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_810),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_806),
.A2(n_34),
.B(n_38),
.C(n_39),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_849),
.A2(n_34),
.B(n_39),
.C(n_43),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_898),
.B(n_44),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_SL g1048 ( 
.A1(n_834),
.A2(n_458),
.B(n_119),
.C(n_120),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_879),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_940),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_841),
.A2(n_458),
.B(n_117),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_849),
.B(n_458),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_953),
.A2(n_913),
.B(n_800),
.C(n_812),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_803),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_812),
.B(n_44),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_912),
.A2(n_45),
.B(n_51),
.C(n_52),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_803),
.B(n_130),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_813),
.A2(n_54),
.B(n_458),
.C(n_81),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_953),
.A2(n_77),
.B(n_89),
.C(n_91),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_884),
.A2(n_102),
.B(n_104),
.C(n_105),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_838),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_907),
.Y(n_1062)
);

OAI22x1_ASAP7_75t_L g1063 ( 
.A1(n_940),
.A2(n_140),
.B1(n_145),
.B2(n_148),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_858),
.A2(n_149),
.B1(n_157),
.B2(n_160),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_930),
.B(n_805),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_807),
.A2(n_957),
.B(n_875),
.C(n_811),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_905),
.A2(n_853),
.B(n_844),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_900),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_857),
.A2(n_911),
.B1(n_864),
.B2(n_807),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_811),
.A2(n_850),
.B(n_847),
.C(n_830),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_867),
.A2(n_889),
.B1(n_819),
.B2(n_837),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_911),
.B(n_861),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_882),
.B(n_960),
.C(n_831),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_819),
.B(n_906),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_819),
.B(n_882),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_808),
.A2(n_888),
.B(n_821),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_819),
.B(n_906),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_943),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_889),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_852),
.A2(n_960),
.B(n_885),
.C(n_851),
.Y(n_1080)
);

CKINVDCx6p67_ASAP7_75t_R g1081 ( 
.A(n_882),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_915),
.Y(n_1082)
);

AND2x6_ASAP7_75t_L g1083 ( 
.A(n_840),
.B(n_942),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_818),
.A2(n_823),
.B1(n_820),
.B2(n_966),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_925),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_934),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_938),
.B(n_956),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_966),
.A2(n_860),
.B(n_919),
.C(n_918),
.Y(n_1088)
);

AND2x2_ASAP7_75t_SL g1089 ( 
.A(n_962),
.B(n_946),
.Y(n_1089)
);

BUFx8_ASAP7_75t_L g1090 ( 
.A(n_951),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_937),
.B(n_848),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_889),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_936),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_945),
.B(n_954),
.C(n_910),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_908),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_889),
.A2(n_917),
.B1(n_817),
.B2(n_948),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_891),
.A2(n_897),
.B(n_894),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_902),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_901),
.A2(n_904),
.B(n_881),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_822),
.B(n_916),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_964),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_887),
.B(n_890),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_892),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_923),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_952),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1020),
.A2(n_933),
.B(n_921),
.C(n_924),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_978),
.B(n_932),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1037),
.A2(n_929),
.B(n_931),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_974),
.Y(n_1109)
);

CKINVDCx11_ASAP7_75t_R g1110 ( 
.A(n_976),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_970),
.A2(n_961),
.A3(n_939),
.B(n_944),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1053),
.A2(n_1046),
.B(n_996),
.C(n_1066),
.Y(n_1112)
);

OA21x2_ASAP7_75t_L g1113 ( 
.A1(n_1100),
.A2(n_1029),
.B(n_1076),
.Y(n_1113)
);

CKINVDCx11_ASAP7_75t_R g1114 ( 
.A(n_1081),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_970),
.A2(n_1025),
.A3(n_1099),
.B(n_1097),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_986),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1061),
.B(n_1055),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_981),
.A2(n_989),
.B(n_1024),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1061),
.B(n_991),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1004),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1070),
.A2(n_969),
.B(n_1084),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1079),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1067),
.A2(n_1017),
.B(n_984),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1078),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_967),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1102),
.A2(n_971),
.B(n_973),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1088),
.A2(n_1048),
.B(n_1042),
.C(n_1057),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1082),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1050),
.A2(n_1069),
.B1(n_1005),
.B2(n_1073),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1044),
.A2(n_1056),
.B(n_1045),
.C(n_988),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_987),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1094),
.A2(n_1080),
.B(n_1051),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_967),
.B(n_1089),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1012),
.A2(n_1047),
.B(n_991),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1093),
.A2(n_977),
.B(n_1071),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_977),
.A2(n_1071),
.B(n_1096),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1021),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1027),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_968),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1030),
.A2(n_1104),
.A3(n_1031),
.B(n_993),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_994),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1043),
.B(n_999),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_980),
.B(n_1006),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1000),
.A2(n_1052),
.B(n_1011),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1026),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1039),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1040),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1091),
.A2(n_1036),
.B(n_979),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_987),
.A2(n_1101),
.B(n_975),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1036),
.A2(n_979),
.B(n_1059),
.C(n_1074),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1008),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1095),
.A2(n_1103),
.B(n_1009),
.Y(n_1153)
);

AOI31xp67_ASAP7_75t_L g1154 ( 
.A1(n_1018),
.A2(n_1001),
.A3(n_1028),
.B(n_1077),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_1072),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1049),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1015),
.A2(n_997),
.B(n_985),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1062),
.Y(n_1158)
);

AOI31xp67_ASAP7_75t_L g1159 ( 
.A1(n_1010),
.A2(n_1035),
.A3(n_1065),
.B(n_1086),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1072),
.B(n_1065),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1002),
.B(n_1022),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_983),
.B(n_1090),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1014),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1030),
.A2(n_1031),
.A3(n_1014),
.B(n_1033),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1019),
.A2(n_972),
.B(n_1038),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_998),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1085),
.A2(n_1075),
.B1(n_1007),
.B2(n_998),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1023),
.B(n_1068),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1105),
.A2(n_1079),
.B(n_990),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_998),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1075),
.A2(n_1041),
.B1(n_1054),
.B2(n_1003),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1063),
.A2(n_982),
.A3(n_1083),
.B(n_1054),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_1003),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1075),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1060),
.A2(n_1034),
.B(n_1083),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1083),
.B(n_1041),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1003),
.Y(n_1177)
);

AOI211x1_ASAP7_75t_L g1178 ( 
.A1(n_1032),
.A2(n_1098),
.B(n_1064),
.C(n_1013),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1016),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1083),
.B(n_1041),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1058),
.A2(n_1092),
.B(n_1032),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1092),
.A2(n_585),
.B(n_1037),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1016),
.A2(n_585),
.B(n_1037),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1016),
.A2(n_1020),
.B1(n_877),
.B2(n_869),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_978),
.B(n_1061),
.Y(n_1185)
);

AO22x2_ASAP7_75t_L g1186 ( 
.A1(n_970),
.A2(n_1055),
.B1(n_876),
.B2(n_935),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1037),
.A2(n_1067),
.B(n_859),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_974),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_994),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_970),
.A2(n_822),
.A3(n_865),
.B(n_916),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1020),
.A2(n_877),
.B(n_869),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_994),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_974),
.Y(n_1193)
);

OAI22x1_ASAP7_75t_L g1194 ( 
.A1(n_1020),
.A2(n_877),
.B1(n_869),
.B2(n_914),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_978),
.B(n_645),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_978),
.B(n_645),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_SL g1197 ( 
.A(n_1020),
.B(n_698),
.C(n_869),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_978),
.B(n_645),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1020),
.A2(n_877),
.B(n_869),
.C(n_855),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1020),
.A2(n_877),
.B1(n_869),
.B2(n_855),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1061),
.B(n_576),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1053),
.A2(n_839),
.B(n_1020),
.C(n_878),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1061),
.B(n_576),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1003),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_970),
.A2(n_822),
.A3(n_865),
.B(n_916),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_L g1206 ( 
.A1(n_1020),
.A2(n_855),
.B(n_854),
.C(n_839),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_974),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1053),
.A2(n_855),
.B(n_854),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1037),
.A2(n_585),
.B(n_896),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_978),
.B(n_645),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1020),
.B(n_341),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_994),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1020),
.A2(n_877),
.B(n_869),
.C(n_855),
.Y(n_1213)
);

AO21x1_ASAP7_75t_L g1214 ( 
.A1(n_1020),
.A2(n_1066),
.B(n_839),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1020),
.B(n_724),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_978),
.B(n_645),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1020),
.A2(n_935),
.B1(n_877),
.B2(n_869),
.Y(n_1217)
);

AOI221xp5_ASAP7_75t_L g1218 ( 
.A1(n_1020),
.A2(n_877),
.B1(n_869),
.B2(n_679),
.C(n_854),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_968),
.Y(n_1219)
);

AOI211x1_ASAP7_75t_L g1220 ( 
.A1(n_1055),
.A2(n_658),
.B(n_986),
.C(n_974),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1020),
.A2(n_877),
.B(n_869),
.C(n_855),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1053),
.A2(n_855),
.B(n_854),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_978),
.B(n_645),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_994),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1037),
.A2(n_1067),
.B(n_859),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_994),
.Y(n_1227)
);

AO32x2_ASAP7_75t_L g1228 ( 
.A1(n_970),
.A2(n_1014),
.A3(n_876),
.B1(n_658),
.B2(n_1030),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1020),
.B(n_341),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_974),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_1003),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1003),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1075),
.B(n_976),
.Y(n_1233)
);

CKINVDCx6p67_ASAP7_75t_R g1234 ( 
.A(n_976),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1020),
.A2(n_855),
.B1(n_854),
.B2(n_869),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1053),
.A2(n_855),
.B(n_854),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_968),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1020),
.B(n_341),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_974),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1020),
.B(n_341),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1020),
.A2(n_877),
.B(n_869),
.C(n_855),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1109),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1207),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1235),
.A2(n_1200),
.B1(n_1218),
.B2(n_1241),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1116),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1189),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1120),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1217),
.A2(n_1197),
.B1(n_1222),
.B2(n_1208),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1236),
.A2(n_1240),
.B1(n_1238),
.B2(n_1229),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1211),
.A2(n_1194),
.B1(n_1184),
.B2(n_1214),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1125),
.B(n_1199),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1140),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1188),
.Y(n_1253)
);

INVx3_ASAP7_75t_SL g1254 ( 
.A(n_1237),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1193),
.Y(n_1255)
);

INVx5_ASAP7_75t_SL g1256 ( 
.A(n_1234),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1191),
.A2(n_1215),
.B1(n_1129),
.B2(n_1196),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1213),
.A2(n_1221),
.B1(n_1178),
.B2(n_1216),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1186),
.A2(n_1121),
.B1(n_1162),
.B2(n_1185),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1186),
.A2(n_1135),
.B1(n_1132),
.B2(n_1134),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_1131),
.B(n_1173),
.Y(n_1261)
);

CKINVDCx6p67_ASAP7_75t_R g1262 ( 
.A(n_1110),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1168),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1114),
.Y(n_1264)
);

INVx6_ASAP7_75t_L g1265 ( 
.A(n_1140),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1195),
.A2(n_1223),
.B1(n_1198),
.B2(n_1210),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1219),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1176),
.A2(n_1180),
.B1(n_1203),
.B2(n_1201),
.Y(n_1268)
);

BUFx2_ASAP7_75t_SL g1269 ( 
.A(n_1173),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1117),
.A2(n_1143),
.B1(n_1149),
.B2(n_1174),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1144),
.A2(n_1119),
.B(n_1161),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1175),
.A2(n_1155),
.B1(n_1225),
.B2(n_1206),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1233),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1107),
.A2(n_1170),
.B1(n_1166),
.B2(n_1224),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1112),
.A2(n_1136),
.B(n_1202),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1160),
.B(n_1138),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1130),
.A2(n_1146),
.B(n_1192),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1131),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1173),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1212),
.Y(n_1280)
);

BUFx2_ASAP7_75t_R g1281 ( 
.A(n_1179),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1152),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1230),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1167),
.A2(n_1233),
.B1(n_1142),
.B2(n_1227),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1239),
.Y(n_1285)
);

INVx8_ASAP7_75t_L g1286 ( 
.A(n_1231),
.Y(n_1286)
);

OAI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1128),
.A2(n_1124),
.B(n_1181),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1163),
.A2(n_1157),
.B1(n_1148),
.B2(n_1139),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1133),
.A2(n_1147),
.B1(n_1156),
.B2(n_1158),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1137),
.A2(n_1171),
.B1(n_1145),
.B2(n_1169),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1231),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1113),
.A2(n_1126),
.B1(n_1118),
.B2(n_1122),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1151),
.A2(n_1127),
.B1(n_1177),
.B2(n_1183),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_1231),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1204),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1204),
.Y(n_1296)
);

BUFx8_ASAP7_75t_SL g1297 ( 
.A(n_1232),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1220),
.B(n_1172),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1232),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1159),
.Y(n_1300)
);

INVx4_ASAP7_75t_SL g1301 ( 
.A(n_1172),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1172),
.B(n_1164),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1228),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1150),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1153),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1182),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1154),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1111),
.Y(n_1308)
);

BUFx8_ASAP7_75t_L g1309 ( 
.A(n_1228),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1228),
.Y(n_1310)
);

BUFx4f_ASAP7_75t_SL g1311 ( 
.A(n_1106),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1165),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1115),
.Y(n_1313)
);

CKINVDCx6p67_ASAP7_75t_R g1314 ( 
.A(n_1111),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1115),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1141),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1141),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1209),
.A2(n_1187),
.B1(n_1226),
.B2(n_1108),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1123),
.A2(n_1164),
.B1(n_1190),
.B2(n_1205),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1164),
.A2(n_1190),
.B1(n_1205),
.B2(n_1141),
.Y(n_1320)
);

BUFx5_ASAP7_75t_L g1321 ( 
.A(n_1205),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1174),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1219),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1218),
.A2(n_1200),
.B1(n_1235),
.B2(n_1217),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1237),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1173),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1109),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1235),
.B(n_1125),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1219),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1235),
.A2(n_1200),
.B1(n_1218),
.B2(n_1213),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1109),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1109),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1109),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1109),
.Y(n_1334)
);

CKINVDCx6p67_ASAP7_75t_R g1335 ( 
.A(n_1110),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1119),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1189),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1109),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1208),
.A2(n_1236),
.B(n_1222),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1109),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1131),
.Y(n_1341)
);

CKINVDCx6p67_ASAP7_75t_R g1342 ( 
.A(n_1110),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1173),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1217),
.A2(n_1240),
.B1(n_1238),
.B2(n_1211),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1189),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1218),
.A2(n_1200),
.B1(n_1235),
.B2(n_1217),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1219),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_1236),
.B(n_1222),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1119),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1185),
.B(n_978),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1185),
.B(n_978),
.Y(n_1351)
);

INVx6_ASAP7_75t_L g1352 ( 
.A(n_1140),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1119),
.Y(n_1353)
);

BUFx4f_ASAP7_75t_L g1354 ( 
.A(n_1234),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1217),
.A2(n_1240),
.B1(n_1238),
.B2(n_1211),
.Y(n_1355)
);

BUFx4f_ASAP7_75t_SL g1356 ( 
.A(n_1219),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1217),
.A2(n_1240),
.B1(n_1238),
.B2(n_1211),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1119),
.B(n_1201),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_1237),
.Y(n_1359)
);

INVx5_ASAP7_75t_L g1360 ( 
.A(n_1131),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1235),
.B(n_1125),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1109),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1219),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1173),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1140),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1237),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1316),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1317),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1302),
.B(n_1308),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1310),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1310),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1245),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1301),
.B(n_1275),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1345),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1302),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1336),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1273),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1313),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1309),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1315),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1300),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1323),
.Y(n_1382)
);

BUFx8_ASAP7_75t_SL g1383 ( 
.A(n_1347),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1287),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1298),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1244),
.B(n_1330),
.C(n_1344),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1336),
.Y(n_1388)
);

NOR2x1_ASAP7_75t_L g1389 ( 
.A(n_1251),
.B(n_1275),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1309),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1339),
.A2(n_1348),
.B(n_1307),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1298),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1305),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1303),
.B(n_1259),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1253),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1273),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1329),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1318),
.A2(n_1292),
.B(n_1290),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1255),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1339),
.A2(n_1348),
.B(n_1293),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1305),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1244),
.A2(n_1330),
.B1(n_1324),
.B2(n_1346),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1301),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1259),
.B(n_1260),
.Y(n_1405)
);

INVxp33_ASAP7_75t_L g1406 ( 
.A(n_1350),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1301),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1249),
.A2(n_1357),
.B1(n_1355),
.B2(n_1250),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1311),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1321),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1321),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1280),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1306),
.B(n_1283),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1320),
.B(n_1248),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1321),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1285),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1257),
.A2(n_1258),
.B1(n_1361),
.B2(n_1328),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1286),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1251),
.A2(n_1258),
.B(n_1328),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1276),
.B(n_1351),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1306),
.B(n_1312),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1321),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1314),
.B(n_1349),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1321),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1312),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1252),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1243),
.Y(n_1427)
);

AND2x4_ASAP7_75t_SL g1428 ( 
.A(n_1274),
.B(n_1326),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1288),
.A2(n_1289),
.B(n_1361),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1327),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1319),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1304),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1332),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1333),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1242),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1349),
.B(n_1358),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1331),
.B(n_1338),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1266),
.B(n_1270),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1334),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1360),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1263),
.Y(n_1442)
);

BUFx12f_ASAP7_75t_L g1443 ( 
.A(n_1264),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1252),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1356),
.B(n_1363),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1325),
.B(n_1366),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1246),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1362),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1284),
.A2(n_1271),
.B1(n_1352),
.B2(n_1365),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1337),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1272),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1268),
.A2(n_1277),
.B(n_1295),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1282),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1278),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1282),
.B(n_1299),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1341),
.A2(n_1261),
.B(n_1269),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1286),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1281),
.B(n_1296),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1261),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1354),
.A2(n_1343),
.B(n_1286),
.C(n_1294),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1326),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1364),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1364),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1394),
.B(n_1281),
.Y(n_1464)
);

NAND2x1_ASAP7_75t_L g1465 ( 
.A(n_1432),
.B(n_1456),
.Y(n_1465)
);

OAI211xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1387),
.A2(n_1403),
.B(n_1417),
.C(n_1408),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1420),
.B(n_1267),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1426),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1441),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1376),
.B(n_1322),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1431),
.B(n_1365),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1388),
.B(n_1322),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1437),
.B(n_1254),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1398),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1460),
.A2(n_1291),
.B(n_1265),
.C(n_1297),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1405),
.A2(n_1354),
.B1(n_1279),
.B2(n_1262),
.C(n_1335),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1453),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1389),
.A2(n_1279),
.B(n_1265),
.C(n_1256),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1437),
.B(n_1342),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1372),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1401),
.A2(n_1359),
.B(n_1256),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1374),
.B(n_1359),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1431),
.B(n_1370),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1385),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1389),
.A2(n_1451),
.B(n_1405),
.C(n_1429),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1451),
.A2(n_1439),
.B1(n_1414),
.B2(n_1406),
.C(n_1384),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1379),
.B(n_1390),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1429),
.A2(n_1419),
.B(n_1409),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1409),
.A2(n_1449),
.B(n_1399),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1452),
.B(n_1384),
.C(n_1423),
.Y(n_1492)
);

A2O1A1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1432),
.A2(n_1414),
.B(n_1373),
.C(n_1399),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1371),
.B(n_1413),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1432),
.A2(n_1373),
.B(n_1428),
.C(n_1413),
.Y(n_1495)
);

BUFx12f_ASAP7_75t_SL g1496 ( 
.A(n_1458),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1432),
.A2(n_1442),
.B(n_1459),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1421),
.B(n_1400),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_SL g1501 ( 
.A(n_1445),
.B(n_1446),
.C(n_1461),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1459),
.A2(n_1452),
.B(n_1461),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1381),
.A2(n_1410),
.B(n_1411),
.Y(n_1503)
);

AOI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1447),
.A2(n_1450),
.B1(n_1438),
.B2(n_1378),
.C(n_1380),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1438),
.B(n_1427),
.Y(n_1505)
);

AOI211xp5_ASAP7_75t_L g1506 ( 
.A1(n_1455),
.A2(n_1396),
.B(n_1412),
.C(n_1458),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1373),
.A2(n_1428),
.B(n_1421),
.C(n_1377),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1416),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1381),
.A2(n_1415),
.B(n_1424),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1438),
.B(n_1427),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1426),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1373),
.B(n_1404),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1383),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1386),
.B(n_1392),
.Y(n_1514)
);

NAND4xp25_ASAP7_75t_L g1515 ( 
.A(n_1455),
.B(n_1433),
.C(n_1377),
.D(n_1448),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1396),
.A2(n_1428),
.B1(n_1377),
.B2(n_1452),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1433),
.B(n_1448),
.C(n_1436),
.D(n_1440),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1404),
.B(n_1407),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_SL g1519 ( 
.A1(n_1418),
.A2(n_1457),
.B(n_1407),
.C(n_1454),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1369),
.B(n_1386),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1369),
.B(n_1392),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1393),
.B(n_1402),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1466),
.A2(n_1452),
.B1(n_1382),
.B2(n_1443),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1391),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1478),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1503),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1481),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1514),
.B(n_1375),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1514),
.B(n_1375),
.Y(n_1530)
);

INVx5_ASAP7_75t_L g1531 ( 
.A(n_1469),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.B(n_1391),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1498),
.B(n_1391),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1391),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1520),
.B(n_1380),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1521),
.B(n_1402),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1512),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1522),
.B(n_1393),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1522),
.B(n_1367),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1486),
.B(n_1367),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1509),
.Y(n_1541)
);

OAI221xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1488),
.A2(n_1426),
.B1(n_1444),
.B2(n_1434),
.C(n_1435),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1506),
.A2(n_1444),
.B1(n_1382),
.B2(n_1430),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1493),
.B(n_1422),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1485),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1465),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1475),
.B(n_1425),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1493),
.B(n_1368),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1494),
.B(n_1368),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1523),
.A2(n_1491),
.B1(n_1464),
.B2(n_1492),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1545),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1490),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1541),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1532),
.B(n_1505),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1531),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1547),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1524),
.B(n_1502),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1526),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1533),
.B(n_1484),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1542),
.A2(n_1487),
.B1(n_1464),
.B2(n_1501),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_SL g1563 ( 
.A1(n_1543),
.A2(n_1482),
.B(n_1462),
.C(n_1463),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1542),
.A2(n_1504),
.B1(n_1476),
.B2(n_1477),
.C(n_1515),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1545),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1527),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_1508),
.Y(n_1568)
);

OAI33xp33_ASAP7_75t_L g1569 ( 
.A1(n_1543),
.A2(n_1540),
.A3(n_1525),
.B1(n_1536),
.B2(n_1535),
.B3(n_1517),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1527),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1495),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1495),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1528),
.B(n_1500),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1549),
.B(n_1507),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1549),
.B(n_1507),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1549),
.B(n_1544),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1567),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1552),
.B(n_1525),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1569),
.B(n_1397),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1530),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1567),
.Y(n_1586)
);

NAND2x1_ASAP7_75t_L g1587 ( 
.A(n_1565),
.B(n_1544),
.Y(n_1587)
);

OAI322xp33_ASAP7_75t_L g1588 ( 
.A1(n_1562),
.A2(n_1535),
.A3(n_1536),
.B1(n_1538),
.B2(n_1540),
.C1(n_1530),
.C2(n_1539),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1567),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1580),
.B(n_1537),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1538),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1580),
.B(n_1537),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1571),
.B(n_1574),
.Y(n_1594)
);

NOR4xp25_ASAP7_75t_SL g1595 ( 
.A(n_1558),
.B(n_1479),
.C(n_1476),
.D(n_1519),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1570),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1566),
.B(n_1550),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1546),
.Y(n_1598)
);

OAI31xp33_ASAP7_75t_L g1599 ( 
.A1(n_1562),
.A2(n_1479),
.A3(n_1467),
.B(n_1489),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1570),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1561),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1565),
.B(n_1547),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1554),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1572),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1551),
.B(n_1516),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1554),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1554),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1560),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1566),
.B(n_1550),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1559),
.B(n_1550),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1560),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1553),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1610),
.A2(n_1551),
.B1(n_1564),
.B2(n_1569),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1553),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1587),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1589),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1616),
.B(n_1576),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1576),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1600),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_L g1629 ( 
.A(n_1602),
.B(n_1564),
.C(n_1563),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1594),
.B(n_1553),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1583),
.B(n_1559),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1603),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1587),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1594),
.B(n_1575),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1581),
.B(n_1575),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1593),
.B(n_1576),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1590),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1583),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1585),
.B(n_1561),
.Y(n_1645)
);

INVxp33_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1575),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1593),
.B(n_1568),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1558),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1586),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1586),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1607),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1602),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1611),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1590),
.A2(n_1579),
.B(n_1565),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1596),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1631),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1592),
.Y(n_1663)
);

NAND4xp25_ASAP7_75t_L g1664 ( 
.A(n_1620),
.B(n_1563),
.C(n_1602),
.D(n_1471),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1653),
.B(n_1658),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1592),
.Y(n_1666)
);

OAI322xp33_ASAP7_75t_L g1667 ( 
.A1(n_1620),
.A2(n_1597),
.A3(n_1615),
.B1(n_1585),
.B2(n_1604),
.C1(n_1588),
.C2(n_1617),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1643),
.B(n_1605),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1637),
.B(n_1606),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1623),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_1597),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1629),
.B(n_1565),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.B(n_1611),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1638),
.B(n_1615),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1652),
.B(n_1596),
.Y(n_1679)
);

AND4x1_ASAP7_75t_L g1680 ( 
.A(n_1619),
.B(n_1579),
.C(n_1595),
.D(n_1611),
.Y(n_1680)
);

NAND4xp25_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1471),
.C(n_1483),
.D(n_1470),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1626),
.B(n_1577),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1657),
.B(n_1606),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1646),
.B(n_1588),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1657),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1621),
.B(n_1601),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1621),
.B(n_1601),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1626),
.B(n_1577),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1627),
.B(n_1641),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1627),
.B(n_1568),
.Y(n_1691)
);

AND2x2_ASAP7_75t_SL g1692 ( 
.A(n_1649),
.B(n_1606),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1624),
.B(n_1608),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1635),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1647),
.B(n_1579),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1624),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1651),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1659),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1685),
.B(n_1660),
.C(n_1630),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1685),
.A2(n_1595),
.B(n_1660),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1675),
.A2(n_1650),
.B1(n_1642),
.B2(n_1625),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1667),
.A2(n_1630),
.B1(n_1628),
.B2(n_1659),
.C(n_1623),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1675),
.A2(n_1628),
.B(n_1651),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1696),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1669),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1692),
.B(n_1647),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1680),
.A2(n_1644),
.B(n_1636),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1686),
.B(n_1622),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1664),
.A2(n_1606),
.B(n_1649),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1692),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1679),
.A2(n_1622),
.B1(n_1632),
.B2(n_1661),
.C(n_1654),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1679),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1696),
.A2(n_1473),
.B(n_1480),
.C(n_1606),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1662),
.B(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1671),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1662),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1666),
.B(n_1632),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1665),
.B(n_1645),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1694),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1673),
.Y(n_1723)
);

AOI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1661),
.B(n_1654),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1716),
.B(n_1698),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_SL g1726 ( 
.A(n_1702),
.B(n_1700),
.C(n_1699),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1706),
.B(n_1683),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1710),
.B(n_1670),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1716),
.B(n_1681),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1707),
.A2(n_1704),
.B1(n_1714),
.B2(n_1708),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1707),
.A2(n_1670),
.B1(n_1668),
.B2(n_1690),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1704),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1715),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1668),
.Y(n_1735)
);

O2A1O1Ixp5_ASAP7_75t_L g1736 ( 
.A1(n_1703),
.A2(n_1673),
.B(n_1693),
.C(n_1687),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1701),
.A2(n_1674),
.B1(n_1672),
.B2(n_1697),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1718),
.B(n_1678),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1717),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1709),
.A2(n_1688),
.B(n_1687),
.Y(n_1740)
);

OAI31xp33_ASAP7_75t_L g1741 ( 
.A1(n_1699),
.A2(n_1689),
.A3(n_1682),
.B(n_1691),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1723),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1711),
.B(n_1648),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1721),
.Y(n_1744)
);

INVxp33_ASAP7_75t_L g1745 ( 
.A(n_1730),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1727),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1728),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1726),
.B(n_1443),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1732),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1725),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1742),
.B(n_1720),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1729),
.B(n_1722),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1744),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1742),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1733),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1734),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1731),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1748),
.A2(n_1726),
.B1(n_1737),
.B2(n_1743),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1749),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1749),
.Y(n_1760)
);

AOI21xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1745),
.A2(n_1748),
.B(n_1737),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_L g1762 ( 
.A(n_1747),
.B(n_1736),
.C(n_1741),
.D(n_1735),
.Y(n_1762)
);

NAND4xp25_ASAP7_75t_L g1763 ( 
.A(n_1752),
.B(n_1736),
.C(n_1740),
.D(n_1739),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1751),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1751),
.B(n_1750),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1758),
.A2(n_1753),
.B1(n_1754),
.B2(n_1755),
.Y(n_1767)
);

OAI21xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1763),
.A2(n_1724),
.B(n_1756),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1764),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1762),
.A2(n_1721),
.B1(n_1713),
.B2(n_1719),
.C(n_1693),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1513),
.Y(n_1771)
);

AOI321xp33_ASAP7_75t_L g1772 ( 
.A1(n_1765),
.A2(n_1688),
.A3(n_1474),
.B1(n_1636),
.B2(n_1644),
.C(n_1656),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1757),
.B1(n_1766),
.B2(n_1759),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1768),
.A2(n_1760),
.B1(n_1656),
.B2(n_1655),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1444),
.C(n_1641),
.D(n_1497),
.Y(n_1775)
);

OAI211xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1769),
.A2(n_1655),
.B(n_1644),
.C(n_1636),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1770),
.A2(n_1513),
.B(n_1772),
.C(n_1655),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1771),
.B(n_1598),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1768),
.A2(n_1656),
.B(n_1558),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1773),
.Y(n_1780)
);

NAND4xp75_ASAP7_75t_L g1781 ( 
.A(n_1779),
.B(n_1557),
.C(n_1418),
.D(n_1457),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1778),
.Y(n_1782)
);

INVx4_ASAP7_75t_L g1783 ( 
.A(n_1774),
.Y(n_1783)
);

O2A1O1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1777),
.A2(n_1557),
.B(n_1555),
.C(n_1573),
.Y(n_1784)
);

NOR2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1775),
.Y(n_1785)
);

OR3x2_ASAP7_75t_L g1786 ( 
.A(n_1782),
.B(n_1776),
.C(n_1496),
.Y(n_1786)
);

OAI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1784),
.A2(n_1511),
.B(n_1468),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1785),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1786),
.B1(n_1783),
.B2(n_1781),
.Y(n_1789)
);

INVx3_ASAP7_75t_SL g1790 ( 
.A(n_1789),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_SL g1791 ( 
.A1(n_1789),
.A2(n_1783),
.B(n_1787),
.Y(n_1791)
);

OAI21x1_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1618),
.B(n_1614),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1790),
.Y(n_1793)
);

XNOR2xp5_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1468),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1618),
.B(n_1607),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1794),
.B(n_1618),
.C(n_1614),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1795),
.B1(n_1557),
.B2(n_1547),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1797),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1607),
.B1(n_1614),
.B2(n_1613),
.C(n_1612),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1511),
.B(n_1613),
.C(n_1612),
.Y(n_1800)
);


endmodule