module fake_jpeg_25627_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_21),
.CON(n_65),
.SN(n_65)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_17),
.B1(n_21),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_76),
.B1(n_19),
.B2(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_35),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_37),
.B(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_29),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_68),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_17),
.B1(n_31),
.B2(n_28),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_37),
.B1(n_31),
.B2(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_17),
.B1(n_22),
.B2(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_43),
.B1(n_45),
.B2(n_39),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_45),
.B1(n_22),
.B2(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_93),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_29),
.B(n_0),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_92),
.B(n_25),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_23),
.Y(n_140)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_107),
.B1(n_108),
.B2(n_54),
.Y(n_120)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_29),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_109),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_113),
.B1(n_98),
.B2(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_61),
.A2(n_29),
.B(n_23),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_106),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_48),
.B1(n_34),
.B2(n_35),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_51),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_37),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_58),
.Y(n_135)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_1),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_138),
.B1(n_146),
.B2(n_91),
.Y(n_173)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_65),
.C(n_23),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_141),
.C(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_139),
.Y(n_154)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_60),
.B1(n_56),
.B2(n_52),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_87),
.B1(n_86),
.B2(n_103),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_116),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_99),
.B(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_77),
.C(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_4),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_67),
.B1(n_73),
.B2(n_34),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_114),
.B1(n_112),
.B2(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_25),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_25),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_117),
.B(n_80),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_161),
.B(n_167),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_137),
.CI(n_122),
.CON(n_190),
.SN(n_190)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_82),
.B(n_100),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_173),
.B1(n_180),
.B2(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_34),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_91),
.B(n_87),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_177),
.Y(n_201)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_170),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_132),
.B(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_178),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_107),
.B1(n_83),
.B2(n_33),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_110),
.B(n_5),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_130),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_13),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_120),
.B1(n_146),
.B2(n_142),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_32),
.Y(n_181)
);

AND2x4_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_141),
.B1(n_140),
.B2(n_121),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_121),
.B(n_32),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_162),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_126),
.B1(n_137),
.B2(n_144),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_202),
.B1(n_203),
.B2(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_208),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_144),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_204),
.C(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_154),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_7),
.C(n_10),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_10),
.C(n_11),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_176),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_13),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_177),
.C(n_178),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_181),
.B1(n_158),
.B2(n_161),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_221),
.B1(n_241),
.B2(n_208),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_212),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_234),
.B(n_197),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_232),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_181),
.B1(n_170),
.B2(n_172),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_181),
.B(n_172),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_224),
.B(n_239),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_160),
.B(n_183),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_210),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_153),
.B1(n_168),
.B2(n_171),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_189),
.B1(n_214),
.B2(n_202),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_193),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_178),
.C(n_155),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_237),
.C(n_204),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_178),
.B(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_243),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_162),
.C(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_197),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_169),
.B(n_15),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_189),
.A2(n_169),
.B1(n_15),
.B2(n_16),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_14),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_245),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_203),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_253),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_201),
.C(n_235),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_220),
.B1(n_232),
.B2(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_186),
.C(n_237),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_234),
.B(n_185),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_233),
.C(n_226),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_226),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_275),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_247),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_241),
.B1(n_218),
.B2(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_253),
.B1(n_264),
.B2(n_245),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_206),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_224),
.C(n_223),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_228),
.C(n_227),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_211),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_282),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_291),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_262),
.B(n_254),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_287),
.B(n_266),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_257),
.CI(n_254),
.CON(n_288),
.SN(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_248),
.B1(n_247),
.B2(n_205),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_216),
.B(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_278),
.C(n_269),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_296),
.C(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_270),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_307),
.B1(n_276),
.B2(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_274),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_312),
.C(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_296),
.C(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_289),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_318),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_303),
.B1(n_300),
.B2(n_304),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_321),
.B(n_14),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_281),
.B(n_199),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_317),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_316),
.C(n_322),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_312),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule