module fake_aes_5891_n_550 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_550);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_550;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_235;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_14), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_2), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_78), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_57), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_33), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_77), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_72), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_6), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_58), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_43), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_29), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
NOR2xp67_ASAP7_75t_L g99 ( .A(n_74), .B(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_50), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_69), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_1), .Y(n_105) );
BUFx5_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_30), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_44), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_63), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_36), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_15), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_107), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_106), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
NOR2xp33_ASAP7_75t_R g122 ( .A(n_92), .B(n_31), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_106), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_98), .B(n_0), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_105), .B(n_1), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_85), .B(n_3), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_81), .B(n_3), .Y(n_129) );
INVx5_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_79), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_106), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
NOR2xp33_ASAP7_75t_R g137 ( .A(n_92), .B(n_34), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_105), .B(n_4), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_90), .B(n_4), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_135), .B(n_103), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_125), .A2(n_109), .B1(n_80), .B2(n_108), .Y(n_146) );
NAND3xp33_ASAP7_75t_L g147 ( .A(n_117), .B(n_88), .C(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_135), .B(n_95), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_132), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_131), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_117), .B(n_90), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_132), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_120), .B(n_121), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_120), .B(n_109), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_125), .B(n_87), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_133), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_121), .B(n_93), .C(n_115), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_129), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_128), .B(n_103), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
BUFx4_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_128), .B(n_111), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_161), .B(n_122), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_151), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_162), .B(n_136), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_162), .B(n_136), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_152), .B(n_146), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_165), .B(n_126), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_152), .B(n_127), .Y(n_176) );
NOR3xp33_ASAP7_75t_SL g177 ( .A(n_145), .B(n_124), .C(n_111), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_157), .A2(n_138), .B1(n_125), .B2(n_127), .Y(n_178) );
NOR3xp33_ASAP7_75t_SL g179 ( .A(n_149), .B(n_100), .C(n_89), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_157), .A2(n_138), .B1(n_112), .B2(n_116), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_138), .B1(n_127), .B2(n_134), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_164), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_156), .A2(n_134), .B(n_123), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_155), .B(n_141), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_155), .B(n_138), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_164), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_147), .B(n_88), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_141), .B(n_137), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_147), .B(n_110), .Y(n_198) );
OR2x6_ASAP7_75t_L g199 ( .A(n_195), .B(n_159), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_167), .A2(n_113), .B1(n_89), .B2(n_94), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_189), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_170), .A2(n_159), .B(n_160), .C(n_163), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_184), .A2(n_163), .B1(n_160), .B2(n_158), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_191), .A2(n_158), .B(n_142), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_196), .A2(n_134), .B1(n_123), .B2(n_132), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_192), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_195), .B(n_113), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_192), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_189), .B(n_91), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_188), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_168), .B(n_148), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_168), .B(n_148), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_196), .A2(n_142), .B1(n_130), .B2(n_118), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_169), .B(n_130), .Y(n_218) );
BUFx6f_ASAP7_75t_SL g219 ( .A(n_196), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_172), .B(n_130), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_187), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_180), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_188), .B(n_130), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_181), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
NOR2x1_ASAP7_75t_SL g227 ( .A(n_185), .B(n_94), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_166), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_187), .Y(n_229) );
AOI33xp33_ASAP7_75t_L g230 ( .A1(n_181), .A2(n_91), .A3(n_93), .B1(n_104), .B2(n_96), .B3(n_102), .Y(n_230) );
BUFx8_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
BUFx2_ASAP7_75t_SL g232 ( .A(n_219), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_224), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_224), .B(n_185), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_217), .A2(n_174), .B(n_182), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_208), .B(n_171), .Y(n_236) );
CKINVDCx12_ASAP7_75t_R g237 ( .A(n_208), .Y(n_237) );
OAI21x1_ASAP7_75t_SL g238 ( .A1(n_227), .A2(n_178), .B(n_186), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_207), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_225), .A2(n_190), .B1(n_196), .B2(n_194), .Y(n_241) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_218), .A2(n_179), .B(n_99), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_217), .A2(n_173), .B(n_182), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_208), .B(n_194), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_205), .A2(n_182), .B(n_173), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_202), .A2(n_183), .B(n_173), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_174), .B(n_183), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_210), .B(n_176), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_206), .A2(n_174), .B(n_183), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_201), .B(n_185), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_203), .A2(n_86), .A3(n_97), .B(n_114), .Y(n_252) );
OAI211xp5_ASAP7_75t_L g253 ( .A1(n_214), .A2(n_177), .B(n_197), .C(n_198), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_190), .B1(n_185), .B2(n_101), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_216), .B(n_185), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_212), .B(n_185), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_212), .A2(n_130), .B1(n_86), .B2(n_97), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_143), .B(n_144), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_240), .B(n_221), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_251), .B(n_213), .Y(n_260) );
OAI211xp5_ASAP7_75t_L g261 ( .A1(n_241), .A2(n_228), .B(n_223), .C(n_220), .Y(n_261) );
AND2x6_ASAP7_75t_L g262 ( .A(n_239), .B(n_224), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_239), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_244), .A2(n_212), .B(n_229), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_236), .A2(n_199), .B1(n_226), .B2(n_224), .Y(n_266) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_200), .B1(n_215), .B2(n_231), .C1(n_230), .C2(n_226), .Y(n_267) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_246), .A2(n_150), .B(n_143), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_237), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_245), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_199), .B1(n_201), .B2(n_114), .C(n_230), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_248), .B(n_199), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_248), .B(n_204), .Y(n_273) );
AOI221xp5_ASAP7_75t_L g274 ( .A1(n_257), .A2(n_118), .B1(n_130), .B2(n_209), .C(n_204), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_244), .A2(n_231), .B1(n_222), .B2(n_209), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_244), .B(n_231), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_244), .B(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
NAND4xp25_ASAP7_75t_L g280 ( .A(n_253), .B(n_257), .C(n_254), .D(n_242), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_244), .A2(n_144), .B(n_150), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_262), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_279), .B(n_252), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
AOI221x1_ASAP7_75t_SL g286 ( .A1(n_260), .A2(n_5), .B1(n_7), .B2(n_8), .C(n_9), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_279), .B(n_252), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_259), .B(n_252), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_259), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_252), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_275), .B(n_233), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_269), .B(n_232), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_270), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_273), .B(n_252), .Y(n_301) );
INVx4_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_267), .B(n_242), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_303), .B(n_272), .Y(n_306) );
OA21x2_ASAP7_75t_L g307 ( .A1(n_296), .A2(n_246), .B(n_245), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_288), .B(n_252), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_289), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_288), .B(n_268), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_299), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_292), .B(n_268), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_280), .B(n_267), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_298), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_242), .B1(n_280), .B2(n_271), .Y(n_321) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_298), .A2(n_246), .B(n_266), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_300), .B(n_242), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_301), .B(n_265), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_301), .B(n_278), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_285), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_292), .B(n_268), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_290), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_287), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_290), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_291), .B(n_268), .Y(n_332) );
AND2x4_ASAP7_75t_SL g333 ( .A(n_302), .B(n_275), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_320), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_291), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_318), .B(n_302), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_286), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_306), .B(n_294), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_309), .B(n_294), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_323), .A2(n_297), .B1(n_253), .B2(n_261), .C(n_232), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_318), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_314), .B(n_295), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_314), .B(n_295), .Y(n_345) );
NAND4xp25_ASAP7_75t_SL g346 ( .A(n_317), .B(n_277), .C(n_276), .D(n_274), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_315), .B(n_295), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_309), .B(n_293), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_293), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_293), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_312), .B(n_293), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_316), .B(n_302), .Y(n_354) );
NOR2xp33_ASAP7_75t_R g355 ( .A(n_315), .B(n_302), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_319), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_329), .A2(n_236), .B(n_283), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_283), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_330), .B(n_326), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_316), .B(n_283), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_326), .B(n_295), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_323), .B(n_275), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_316), .B(n_283), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_310), .B(n_262), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_324), .B(n_275), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_310), .B(n_262), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
OAI321xp33_ASAP7_75t_L g370 ( .A1(n_317), .A2(n_236), .A3(n_118), .B1(n_281), .B2(n_258), .C(n_256), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_305), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_328), .B(n_106), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_305), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_328), .B(n_106), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_324), .B(n_118), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_308), .B(n_311), .C(n_233), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_369), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_335), .B(n_328), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_372), .B(n_308), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_335), .B(n_311), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_348), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_350), .B(n_310), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_375), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_372), .B(n_331), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_356), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_331), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_374), .B(n_339), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_370), .A2(n_313), .B(n_322), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_336), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_340), .B(n_331), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_356), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_332), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_355), .Y(n_395) );
OA211x2_ASAP7_75t_L g396 ( .A1(n_346), .A2(n_321), .B(n_333), .C(n_322), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_338), .B(n_321), .C(n_332), .D(n_327), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_360), .B(n_313), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_374), .B(n_332), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_360), .B(n_327), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_362), .B(n_327), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_367), .B(n_327), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_342), .A2(n_322), .B1(n_238), .B2(n_333), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_371), .B(n_325), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_371), .B(n_325), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_367), .B(n_325), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_349), .B(n_320), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_343), .B(n_307), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_334), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_361), .B(n_333), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_322), .B1(n_238), .B2(n_333), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_337), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_344), .B(n_322), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_357), .B(n_106), .Y(n_417) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_358), .A2(n_236), .A3(n_234), .B(n_262), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_363), .B(n_256), .C(n_7), .D(n_9), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_336), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_361), .B(n_307), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_345), .B(n_307), .Y(n_422) );
OAI21xp33_ASAP7_75t_L g423 ( .A1(n_376), .A2(n_118), .B(n_236), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_334), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_350), .B(n_262), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_364), .B(n_307), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_352), .B(n_118), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_347), .B(n_307), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_357), .B(n_307), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_418), .A2(n_359), .B(n_351), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_425), .B(n_352), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_383), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_380), .B(n_353), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_395), .A2(n_370), .B1(n_359), .B2(n_341), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g439 ( .A1(n_403), .A2(n_351), .B(n_341), .C(n_334), .Y(n_439) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_420), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_419), .B(n_353), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_382), .B(n_364), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_379), .B(n_354), .C(n_351), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_409), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_406), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_417), .B(n_351), .C(n_233), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_415), .Y(n_447) );
AOI21xp33_ASAP7_75t_SL g448 ( .A1(n_423), .A2(n_417), .B(n_391), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_397), .A2(n_354), .B(n_337), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_388), .B(n_392), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_398), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_403), .A2(n_236), .B1(n_366), .B2(n_233), .C(n_153), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g455 ( .A1(n_389), .A2(n_366), .B1(n_368), .B2(n_365), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_366), .B1(n_153), .B2(n_258), .C(n_337), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_400), .Y(n_457) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_414), .B(n_365), .Y(n_458) );
NAND2xp67_ASAP7_75t_L g459 ( .A(n_396), .B(n_368), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_427), .B(n_5), .C(n_10), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_394), .B(n_368), .Y(n_461) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_416), .A2(n_368), .B1(n_365), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_462) );
AOI311xp33_ASAP7_75t_L g463 ( .A1(n_430), .A2(n_10), .A3(n_11), .B(n_13), .C(n_15), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_379), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_425), .A2(n_365), .B1(n_106), .B2(n_153), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_401), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_404), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_428), .B(n_11), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_408), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_422), .B(n_16), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_421), .B(n_16), .Y(n_472) );
AOI321xp33_ASAP7_75t_L g473 ( .A1(n_381), .A2(n_17), .A3(n_18), .B1(n_255), .B2(n_250), .C(n_21), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_411), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_413), .B(n_17), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_390), .A2(n_245), .B(n_235), .Y(n_476) );
XNOR2x1_ASAP7_75t_L g477 ( .A(n_475), .B(n_425), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_444), .B(n_391), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_458), .B(n_426), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_460), .B(n_399), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_447), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_467), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_468), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_443), .B(n_390), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_457), .B(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_432), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_449), .A2(n_429), .B(n_386), .C(n_402), .Y(n_488) );
XOR2x2_ASAP7_75t_L g489 ( .A(n_460), .B(n_384), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
OA21x2_ASAP7_75t_SL g491 ( .A1(n_472), .A2(n_384), .B(n_427), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_438), .A2(n_384), .B(n_407), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_456), .B(n_385), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_444), .B(n_385), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_452), .A2(n_424), .B1(n_412), .B2(n_255), .Y(n_495) );
INVxp33_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_454), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_436), .Y(n_499) );
XOR2x2_ASAP7_75t_L g500 ( .A(n_461), .B(n_18), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_469), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_455), .A2(n_424), .B1(n_412), .B2(n_153), .C(n_250), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_474), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_466), .B(n_243), .Y(n_504) );
AO22x2_ASAP7_75t_L g505 ( .A1(n_440), .A2(n_250), .B1(n_20), .B2(n_22), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g506 ( .A1(n_471), .A2(n_153), .B1(n_235), .B2(n_243), .C1(n_250), .C2(n_249), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_437), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_488), .A2(n_473), .B1(n_463), .B2(n_462), .C(n_431), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g509 ( .A1(n_496), .A2(n_439), .B1(n_451), .B2(n_453), .C1(n_445), .C2(n_470), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_492), .A2(n_439), .B1(n_446), .B2(n_465), .C(n_448), .Y(n_510) );
AOI222xp33_ASAP7_75t_L g511 ( .A1(n_481), .A2(n_442), .B1(n_433), .B2(n_435), .C1(n_450), .C2(n_459), .Y(n_511) );
XOR2xp5_ASAP7_75t_L g512 ( .A(n_500), .B(n_433), .Y(n_512) );
OAI32xp33_ASAP7_75t_L g513 ( .A1(n_491), .A2(n_446), .A3(n_476), .B1(n_234), .B2(n_28), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_482), .A2(n_476), .B(n_235), .C(n_243), .Y(n_514) );
AOI221x1_ASAP7_75t_L g515 ( .A1(n_505), .A2(n_222), .B1(n_209), .B2(n_204), .C(n_32), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_493), .A2(n_249), .B(n_247), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_486), .B(n_222), .Y(n_517) );
AOI211xp5_ASAP7_75t_L g518 ( .A1(n_495), .A2(n_209), .B(n_204), .C(n_247), .Y(n_518) );
NAND2xp33_ASAP7_75t_SL g519 ( .A(n_480), .B(n_19), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g520 ( .A1(n_485), .A2(n_249), .B(n_247), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_486), .A2(n_23), .B1(n_25), .B2(n_37), .Y(n_521) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_489), .B(n_38), .Y(n_522) );
OAI322xp33_ASAP7_75t_L g523 ( .A1(n_479), .A2(n_40), .A3(n_46), .B1(n_49), .B2(n_53), .C1(n_54), .C2(n_56), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_477), .A2(n_193), .B1(n_60), .B2(n_61), .Y(n_524) );
AOI21xp33_ASAP7_75t_L g525 ( .A1(n_505), .A2(n_59), .B(n_62), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_512), .Y(n_526) );
OAI21xp33_ASAP7_75t_SL g527 ( .A1(n_511), .A2(n_497), .B(n_479), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_508), .A2(n_501), .B1(n_484), .B2(n_483), .C(n_478), .Y(n_528) );
OAI211xp5_ASAP7_75t_SL g529 ( .A1(n_509), .A2(n_502), .B(n_490), .C(n_494), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g530 ( .A(n_513), .B(n_506), .C(n_504), .D(n_494), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_510), .A2(n_503), .B1(n_507), .B2(n_499), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_525), .A2(n_498), .B(n_487), .C(n_506), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_522), .A2(n_193), .B1(n_65), .B2(n_67), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g534 ( .A(n_517), .B(n_64), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_524), .A2(n_193), .B1(n_70), .B2(n_71), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_526), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_535), .Y(n_537) );
NOR2xp33_ASAP7_75t_R g538 ( .A(n_528), .B(n_519), .Y(n_538) );
NAND4xp75_ASAP7_75t_L g539 ( .A(n_527), .B(n_515), .C(n_516), .D(n_521), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_532), .B(n_523), .C(n_514), .Y(n_540) );
NOR3x2_ASAP7_75t_L g541 ( .A(n_539), .B(n_531), .C(n_529), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_536), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_540), .A2(n_530), .B1(n_533), .B2(n_534), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_542), .B(n_537), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_543), .Y(n_545) );
AOI22x1_ASAP7_75t_L g546 ( .A1(n_545), .A2(n_541), .B1(n_538), .B2(n_516), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_546), .A2(n_544), .B1(n_520), .B2(n_518), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_547), .A2(n_193), .B1(n_73), .B2(n_75), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g549 ( .A1(n_548), .A2(n_68), .B(n_76), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_549), .A2(n_193), .B(n_536), .Y(n_550) );
endmodule