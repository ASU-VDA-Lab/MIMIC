module real_jpeg_29684_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_43),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_56),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_57),
.B1(n_59),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_5),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_87),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_87),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_87),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_8),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_57),
.B1(n_59),
.B2(n_79),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_79),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_79),
.Y(n_190)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_57),
.B1(n_59),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_11),
.A2(n_52),
.B1(n_64),
.B2(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_15),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_15),
.A2(n_61),
.B(n_65),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_57),
.B1(n_59),
.B2(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_63),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_15),
.A2(n_45),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_15),
.B(n_45),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_15),
.B(n_81),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_15),
.A2(n_26),
.B1(n_37),
.B2(n_201),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_15),
.A2(n_64),
.B(n_217),
.Y(n_216)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_17),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_22),
.B(n_105),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_99),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_23),
.B(n_99),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_53),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_54),
.C(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_25),
.B(n_40),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_26),
.A2(n_35),
.B1(n_38),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_26),
.A2(n_101),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_26),
.A2(n_117),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_26),
.A2(n_37),
.B1(n_195),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_26),
.A2(n_117),
.B1(n_190),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_36),
.B1(n_95),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_27),
.A2(n_36),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_28),
.B(n_48),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_28),
.B(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_29),
.A2(n_45),
.A3(n_50),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_36),
.Y(n_117)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_42),
.A2(n_111),
.B1(n_114),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_45),
.B1(n_73),
.B2(n_76),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_44),
.A2(n_64),
.A3(n_76),
.B1(n_218),
.B2(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_45),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_46),
.A2(n_47),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_46),
.A2(n_47),
.B1(n_176),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_46),
.A2(n_47),
.B1(n_143),
.B2(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_92),
.Y(n_202)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_69),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_66),
.B(n_92),
.C(n_93),
.Y(n_91)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_63),
.B1(n_67),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_60),
.A2(n_63),
.B1(n_86),
.B2(n_140),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_72),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_65),
.B(n_92),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_80),
.B1(n_81),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_81),
.B1(n_138),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_75),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_75),
.B1(n_97),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_71),
.A2(n_75),
.B1(n_158),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.C(n_96),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_92),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_124),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_118),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_116),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_111),
.A2(n_114),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_118),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.CI(n_123),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_163),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_146),
.B(n_162),
.Y(n_128)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_134),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_134),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_141),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_150),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_156),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_159),
.B(n_161),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_160),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.C(n_166),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_247),
.B(n_252),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_233),
.B(n_246),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_211),
.B(n_232),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_191),
.B(n_210),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_171),
.B(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_198),
.B(n_209),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_197),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_208),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_224),
.B1(n_230),
.B2(n_231),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_223),
.C(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);


endmodule